��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����`��B�㓪F:��ew���@�C�k�.U6�vά1�xrl9��Sr?$R�t��M��~3pwd��<�i��w_�)4ޟo$#)����4F�1s[�p;��Q�!�~D�����ӘFy��P�1�ɂa�Gi���h=�T�?$��0�=�8�oN�l'ߧ��S��P0T�\"��6}8$�ل0n>+���U>Ö��7����q��?⨴PE�����et�/r&T.7�@�uv O?�`����+���#��F��O9l.=h��`��]���Z�^�������hğ��v�(3c���7{������;���Q������2��˖�+���i���}������9ݬ�����V7ARʁ&�D�5�x�p2�����!���Ɨ�՘tޙZ�d���o��c�k�f��ʝ�$��b��1ʤ�n�X_���D#0k�i��mf
v���_����rya�~O�@u�����u�\�]��=n�D�4�ڎ��6���$M<~?�xdP�sҊ�N�����OG��l�v��P@�o�}RBKn�#9�5
Xx/�	�jR�ٻ���������	��tdg�������):���![��%K�L�'��K�9�:1��0[�(�.����4[��n��$e})M�&?��4�]1��13�8��K���X?�TDj7|���R$��ʨ�yy�'i�b
�R�+0���YVW�G�ANД�o�I���?H'엇��&����:��m���'�rr+s/�9�����{�!��5V,>�AP �la(��`�c��ˇO�?�-ȓ�L�6l:\Up��ُ7	�I�M�k���L]I��&m��f7���:���ܴ�+�,��N8{Aa���iۓtEP��m9�b ޶g�qe�������)�(F0K}G���ޥ�Y;�\y��v@��ܵ�3'8r��6ڇ�\�+$'��A�e- ��O�o<ѩ-���|���[Sw���*;3�,�xLV�%vi~�2,� Al�=�F�?cS�KP�3�`�a�/�I�`�>z�dW��="BY	ᡶ' ��˯`R8� +civ���l"M�������L8�\�dD��M�x(㙾6�����`����FY���԰����Kos��	3Ë����m8�8��W����5��o0�j��N)�ٗ�L:�t��;���8����J�Ԧvka��a�x[�5��a<t�zK��|�1�?�܌�»."xV[�G`�����Sm~ɶ�0��Ĭ1@o��pK"�Z̫�hS��:W.�iLw,��R��MZpQ�CQh{�������Un�������MQ�"�0�xn	�)oL��$���L1�|�v�����'�6��ޤ�i]��jC�kg�Urx��q$pk��"��Q,N�o�p�όi��R�6�m6HI�k�	|���+�T���Νh�"��|���X�
�����`��1�x�\��
!C��\?e[~�q�BH:+������C�E�dk(-�?�<q.��ֵ��Q����{ٺs'�?��/���x������=Q���>��Y� ���Θ���J:�I*ō�<�IO��,��GƮ=%��s3��Ȗ��p�x��];&3�'lT#I䮄�܆36����G�āV�����&	�@���Ж���S9����p�.n��ov!(xs��u��w{� /�ʀ��"��!�ޚT�(h����?=ݭm�I��G)}����)˩�a�p�j��?u��M�'U�*,v���j!f�=\^^E�O�Sc^��'Bi^�K4�v�1���Z ��@)Yex�	���գ(����8D (��7=Wq;��!���-$��V(H��GK�Z�u���.����KR-���h���E�nF��Ѩ�1@���-�@�Y�<��S�D�W��>���P�M徾4]��՚�0)����nC�b���V�����Ly�-2p�S��r-�G^������F`���_q8&b:&���4\}y�:�n�	��"̲�k-����a$Z{L�Y�$�@ז�}��h��GQ]�&��RVKNv�K����?�݊�ώ=� ��tƝs��I���1Ԟ������p �7���s���!����"�]XG� !�0()Y<i��^t�� (�Z���ۦ1!�bQ�PP)���05wڭ�1|b�?��s����i���=�7J`�LbR�İ�	FoY-�}.��M)����W��	=�G�������%>'���v�_x��֙���}�&a�P�b(���:���ْ=���'',�
-e8T�q��w����D�����$릟��ܡ@-��G�̨��R�!�[���47����j���V�f7�4;rӜgǔb ��w�l�7".�����F�L�����b�T|8���~��w��4�^���Ǥ\T.�J��30u#��'�(�>U�߲;��DЎ0�|Z	��:Y·�W'��m(M}�xݓ�� ���GL����2�"�i�ț�y�s^�t)���t� $������}*V����T�1!���-�E#p��$�q7y���������Kx�0֝fKQ���QK���C��Tt�#l�B0���/Q9�yn��s�g�+���~Md֔�W����O�-qe�~A��II������� ��2�U�v�	R1���%m�,Ti<r����F����AQ�����i�ͅR�P^��;a*ޯ�f��v+s�
G*c������_C�r�u���T|R�Z��X	��SdP���"$.�e��*eQ���GW���C�c��(��3�kϢd��U~EV�4f��^��4�P�od�hr"��L!�1N���r�<e{��t	�:�������ʟ��K��C���v�"PԴ��� �_׎��ז��0f4xk�BK2:bq����qs���[��2�I��1w�2Q})D����"��"ۯ(�N~��TA���;Ln���l:R�{�������A˸�+jUe��
b�ͮ���a���I	��枘��n�h�ɡ�&� �e�qc��x-vչ
^r�c����*���P��h��?u~[���#?����C���*��.ֲ0i(d���B��t��%e�A�Z�U��'A^��x���j�&�높pp��>P�B��	��,�<�� �p��̧���y9)�l�;�[�5 ���DS��DH2qr���؂8����w�c2(�%��Y�W _�)��+�/� �1�G��O����LvrGi�`@��|�w+�g�!~>{���mQ8��� ����5�b�AY���|�i4U���ٞ,A"�^�b%K�"�P�wv�6������s���x��i< �P �@T��=e?��[U��٣cZ�{)&&��X�h'5q^L�2=%�*'���F���_$�
�������f@*��g>�÷nCR��F��pNw-����t"2��SC	�^����C�<�&u�v�(D��d��i�A_Ô< RP��2�E����e;�Cv������V��D�@�=�l�"�Ϻڽ����mn꾎�`��~��2>W���-%���{mz�/��>S�+��A\Y���X��e�H�/�A6Fy't�'!�ˢ
�Wi��>����J��9}�_����}GxqT����56Б�H&���r�P�E�a]�׻��TPT�z:eS�#m|��zQ�����
>�}+[�6�	~$⭪������h%})ն��PW�C���s��pɏ-�(%� r	���ۤ!P��n�����u��T9����L�@�/%����BӍ�3��+=�Ci0��A���X��BNj{v��0-/�	��5Va0���	� N�J���n`�U��9o�O��_��I�C�?ŵO��t�G��]EH?\�L)sE Z���o�H�<_(rNC!�x�:�{�f
�1Eșk�x���?(F�R����R��Y�SH`2��;�PZ��S�ɡA6���#sn-�V�ɵ��x�D�)��(��*�dC��7gXt�C��?x��O��Ǡ'�*�:M&4mv��+ctb?�&�����(�\�¹����$FB^��H�b�-�6�4� w�����ʼ֩�q�@}�"�4Ty�O9�X�`Tm�[�l[݌�63i�9�;6�c���'D����
����8D<\�`�q�M�����h4���I�C�a{/���1�l�Q��v!�=��V� YG���w��yb7$Ǜ<�zs���Pf��&GpSO%���q��r�,h�

��<�?��������@�E���[�_XV�i��7:{��  ��F��e�2g�V�ޣ��u���7�6�QǞv�aƬ8!�<�ࡶ�u��xia'�V��-��Kj'�V>r5ʱ*K{���j�&c0׻F�1q�nM�������T���.�N�`�����vw�1� }���'!@"���H%��h:\g��;SM�X1�~z��8ܓq�f�``��-�edR��V+^�ǥ�0�t���Eȵ�z�H2���O ���M�X:4S�����LBJn
)�H�{+�L\ǧ��R�O��@m ѕU�N�����^���([�VV��?��R�ބ
�t	��!r#�K�9Y�k�)s�:Fi�������˯V�M���A'w�e�/�T���@������U�9����R�-aS^���$��/���
��jw�)����8�X�	Xv_�뭬5�AR�6y�I�ξ����� \�o�[#��V)���0]r~|z9����F�ek���
���(���b
��]��+�%�R�V���U�	g<�g�ցW�1xֿ�U�K���V��ǹ��������|a"W��zc0����n�+�^D<�h����Jg!�['і� �����#Ό]�Q���\�~��u�������S�Y�� !G�\
Hr$��A��`�i�����ӿ��!&��17���m+d�[�G��?� ��8V��z�l�A�XǨz=tfK_��O�|s��qZC���c1,��9����5���h�d2���~�l�yx\����@��Ѿ=E�$���d�y��=���]�۟��(�~T�g��'b��}5�l�n7h��bCduѧ����B�tt�Z�����Հƅ�0�I�f.y�q����'z욗`V"Y�T}�rw*ޗ�vl�K�k�r��$�H�t:m��5��a.l�E�,_O�I�D�w�f���g3�t(L;a0u�� �^E}�7{غ�b0���B���/�?F@q�����B�$���Ƙf�İ�(�Nr[�fb�� ��D���q������^��)*_~���s��Q`��5���8�C�(F��B��bg�r ,>�C��#E%�m69��]Ú�B+�6Ro���I�F�y��I�t�o�����a��?�c������D��>�	�wAۯ�Pxc5��'-�:^4�	���.�z@T�j�*��4��i0���x��Ȫ���s$�ޓH�q3L.�]S��q����Q�M|�Ϟ�x�z��t7E���������#�x�o��&M��6-���_"՛-�i�d������~��3նF�N���/7�ꅅ�dR�5�5��״����R"��n�_y�ۘT��:��������-����f�����g8V�M>��_������kF�f*�^�]�G�ߋ����e�h�ĦV6�e1cf�*R����N�7�G:�",)���־4�����l�RIzZ��KOv}Q�[����5�n����������tnx?I��y�CC	H_ϟ��E�C�`�Qj{���U�
�3|*@�P�c#����Ս�$��*�dU��+bL��IHŚ�XW�,5P�եAB��Z*�YR��q[�!�R9�kv�e~�~p�^$����GR�OR �݌��U�E���L����V����@b�6 I���}�X�;���ݢf$���2�DS��N���"�o1O�Q��RP<��vM�#�������_��V����z�+̵�v�U�����S�[V`��-4!d,N^�0�'1"����
Ɣ�~ ��5P4R��ߤ����.��C}H�Ώ9T�2%	qV��Y6��;3���i��'In�Q���a"�Q���E�Hj�m$��B1�:�)	�xqu��_��mV7�*�����Eȱǋ4(RݙQu���}*��,�CZvwN�|��*�X|��z�O�95l�Y�y�T�iH缉E�=攰��0���)���@lq}�-��L��!�)��>����k&
p����K%^�]� 5�*F
�z�I^�l������UHF��<�E�[��ִ��7�p�տՋ`�H;��
���E}��s��\L��?��4�u�pL�7�����P���Ӷ�e��ޮ+)'��rr%��!&I|G��lkP#��V�Tg��g��AW�b���V�����
i$�ى��}�I��&��4<�Zq��F�/�b�dvxx�뉂�j�L�!�K̦�S�ʍ��g(��-���D�;N�� n�T">�6���89lH_)$�!�����e$"���ZP	U�^��zF8���o����s��RH������pɩF�K�2��*��&P��^�DW��!�������˼\K0aB����v&�ت�[ ���XI+V�=���Y�����wI�}�ٹ��]8d�����{Vo�<Q��o�q��n�e�,�7���sKX�{�ℛ�C� ���Dÿ�6V�%��H�''Jѡ��bo�o1 �2[�qu��_�c��,�!���q���b��t��u�	�����6�`����k��~%b �4�2�Dؖx�Z
�����{C���.k&@���`m�m4��3&��s*G��M��6F�E:�s��R���eب�����/ �f?�W?��
���聐��l�����E��~N��љz�K���4�^�T�"g/S��ڛ�	���Qt�j�+c�]��eq��D`?j�uj0��s����P�xmeQߓ̾��ȱkk�ӱnC�6Ro�Kf�w�;�uiu�K�G�I�p�z;�ܭ�c�\��m�����ex%]�p�I՜��ڠT�"�;{���c�J�=��xYR>TBT������C3:=z�U�ӵNj�4<����t��_6ʦnz��Z�&��I�=���\��a�� b�̅�$";A�;
�N��6�1Ui.;�j�y�~#��0g�$M|ژ|m���w�	�;���]XFo�cF�����,#g[�&@\ݦ��Z
e���FߕLՅKc`��x��U"c�@�ٜ����[�6^�Am�<U_��]��}w�y�6�)�~� �\/�1��.zƋ��6�$��.#�8����YD��Dg@3��otf	u!�)+	���R�m���+��,�Ը]�.3&��ط���=����BO��A��`;�ϭg���$�B\v֤�E���C]��Zk�]�q6��fVEE�G�� �Y��#�@O��ц]�����׉�.�U��(O���e�+��f۸ʧ��4P�I�M���y��CQ�]�o�YHLOv�V{+�+�;ZsϹ���D,�[�%�#ߺ4ɀ���H����ݾ�+@d�5�LBK�釻[�ܤ�4����Q|og�����v����L�&�%�*�G�����c����އ�eKVo"iGiѴ(Ҏ�(��7��x��2�BUH�M7Tª]����[j��<pe�=9�b�en���'��F�፨r��
~��s@��B��Y��-^��hn�g�<+�_;�K�]���j��֞��}~��Eo<�A����ӗL�_�G ��u^�3�����e��F(�'`SP�T� �$��W�u�{�B	/���d��2�.{�-�u�����%(��^[�,;��qS&L�i	���m*҄j!��/[�	y���;A��^�)�rs�Ed����C`�s�2Wb����@����Ŝ���((�*[�}�Ú��N�����#f7t>5ǧ�R׽~,�2<�3[V�U�A��r��7j�i��E2�~���>{�����.a96*��H�*���R���%0�����ĭ�{��k����)�t5
p~NDTp�N���{���	u$n���Uh�=Oߥ ��"�����b�u��9b����;�(?�)�"����z�2��G�?�#�<S�t�W6)?O�`�_Y��eS_z�3]Z��Cq�p�Ŧ��h�s��L!���ht.��q�z��S��W�$��(��w(��cv�ϔ'�'�ahQ>���&Ln��E�ՠh	QOY@�*ИY��P�;Y~yg��{h=?���h��ǿ����6���11~v��B����Ao�cZ�K� 1�s7+~����$���US[Qd��#�0$-��#*�-4(%�~�v)w�5�ȣ(X
���E��z�\�P+�7�E�=��zAUD��/���8):`��^)�_�D0��暊��B<Sr:]�{[�
��ۏ�n��F`g|픴�����+��+
'9R�'Ł,�"ӏK��=�.U���"w�M �&�o@)�=`���!G�(�F�J����C���kq�"�V��4>�o�.�2�h?rL��,o$����O��zh�%{k�:�������")y�-a���*p(!���l��ٱK^���0�]m��&�ͫ�h>�,-|�2�u��tcZ�� � 0����0�f!��,�>�Ί�'٦�N����o�y#('CT�����{���oF7��2l��[����=�bM`�h���l`*�\�����]��O�a:�\5az%w�?�+:�OӁq���n˸ǭ��f���\�P�Md>U�0�ϱ�L�i|	�\p��W'�}q(�GT��ts{�ٜ����*I�e��o���2,�����-y�m�5��,`�W39�����7��������?���9��-jԒpnӺ��)2oR�������	��a�Φ�D�"|(A �5���V��&|u6�a[9��J�z۰�%E��̻����%�f5��n`�2;b�v3,�n���cfڤ騝'����Ҳ'�76 ��V��B�x@n�X����޷Q�A˓�#%~�ʢ����4 ^.��_��~w�Xg�A+H�MP,g-�:j�|�X��|.��j;�/��1B����
���Mϓ��h�*�j/_Oy�@�w����'Ί���㌰�Y�t��Ga-�l��k��8�%ߥ#�ʜ�ΒOw� X��{���D;�O[��J!��:=x�|fKl_C��'dU���*=�Z)geo�o	K��/��R�F�Ik�� �ԉ-ҵ�!��r�%���[��H�����I��]�t��u�;6�=�V���|��ھկ�����[�.N����ӽ�݈?\��NҴ�4��4�����7>�`�z�}1"m[>$��*?d��9�E�V�B������G���R�q^W?-�
�r�r�ĉ����� �VZ$(;������L�b,�7�*n�+��n���a4�[-��� h�j�_YZO���p�@��<�s�A�%6�����l�E���b�p��1^��
đ����m��q ��g8oY�1��������[�M�9{����P��u)�pu�D�cԽ1�Z���Q~vv8��&���~ݢ�b����gY�O��"��*�NA@n*QGLV)�~F�R">7 �:�m��K'�w��Ke�k����=�:η��Ŋ�)3��!��_���Ş�0]�h�88m��r�B:kӛ���W�K���sK��Q>�&5�D%/����UW}�ZZ�: ��{g�N�BǕ��,�Y`5U��{��C_�/a	�E|�ԁђ��?ĸsW�����)I�������}BВ@�JF�T�Ft~K�]a�Y�U0W'Ѷ�E��*K���3��E�{y�����#,0T$��5n�]H(��T��|j���h�_)�G�$���d ]x�e�rb��#�����f�Ƣ�`.��Y��ɟ����M�	���S��å%l�֜���mc�Y?|��Er���w�EJIp��G�G�νX��hh(Ώ��usY�3�J"�r��'6�3���b���ǝ�q��*��GP�*�D�cM4��%i�������biw9�_�kV����T������
!樒$Ǉ#L��ܡ������]q�ņgEo6����Զ���:��l�"���X�֗�����=�?e�9�Msܠ�0��m]�D'z��`4��@��5��.��6/�J6~��1���O]pb���1��n?���$��LB�� m��>�}룾��n��ȏ�N��>��j
���B`j]�Չ�RB��7�aY����6��c���`#�{~(B=�)sIH�QIY�*�5�ܖg�����i$Y��MC`���H��s�~W��7�.���<v�dX��)2Kbe�d�%�bؐ��8�8c�a*��� ��K�����"�އ���t��Bd��{�����FY�@2��cf۠�m� ݙ��,ҴʗI�㗥�#`UM���s~
���B�G+�\^�R_z�w����ɹI�,UH���D�E`m�Eo&.�,݊��W��?��(��v�!ؤ;M����dG-�2 v�،���|�/�,ڻ��i����{�^�]$����G[��a�
ӿ�G�ư�=f���)���2f���MŸ�gH��^��ߤ�%M��~#R�f�Z��)`�L�o�~�l����u� xEyπ�$=���y� j`5cd껛k[��XҖu���t
�8cL�'yLG{O�kLQ��~�ݖ���I���]�\�r`ʕ��u�<�
��c�i�,����8����a�W/��R������Z����CJ���:T�Ǹ_��:~~����ö��ѵ�vR�x4�<�醰�V}�
��p�S��yN��z\-�y>w�;e�x쓥'LC��F�EbU�t�|l=��+���'`0`�<Z4 �gû��L���	aT�Q��ƻ*G1x�M����lJ7��>@�0܄{+�6���@� ����r��v����<-}��P� �	�;�y�F�)i!����Bk���h6���z��H!Qf}Q,b7��!�S�2��ޠ�Y3`�b�k�/|��s�I�lP���?����?&��Mϸ���n_����]-�%�DqK Ȥmo:u ��]i��Sb//�N��p�Bk:1E�7 �Q K�+���5Й�("�LżL3�3�0ܧ��O	d#I8��?�C�[c�Q��e�����c��T�Фn�̗�����e�EI���U8�Ͷc���N����Tj���<^�����{����t�|��0/�,� h6��rFv(��Ʊ�����V�h9p�~�6S̭ͯ>fk�*"bT����oK�c�g � t��Q{�2,�|c��jFQKS9a��0�n+RÏvQm���RmT�{p��Wm�yٿ��\.��xV��5W�'�^�3H�s%e ˣ�h�b9?��ู��AU	�y��7�\v��XD2�҉�Y�̯�W�l�����2��������&]Ǡ'^����h�4�[�#����9��C49u�����&S�i%���:����_=ɰߧ�Kp�Y�{��g�x~�ZSm���a�C�,�`r��Ԑ�F�+$=��o��1��E��������b;zǌ�Р�ɒ=4{:6�i�N�,���sƿ�)�g��ğ>g�tf)�?~���h�Si"ps�n����wL0G|sρ�:&�ƣ��;~ɚc�Jcq����(�m��(�V�`����i��XQD��t��2���}W3�{��a=�;$�a%�n�$%��P
 Z��Ĳ*�nF�OG�O��0V�qw�>�#�F� ��%��rIƲ_��~���Tq0ڒ5�I0�,�-�ԨY��ÕwMӠD�r�S�s�Ѧ��\Ktw��\(�ؔm��SY�zݥo�ȗ�`���Z�*G���e�;���)aY���	��)W�eZ�{����v�w`+�K�b�~I�u�O�����IK�t 8���nʑ��,�{���TΖ1��/��0ej����D"L-�p_��������{bK�ڥV�����dpufʞI��=�z�X��/��ܳC�B�^��Ot�R���!�U���}��H�({��-wZ�ە6�cU��̂&?�塳V�3��%M��\���y�87��-�]��iծ�Q�>Mm��D��=&�� �^xv`+7�F��Ty��J�>�s,�-��6_����:�l�'PZa�l�s$�W�&��YYFEL���?��tY�����[�v��u7�|� �:���|��Vj}� 6^L�6��_g�L���D������ІOiI6 `��Bڟ3��F�ذ�S�H^�
�{Mњ�:6�R,
�M�wF��jjZ�,�
,7]-S!��NQ�k��5]1�F��Č�#��n~2�]�8���r���$��0�$o��y4�?��߿��9��%KӇ��_6ɍbEp�ͯ���R�<���� ������Y���Y�J?e�h�J�����E
���R	B *�+�>;]V���93��{���?K������֙)_I���i�	l�6t1���m��"�kS�k��;�o���E��U�]^�*_F�k)_�RX5>�����|/Ha�vRJf�ه3����bF6�C���u�CҶ��Z=T���?rq�y{8�h`��X�����:�&`�!��39�<��ãn'��F�ۊ���4䌘�B�7�Y�*h�q5h�dO��-� $�W-BVܫF_]�����'�=5�$�<�G�J�����w���4Vp"сu�Q�H�\E�m�/���nz2�|����P q��I%�Q�e J��}	�?���aa��P;�,��dXĒ^R�o�"�� =	��������U��9���]Sf�����nʬ���m"
��	Ig����Q����~��� ��s�d�O�4�$�Qd�X��x������M�2�Ĥ��L��)���p|����%�#�^��q���������ne�Ԡe���`��T���:��O���r��B(Ptt��vaT:k�E	�\�^ۋ$����۫�G3�u�v��b쳵G�:�!p��L�e��k����T�Q�ݼi�*c�����Vu>�s)�}��4/\6�>�v5X���^�;c\j�א{.b��<�;��v���@8�ȕ�4 �Χ�Y !����La� ��j���'��2��?R˾@��	5ׯ�����@�C�*�ڧ�x[R��b��7N�wt��.2�=�o��R�=�kO�7��6�T�Y���jW�R�Zf����)ҠS^�A�13Lb�P�Ij����am�[���H�:�HV�7�\'m���<d��i#t̓�����}�qs��A�k�� f��U�<��>¿=�~�z�{y�@_s��)˔��	o��)��g�\��}��; �p2�|��#� 	��JW
����{�Y�/�f��I�hH��/��c<f��Gte�v�3���
k�Up�T���f�-�z�|�QIe-�������≌����uޫ<���P$R���+�΁v�UnO%*��C��MD'�(���J���/>�t<1$n��<l>&ЖD��t�S��{�s���\��@��­�"J0I����D�����*{��e���c�WQ�a�U.<�:W5��!��q���/D!E6!{��`�F��C�E�+�^6*9+1v-�(s��d
�n�u�r�D�ϵ�s����.��s����#j�0�P������b�淂����?�����Я�h����f*Y�����@�V�JO��,����	>��b���?�d��j�h&��~� )u�^?���/�W�Iz�<@˃��h0�fC�K���0o����"3��|�҇��6���Ѣ��`;����d���Y@���X	�@��H���#b��'��G_2�5
;�y����~I�Ï�v�Ƞ ����ۀ��H�`CZ��K��̃v4�E��SU�� ��Ow���!㩗�z���D����m�G5$+�P���h��}�ۘ�lrڭ��s��U�$�$���ቭ×��ͦ��.8I�y��g��~~��R�ʤg�T��!<���p?aT�*95�j�e��=�מ��ձ��ͤ�wc���&��t�#[�d���k�8�h�O)&\��-�x����)��h�eDr�#5�H��q�C�"�*�|t�?��l��i��s}����M�9J�g�`(�Db�2t����.[s�	t���ī�Og�@FAV�z���iX�nc�K#a�t	e�|��l� ��p�xk��F_sYm�޴f��Ye��=*����J���|l P�/��	==�*(jjA�Zف�C&0�z֓���4@qț��:���ʌ�1# l/?�jL�;ܠ�h�b��q�j�uT ��r��"V%�u���9��ˠ�X��3ZU��d��?��Z\˭F�v8Ȫ��J+��J��K6e1%ܔz"��?�%��'fI�v�؀aU�&���R��q���h�r�Qd,���2�˹�H#!���km�)�3(	�o�C�v�؀��߸x_�����5b�Qu��Ŋ"�6��;F�`B�����Ŭ-��M���v�4`��ږ���
�6iR�<�m�I��c�����J�o�����>
�$�l����������gū��	<�������c� !VD5F��;��=5��*���z�	/��S}���+-�v^�D�s�5��&�=Zhȣ����+� ������1\,�(�5��+����f�V�wh�<�V�K�h�����$FWyu�q�Z�+G	��7ձ��ABz�z��pq��~HVLe�1��.
^��@�����No��1�<����o�� "/��1JA���K����O��Q�;�+x��|rɢ�-�t7�VɧWg5:C{G��$)��簨H��ͥ+/�C�'��&�+:�w%W�T�y��R��T�
�3x͊�*#�� W�&�Y-kû1�Z0K�å�P��;iz0��u�9��]�h�>����w��P| ��N:�U�F��&6�B��g�뉻��^0�-��h�`��n|%/k�������j�&�1�J��������Y�hT��A��riQ�)፳K���s��1k���ŀU�o���������[��::�*���~��J�%�4��(�1�d�UHA��j@���5�r�g�x��2L�6N�*akȫ
8`��r���`u'��� Ob���͹s�Y�[�R���[���AA�;��%�H��v�Ϊ����O"�`ַ�
[�y��3�p����#�j�� �g7��/�ŐE}D/g���)a�z��2�M�
<)�[L�I)^5�v��̞����&	�-�w�K��T�&�[r�%ʔ�Ux�#*�<^t�')��B�x5+�g��k��r�y�Tz�6�꼐_L>�⚢~y.v�]X�k|�ka�we��-8f ����%����D�=n"����?��=�D�Kp� 4����Na
��Y�  �����X[�5>�R78Y���z�m���<^%�t�;	�I������K0��jp�!��oD�_��G�)���a%R��c,ƱA�X{�7����	�W^�V������
�.7�)t��E��@�E$w_��9��՘(�fSm��yC�LҤӼ\���Q5�k�hѾ�t1Z�
D�(U�B�܁{%腗�Yo���3�*������K&�Z�	�.@���Ŷ�L�5��}�`}(T�gx_�*�:N������Q2������n�����:����}�l��!���b��:�N`�C֮mU�}��y;&�(�<�:.�E#����4!>�>_�ܞ�����!�c�����Mz!:����΋ɬ�%���Oe�,�%Î;�,e[�=���9�DkA�L� �)u�@Щߧ��UuQ�c����a(!w�ugd!S��>@aJ��^�<v��
��/]�=(u���[I�`o�󮅵�~��3R�K�J�%ܽ���ܳ���(�
�?&xr�md�1�nz��,U��#�ǯ��֮�+aS[h�C#�60�O/;X$en���0�������=w����G��p߃]�?e��9b����(�z�(��vJs�!�+ȃ}����n&L�<#X�#�<o҆3�cDQ2n��$ߟ).��YHL2xb���\�(����D����o�_�u�<"�*�c�,�ٜ�l��s7�*ʟ��=�N�b��{:��CK�~�d�%�Bz�qA��"}� ��w.� ��l3O$tJ�����ho��׀AB��7�)�Ň��n��>�c0M�uʬ������&����_*�Be��(n�n�:\���KS�5w��R�{��ǔ(,�+�Į����ߣ1w����i���m2:�����+^Kh�.g?q,/>�!GG`��g����H�@�_х����N�ɘ���~r\�b|HQ�گ*�tN}����k�B�����i��͸�?(�g.ì��4��?�vٰɑ�ԅ���ܓ5ʑhr�6K�e~Qҁ�['�Iuk�_���
��YC��=J�gH�&Ԙ�ѷ�B�.m;�f�Z�JoΊ��R����Zw��s�=yS���n�y���X�tW�*��ѥ:n�ӆ���;堤� �\��=�ϫ�}��o�Э��m4�L��ia��Z���m��O%���~�?POqz�����j�51�Vn������X:��A�a~�P����nA��}�u9��E˕�2F�8���>ǌ=�q����D�����_.�Bq�%�*Lg��H�����6�yY���%�G"�ȓ�[��i��?��6=ůٌW��uJ.�g��^gk�tUlOQ�0)�!�;��E0�^�b�����̧(�nr��w���˻]	�X�P�AIb�Z�:ѧ�j\��������7�h����(�2W,�TГ���I�!|@x�@�Vi��V��O.57�y7_�( 	�M5�j���𚨼	H�߅u�vK	��əIrU�s
���]��O��~o��׀oU�_�ձy��8�{�]��[��^���p� bg�̑&�7���H]�v�����5������XL�/��祱�H���a���j,��3h-���]o�q�9r����w���6����C�qߛ� �g+&m����I��kL�����^�R)4&eV}� �A��O>MD��D�˙�rQli�@��:.}IQ`���0oܘx��8����(k��CNaK$���1m����[�c���;rs��/Ĝ����^H}|b��O
��p(��r��9�V��9Ѱ��sɗ�j	�y�j��m1���]Ц���"��C��MkE�-�$��"�Z̠sUN�˩�(pVS�Zn�.�B���U=+�y�ܪ�C��>#��Ue�w|��а���9�m����1��C bc���eY��[?~{Yn�sI�2��_�O?/�_3���g c�Ą���S�Hq�%��H���]Ʃ��������zUy�h���N5ŶZ]��Ĩ�$�1Ӊ}����H/j` ·�4L	���б�cb����ӂ��� y\��V�2/Z��a�t���ױ�D�@�&<���^�Y�J�Y&��z���9LGs��}��X�ʿټ�f$�A��l�'�K���������=1��r�k|���m�NW'9;��������s�����5�pb��l1K�3*�5�Z��,夙}9������Lh�ɥT	���"��w�Dߍ�؅�T�{I#������� ��r��	�'�R	�@t��,��_��:~�,�u!�t���O�(��m��t�kǳl��hX_�VS�ŏn�[a���H5Yd>�}��^|6ą�- ;`���LB��!DF����w	�B��-nݏ(���!��ݦ������1�F��2��gv�O���Z�@�R<��f� ߠ)Cè�)�ăƣ 9	/{��Y��q�"� ��<\�0�Q�կeq�!"���`_��,�[	?����W�	�8� '�۽p\�Zo���s��<a�<���3���9��Q����$x\���΀��!��{�!�U]��z��ri<S�S�&� ���E9��[4$k	Ger�uxxCKЬ� 2Ti�
$�C��6�o��?t�Z�$���z{䵶(o�9���@�7������;Ve��#-����s,R}_���_%ŧ�m��=�5+bP�&,.)^1�c�:�����+���H���g�����A"��e�ٽ���x�$0g�.�#!����!S~柱��?����谵j�z۾���|JK��'��ND��:�ţ�����ߢd�>��TE�ö#��Vq��y��2��.hj�[���K�e�����©@K(x��%~�����S��h�� A�,��:�����ʃr�y-!alE�Oa�2��Z/�<!B�,��=�,y_Ex�sM��8��l��`�/:`�M�AAs��n?�����.��t#I��y��\���3)��m{�R}��-3�����V��nc��Zm�@�Y�O���;N��צ�3�e�6g����i���&�_�{��H�Q���(Y�岄��R!�T�u#�ȿ�[�<)I���\�
�/GH���B4�138���T.��Kp/�3�Q�i�|az�dpN}�φ�v��Q�����WL[��ɐ�0�����g��0�D�91��zJբ���S��/Ά�QUТ&�/�)۔g�p�K�Y��?�&����w	JuA�45��ZbJt��;�[�/XԨ�u�'[�����.T�EM�6��U��5E��%�-��9�����&��~�EH��rv���9�|2��nܓ2��b��Stu��Vt*d?���)��Fς$��X�^x��3R�IJ�4�)E��V�!�9�e��U�䷍����<9c
E��զ����7����r�[�&������1�5�v��lYL��E�f��'��~�ꁦo�9Z���b-�MY�DߨC�8���[4zL���v2h+
�^ڤ<o<�x2p	�s�i�f���.���,̂U0�t�	���!�`sߊ+���9z%h����vq�R\�蒿���{��K���V�o�2(������S��ō1{Y��6�� �>��,s��{���d��A{}�9.��(-��9�o͏"��1�\�$�2H�2d�-�����{>YVJ�˸ő�&�$�|��z�	w��ϩ�r���L�
O��v�����ji ˼]a�����4�ӦD�A����o�p)�H���Sx��%qY�b+�E����ZQ�R�:U)�@*K�I��<��d*�<�!y˱����_��G)��Ռ(����t�ef������!���}���׌���=��:����z�&fC�R/���\
�9�(ť^XW�~�'��x��q���^�V�Z\9��g�r�*�P��ΐZ� 18'��$�/�ld%�U�[Vv��}s�<6�jw���Hg��V3��w~;���e���$B�����+�;'�d�p�*^�2�4 <u��~&O�*$�%Ys �(�PP�7Sz���8X:��]t ��B,S�C�FEcm�O���~�V�UiP�¼���Z4��e�����=]!u����-fA����Q��';�f�r�萠m��d4D��!���?�q���94OǨ�Zu�����6�
��o��ɚ�v�-x"��Υg��/���I�M-JdeZ��ɒXmq44sS%�m03x�(�`���%�ǽY�cg./���}i��p�RE�n��0�ӌ�Aw�JbǛ���I���E����o .x���q�z\@�mPL����T�rf��Av��;
�����F��0܈�c8 ��.�0��Se�$g�����@LAr� ��|�cR�$�6#�%�������/F�wX���nO��kSG`��z?g���,�MvQ(�Y�����uݬ�/g�e��}�a��Ԧ���}gM=\��ߕm��ȄO+��V��?�$K��7p0@���	!�K꿪������o޻@I� ����7ѭ�9+P�v˹��KW��L����V�A���f����+K;�&�F��a�/p���ђ��[I�ef� ������/N��� ~$���n��6O2XBg������oe(5.9���f{��?xC*�ġK���@I�4���'o2���"��n�g�_���d9ժ��b�x%տf&�dnb��b9PS��Y�}d��co�tp,�PX��||hJi�#�^�����!W'�v�����R��V���E�TY���0`��ۆ{����)���;�s��� �C�;B�~t��"L�@�PP����ݥ\�sW��? >�/�.��ck��z�RW���W�|��������˲��"WY��܀��y)�V�'@�i��.�l�a焒6/�Sm+��!����"��	5?$h2��7����� �K���
U0.q���w�9���: �� ���9Y������9��PS�G��7ʓ��o겟(��jTS/g��������� i����2ʾ�sf�<��3@���nށ�x�G��2���N��z�AǨ�b������< ni���)b���*��Z�gQ�,,[�������Zh�a�,|>*೺��_5�I����(��(A����~�R0kW7v�*���m��G�$hl��d�w�G'�"�p4��O1��ET%�v�k0&Ȍ���B��/��6�O�B�a��~�uW��fus��ν:Rti�S�IN�!�H�B[H-Z�LH�8J�cK�˃r.W|H /c�Z�F|�+Z����1�!G?�.���P�<�Ǆ��������W�_���[}��
aس����EM�+�����F�Y����|tl/¼(��yYG+������u�1;�f�isdx��I�%��,���ٿ�)�B~�Ƹ�0�Z�-��fk]Q�]�O�L�[�7����/��p.aϻ>`֓{�Ћ�{�֓�q�����g�O6 �$y������@�^��C����g�yH"6��!ςy *T�~Ni̐6�o�j�V�f�l�����¦�����p����oay���+������q�K{���G�����T���H����S�� ��V���7�G�y���-٤s����Z��#=��M�R��g������}�����m�3ӱr�<�C�+*v�	�j��Vz֋o�[�g�T>~�QˁU�)|��>��WLK%bl-���������V�������;��H��'�����P���@��վ��UG?��R+�Fm«��
�~�
�ؿ���1x�2	` PŬ�.�'�������ձ�6W��� ����<��'����C���j)Q�n�l��L���I2�����H8��\5]�F"��nqp75N/����p��=q+�Aݗ�b���:�f�]�*�NDY�~��߭|�(�ҡ{[./��������]o|��z$�7�^�d��]'�>�����[�:�i@Y�<]a�}�q��h<J�/�~x'"�$.pC���v/j����V1�B%�`[1���g���q����[Wu11W�-mB���}eЈ���l�E�q���������*�x�ˠ�F�Ծ��<�v�Y8;![Ύ����,�BT5����"�e`#��E�&#����
�DF������&�&5��D!�ft�j�Ʉ��ی95yJqLF��_�q�wC�D�%�`�e�<���A �e@�wפ��4B���f�G�I̛`�*ߜ3��.k!��^�"c;S-�y&[����7�nf�m�#�y]����bӮ�9��t�Z�9���i���(�b�Kfk�Z٪��)�KRD�8�f�u MK�_�Tr��}
WiL�i6��5Ͻ��r-��7aJ��&'��{���؍��&a�ƺ�����l�n���+ŭ`�d���TJQ����]pJyӰ�S�hM�h���=]T��h�4
ùѨ�p�Xj�4��8��!(�e1�0��X�^i�t��l��X��������(b��_Z�Z��;����u�7o#0k���]L����A*�*[����R��Z���W��C��ISf�<_qWm�98b;4Cq�{p��<�~���a��g.D0��))K)ŷ��ãni�<�y�d�����$׳W{������̈��Gx�%9HjMm��~��m��4�M<#L�G ��%�*dy{���:v�l���g*�L�������5[Zo=sJz�3�X�/����7sD.sp�a)�:%����tm��5�+��2@�_�x���F��$r;\�(X����A�A@��^�] !	�'��}j��^�>r�l�A�[W�� �G�i�%d?`�u�ApR�g��[/�J�7Y!�r���Ǣ���\Ln�ɪU��%Ȏ�Zu$0�M�J���p'f������8䌞�>u�9s�G#2�~��ƌ?p��f�����90��W�����{����y=��v�#iH��g��,�9�l���@�Cv�����w��_�V;�ȔE�:�Q{�f�ɓ����4/oj�YZ��FB�����`�4%}�+����ag�\��r����_F�O^@m^�>)�|��#��A��HQ�۬[�4R��Ԋ�1/2��=1W/�b�=������GW����	��_�1��ߺ�[�5>s)�x�<�~H3�⍜�Tg@:,{�T&��>q:�H��O�&|�N�⺹�G��cظ�x�=̳tBw&��lPR,N���:g���S�;1H�ą7��w�h{�w���Rpt�d ���}?.���˙><��e�S�S��Y�ADz�k�Z�+4-���yEK�W��#���#49�������g��5<cҽ�S�m�X?�fU��%���[�� �>���}�󘗴Y��c6[_l̪3��Wf�zbJ��g(��9Ō�ɑ���3/-�A0��4���U����}�)R�є��A�!��7�����S��9Ա����z�%�gCKMjL'�Ͱ���:�;T�&�}/����2C�i���U4F�'s��s��r�J��zvd&�/rB.�_�u�v��أ-��ǯ��7父ȴ�v�(�B��s�����P�U��ѵ�p�)��h=
��g;���ΐdW����΍|��;
EM�3�'ɿ\	b�?a��[�~����&� ��SOă|�0��7��3s������g�P�6o��y�Ow\�z�?!E���H�'}[MC�g����c�������y�z���H")�r��|�0P��O�?5�<��oi��"�|a�X p^<�z\��г����u���F'L;iȣ��E��1����`��"����'Ŏ�k�O���-���UE���:՜~P�a*��L�~��d��
�y5'4K���ּ�~�<P����"ͬK��ui�,����tn��x������5��I��,{�0����Pn���&!}O� ״��Xl3���W3[����^� 
1�0g�L
p=����)e`xq��L����������)ס�QHѦw�¯�I۴u8I��:�I0���=�����5D<ړ�9�J�U��¼X�v��hG�������	7 ��Μ..#E�k���M�vyi#i4���YA���"�aP:�̶��)���(]���\��gt���:M����.%Q^���Y��eJUx4HL��E6�"aC�
�re�������������h���N����c��?Ԃ�Wp�e2�MaǾ��� �S琤�D���YH~���m=:�u>6��]��&�����F-����M�v�r�R%�Zr���&
��F:�e;�K�x�{f����.�e�l*
F����N��]���$zCx�Bsq=��\[4]��^�jF�!�vpS8s��f���d!��".$�;J���vh���^�q!�u�Ƚ�p�')e�,� Oks�	���9��<�܄�M�no_�L��3�q͌�7�e�љ���GR�r��:�!����a�	IߋJ����������n��6|�>��^�U7���M���{=� �L~+�ͩ�i�K�ߞ#VJ�&��/E^�6eպ5�*>����}�e��O���Nk���a>D�oE2y�"u�<�	�=�� ,�e|��o�%�ܛȜ�a�c�k��[Wב����m�p:�J�ˣ���1��L�u�{�w9����MSL3U�X�Q�4�$�I�B����B��Z%%�3�%5;}ɒ���&1�)5�����3����v��@�&�fW���aX�+Z�x�o���eE�98ۧ���*�V�i�W����R�3ٶ6X��姻5 ����DWշ��2S�{��=Urak܋����4g�.g��ZIjb���T��1��a@�|����u�th�E��_z���G(����Y3����'0w./ȟ����}�SH.�X2���]���;��7d�ޣ+���64oF���7.�#i�x�ЇD��*���1�K&F�<����ҫ����'�0r���ޠ���RX�����>[�#)ʏ�0�UhR�y�����Ș0\�!'WJ��D0�Z�6~�_�����y�$�|D5l���)��E��,G( �Am
�r?�Ql"�~�Ǭ|a����n?-��*c��9���X��4�
R��e<������ʭ3��B[��Q+�|�|��5B/�[��\`N�Ӭ9b���a����mH����򚹢�F�"��ڲy��[D�W~��x��ᕸ�R��T>�}SU�0��R࿆;�e���X/�R������V7Τ��J`:\�a�(�U��(����tL7���%��@F�����H�����U�P�0��ᣟ���}{U��C��BA����q�Y�I�K
�,"y����ۧ���5��b��c���lg�{M�I��9��_�gN�_�<���m ��W���BS
���<f�@X������<�'�%%<��Wx1� 	�QppU�8l���.�uͿ�)I��p�o�a����P�qc�1фj�*�d�.�� ����ߥ���	�,z�o����p����SF�u��rD%��[B��?��h{���F�>�4�\|K�̿��052f���[O��K ӊ�ĵ���u�Ŏ�jwg����.&���Z˛�b�q�qV�
��EN$st��ļ�X/�_�R�S�8���Z�DP��q'���h�� 7
ؤ:SЪ�X;WH���?� "�����T��/���m{Z�V���F��@�؟)��H!�.ʽCa�j��O�j���,�5�)��2���*�Dغ��҇�*�{�(��[
��x�>,�5�M;8��Q���Ā�h�7��H8���S&A�B��P �
"�*����T��X���?)���o#л�e<���+ ��x2���<G��\�L����4AoBZHG��+� ��Δ�]Q竫�����>�y.�L*������+��Y��!����`EX�XX,בjn��r��Ĝ=!�Y�^�{!�����Z�C%�����%X�x���ظVd(��!l>�<Ra|�N�j�x"ںb!*9'��a+{�WA��5�U{�!�~�C� 3���1����SW-�t�C��Q���ƪ]�ơ�%j� ��[�1�:3�m�ug4��>�. |�jD��;���?F���pБ�w\ԳeF�NO�h�oל��?.��1y���%�u�������׭=�cV��"��Y����2�u�ab�o�Ԃ��G���5�]���o�gzg����-�LE�:k*���m�	���:D�� zX�2(F�����R���d�YXؔ�]+!��F}���nʹe��8^Vϝ������ā�~K�������F1#��W���>:ؽA�9ۚp����cTS�FUJb����'�^݂�.�<׭��X倚?��0�H��MFU��Q��.��Z��ku���-�74�OHS�a�U5�DDz�.(�j$����u�^���V,@Z/��0��_ʜ`�PC)��d��يrk�[<��Mt�-1uj?���t%џR�)RQ�oü_<Z���@��p�e�����ҿ�pP�S�Գ���|��!pT�Z�q"�,�pR�q�dK8_@z��+,H�)�4������YL��k%����k�PE6;7r�o��;'o�8��TP�;��tܧ{Cisg;���Yp��H�8>	� .%'�{�*;��4kv���ʧKa�dgJ~�ӴZ��)H��dl�+����.�M1�?��76���2�=W���<��c;���U��EݣCꭚD& `�����y����i�< Zy4g>�Ј��d��67.�������.�l���w%~�#�<�Bw���I�.5��r�&�Kybш�r��_������"ߋo�CĀCh�cI�%7�����T
xql�ހ����W����?���yv�V]�x�M��ā(�+kK�ax�@qVPq���n��d�F���A���X�G�遆)%��X�8����5�jL���m�����-�G��&�,<U��ǵ�vI��bZ��'�c���"���m��R��h���[�ba���I���6U��nR�^ߘ�Ī�*�}o��|�F��Z4WF:3�w똨|3#�I�5-%:K���p�V���
8�I�5�Z�/��]�H� O�ߔ���"I/�t���9;��t3�O����F������jí��@��f�eI����4r�O&l�A�e��H0�BȧJ�T�+R3�A�%Ӿ ڍ*x�Y��ʓ���k/��7U���|�3W�ζ�wف4�3��Oi�>L�L7�K��K���TP߈����M�ޝ露�E�R&�'�Gv��P�n�G08Vڝl��~P�0���Qg� �E�.�v,�En���������P�U���m.�Χ�\�� ���HG�r��ge�Xpu[ΡHU�=#�Kp�EL�z�H8T��RW�'��ηm(�p�*�<���Q3��'n@�l��瀥��(��wh�TH��.��Hb"_��}�p�X��[p���o)1s�o�G�%�s�������e�Z�̱�>��b�ӵ ��Y�L>q�"��di]͉(�{��Y��4�*��$]���K@5������OT��P;.=������FC9��?��)����Š�3���^y��Ҕ�{�0�3.�#g�h�s����d����l��������D��Ş[;SA)���i����G&�I=&�[P���L�D|��c�`mj�C��5�C�������	��[�JG)�F�"���3��Yhs�9	���f���d����N�܄�:I[\V�j �Q4�h����]��#'(v���=�5�KM^:sE��P��v�.��[m�"�[���ŎQ��Кk�P�(5B	
���i�M���<T���+��&�&����u�? !� b����˒�*v�;������v�I��Lk�\�-�F�S����Oa�w{� "u6	���cl�k�\��v�cȎӅ:�*��(-7:L���5�[�Z<R,YY�`7��C�b�<����.ց3~(̟~���Yp_�K����Ż8�I������'	�Rc��v,Ð��q
<7��I����&���ď���~5>�N[������D��A�/3�8\������&s�FůD���~V����U[Ę�eE{��k*FS�5H�W&��� ���7�`�� ��"7�e^\x�?��F��^k��w��e�J�;�[���vǎQZ�`g�c������P�=nxO&]wg\�Y�,�����X<*�85
~?m[e}�_c �U���+����ľ�Cη�5*�J�+5�7K��5qO��lm#�!����]���Պ �� j�(�����,?�����锵�j++���40��{�*�H�r��T"7Xc����m$Kܽ����1�-27ř~Sv�\<yu?Ze�F���ų��qLsEU�/腊*�����Ay�]�6���`�H<XG��<Zeq���p�mO���d_U�P��;.��`����Q&#.��z߱�A/5;_D��Y��5�L�H��X�hҠFN�8�]�!P�sL�m�d�oyw�J�"h�B,-����V��-���M6���2i }'a&us#�
w���W0�Ǡ�nH�4+V61�#"��C��e�BB���.'��en��ޜ��tȢcx�1(�RGaF�����L�O�����A㮸s���U�"|�xuj�Bhh������J�>MՓ�4��{�R(�d��slEm&kT��@�IJ�R��?z�l1O|��ѳr�(�XI�®pR{V���p(
^�2�o�-z�ݺ��}��f��C�D��7ۭ�Rݮ^����u	�p�O�جݯ��Dt��m�~���,o���S)�)_E7�)����ͣo@�ۛ���EpWud������U� ���ы��wo�<e�0�-#v����4#PPu�	���qk�pTJX�o^�UqB��E�d�󟷵8��^8[h��&�#�6T��_�H�"���!r����M�nwJ}�� t{�xMI^���wI�/�S��5 /��I9աfH��B�C{�G!��p�r$UY���i�(�q�moL�$�K��;�A]��2dٕ���8��59®c:Pt�k�u'd�L�U�Tx	�>f���Z�߱Ҳ��V��{_���귐6�xм��n�w�4t$�s;��.�NR�vk������F�K��c�731bH�<='h���C���i/�����q���Yy�b[����]��d�4��]N��$��g5�R����[3"-P����9�e�����IJ���f�Km�_O�P;�M��-D��.=��$f�<��F �H�V�zd�9�������f�jxz�	��6eG�~�-�?��Bʑ������� b�r��&by�)�7�x���x�s^Sh9;�^�!��a��f=`����I,��gw�)g(��c�����>Z���&	��Ĕ�0�,�i�����I�����I�Mv�#ܭ��!Y�i�
m���?��)�K)��S
+��aX�wQb1 ����ҽ$�o.�5Mz���8-)a��LJ�G�5D`m�x�@�ΟΫ.ҷc��"�Bs	���O�W�̪�?$]��/ x�L�&���2�#�~�n�� j�����q�6��h���O��%�p�Ռ��
a��!b�A}�X`��ȃU�<d�_�W����+��],���|�S1�j͍�n!�ƫ*Raq��pC����8sZf��k�,OwĴjfՙ�G��eD�ض���m\�p���pZ�=�A�*�L!�s��f�:;5̎�t�}Y)w��~�r�M~n��b�*i�e8��5@BW[�z=�����DO-n��B ���+F.>�ͨ����"Cx����	�^.\Qf��e��Rv�ǛW��ʟ*�ϣ��<*/cǄ
���f�0+@����2��1���kE��ui�%ޓ5��"!��9z:Ȋ����30`���I��"I��W�JJ�Ђhk��^܀˶��En�Ì���\/�5������ys<����DL8�1��
��_���,wܰP��̊�x��z�W�\VH [�:�o=�1���^��y��3��kă�m<
���;uFɽm�ډ�ر��y���d;�y��_�γ#碬�"����]��e-m���� �� ����R���?�(���;���0����;���[/��_`Pm���=$�E��%K�%����V��v�pT��:JKl����nz���.�'��Xq��:Fa����K�{��B/��0p
I	Ǜ�햠��M}�E�.��C�U��6'��� mرx]Wt K�B�-z�[���q˥���V�O���>lh��
Ȱ������m�[��pJf�.�܈�90�7h��j8 kyA����)0rG;$฀�S�;��%;��;u��Q�O�zR:��@��I)�����K��-��|2��޸%�ܰQ�W���90_�M�d�{C�L��N����ǹ���9���5l����ٶ�Ə�W(��p�O}AΖ�(�6g�;>dMir���䡊�˺R��|xy`��+L���1ZP9�>���A�E�83V^TH�5sSA�b��2�է��\��=?����k��8u���r�����{�NO���ꢝ8 F�u���Io�/��\?b�[��ȼ�rkwE����-Є��q$��0`�/�4`�&�q�gʿn�����T��_�֢�s?��[+K��
9���b��������=� ���Be�)��!����T�c�$�A�ʙ�$����c����;DMOdT$׊-^���ǆ�$�$��iz���B�����:w�PQ�gx�����E����4����nt%I��se�N!�7�5����PT���j��i�v	w�Q�Z�L���2���pmt׎ �X��(f�b�."K��i�x��������?iS��RQ�Oe~�:���n��2�X#ڴڽ��J�,�c���ͻ�K�:�� ��H:�� 3�TL��`�?o�ć=�� �w���n�=��,t�^}�&Dm����m�+�qY'�p���y���	��و��;g%E����g��:'�H�f[��=�����e{F3��^H�)}IZ���+;���&ǈ��?j�p�?_E�Y$ �_��W�������*��'$������ɲdд��9�E��)�Fs#��!18+dC!.��T���o�~�[������� ͻw��Q<<��vx�MC�Q����}�o�*��Ō�\i��ʤ��Vg<�J3H�½�:�W��)b7�{t��w�r-���:�3T��'S���6L��^�	��QD#�Ԫp�ƅ�T]�Y�1�q�宭yim�a��&�gנX�x��^L�:�ßH!g���<+�t�cm׎<��ǉ�7e��os�o�1�ټ��W�[o����	�0�Ý��
킺["8�	���x�3��E�lȔQ����9̀E��e��-]%V�2����H1q�C��[4w-��&*���W�zog��P
J�y5��d��V�}�,|ƹmѹG�L�Y�ok��q3�-�U��x>��4�Hc����<�� ��F��V�XS�1H��L,f#H�����D�y�w�ǳ�͟[��R��C�]��_�Y7�q����0aG�[d��R�ɀ�����ʌ�A�p���ԝ3�X�-:�������d��py���t0�"��R�>�}�-����~X�,i|�=�A�/�&�ʸ��pS��9�Ҳ�>a馋�lѦ�#�4�z��s�R�Ԙ�F>?�`����w�,����6�Pg�q��Y�~�3(���x�&��1�X!c�r�ӆ9���yZagQ�|��*9e�|]6��8�]��{X�W�;@ ����'��[�97������@^t�p�ԉ���ZF����/`�#[،��`��{n�ee��#��#��Ϫ���L�R 6���G���,}����T����>��B��[N%��T)��k���k��)|��^����sy�
.�:rH,~� Yݺ�����O���*{z M�ktƸ�d� R.�&��t�E*Tp�����F�ހ�M�.�Ϯ����Q{�	O.�'E��G����3��׽�fu+�4�y�}��MK���v��F�zc8}�\#�ҡ�t�s��Q��q��j��5��6�����(������|5nH*��VQO�qL.3D�V;@�CӔ9�Y I����\�W ���h�BF���ݕ���+��|ɰ�L�ڜS�u`
$.�v�g�a\�M��@t$n}�bXa�.sࣕZ�v�YP)��_���yF\ɝ�Q�N"Ta,<��wK�t������Զ"��(\���MM�k�Q�S\!@E�׹��ʧ����@6g�0�Q�q�"$6��W��l��iaQ;]y%���o�ý��V@��&j�<]|�,���E�ѕ�,B_�}o/�.2����W_�.�@u�MЊۯp���h�����*�)ʫ�f��S��ìk��=C#�/�U��o�P9%H���N�A�
��2�[��a�H"���l��E�qp�j��#H�㈦8$9h�ƿ`7E�t�>t5F?�#]�z�a�&�c����a��G�X�S������Ld w���f!z�]�\���Ψ���bcƾp�d�_����^�|��Q��e����4z-^ZZC�ќp��̱��Յ�[%0��B��qt����L�A���]���&�c��e0ȓ��OH0z���/��m�Y�hO��dK��:V�at qr뱬5/��?aCӅ}T;'/~fStiA:ȵ����Q�7*R�e��s�s�� ��y���~r�X_�f����2�l(�A���Y�Ñ�_�9E��ߡ_/}Z��� ��dF���$h�WL�<�x�@W�b�a�H�\��7}e qS���p�2q6l֘��:F�1S_�d>9
�Z�������	�N��+PxrቡD���nز���V%��H��W����S��ឳ�+��x���Rq����v���Xg1�Of�u<�d�D2J�+dE2�x�|�W٦���ѥ�4m���8�RR������gK ���b�p����~�]��a�S�ܭ��a}쾙E.�������=�D��T�c�Q/��<9�QĠ�Qͺ���4|��U*_��eu�őY�>sʧc��d�BݶCD�>u1��^;�g�!�'o%�;�&�Z�q߿�p��r�������ŊF��f�A�>��S�B��0xh��pr.�[��+s3�#Yt�.�w}�C\�fJ�����]н�KQ��Af'��e�N2�jxqؙ�cq��E���/S). v���G��w�h[�H�j ^J,��v�YӐ�$�Cu��{9��mH���"J{*�I�;Y �q�x�9"��ငE��4(��WQ�o�2,d�W�B۷�p�VT��`I*J�1Є��6�4��ߩ��y�/�H��K�yfY�5O���w˖�B�c���D*J`;�g����U�%����:l�	dq�;W�ty���f��	j~d��o�ɶT8R�'1�ž:�GS�e�%f��S��+�*�~���m��K�U����jAn�����r�����}����6�r�!�0�[7�FU�!+LV~1r,\�t@��6�}F?�~4#z�E<I����P�����q�1�q��;�e�e�����%�� ��L��H�����#�U�۲7�-R1۫˱�{�6w���ũ��jEІ��|�L���_���k��BtR᳅Ŵ�h!�6��В���Р���E�Zxgu��&�~3�;�ԍ����G��}��Ȝ�q����u�� ��|�S�l�=��t\�
Ȧ������95�o��_8�����;����[�sL*c�s*����oc�1޳��SU1�I�΀�:�����HR�Ҹ7a�\.��8
�%�;��V
�Dd5*��.ͤl�)B�QD�����`ޛ"�Û��T�9�2�{J\&�Ð_�}��Z]~}�bJ��<�}���O�}�f����4w{j�q3\)I �:�6<j�9ĶbkW��]�|�S��^��4<�I�s��.NGm�Y�r�%�/��������*�*�+r������;QZ�Yh�6	ϩ�yla=FP��QxLY�G�����7,0/��oE[��ɓv���`Mr�鋔Thy)*3�|&����/l�S`/W㕴z?=�48詝j������k��Ms�Ʉ���m϶�i҅�X���Hm�s�E�i&e�@:��c�^��4�v	�DN�?��4�6i+���sa��-��!������zf{�[~x�Z��I���Æ�}��
 ����i����H?�~(��+���{ٙ�-#�ߝHn�	����L�7�4I��%Y#���X����b���Cr��
�l�y>6ʘ6Z"t(-�aW��RK���?�	|��W�9�]��;��l߆#S�5���3LzKo�� ӗ4��M���X�j�����y��R}� �|���Z�Ӣ����uW"��s)𓉸�>�e�N�-zU^3����5��g0�(�?�� �BpTZ��`��H���U񬥙D��,$T_�
�8�kw �aڐ���O%�6�GPI`��^��XY�ҿ�'`'�x�$N~kl&'��\8 ��A�ف����N��v��nM��R�U�.������d�L��j�"{�L!2����{qn�X�X�*�M��*'�;�r��cF����aqU�<<�]����F�Q������0�N#�7Q��<�~���S)k��`�B��?�j���L%�[W���W9#v�H`���h����$��i���д�����=B�;(���H��������$�OU�=@�ZE�d���N<�w�f<��?������7�ɑ�C���X5Q���V�3��phef9yRE��������!�s�RJ[}7ϰ�m0���8|�c��3��ޝ��-���"�2��b�{�rxr/,L��l���gF���`c�^�����=	7t�H�w��+?�. ����P"<<��
J�F�>����Qr�=�XE	�X����iEXS�jlD�"6x	3��?�Q���d�!��',~��KO�-a�̈��Q~�*z"�dqቝE����C��>�U���fMKF�ri̟2�Q��1e2��Ħo$ʗ�EZD��"��&ۗo��?5��Y}�&����ㄟ+j�R4��ں�%aj�p�ᷟ��yZͻ�M�)P���7���Y���R��K��ҽ�p���Xi�z��C�������or��M��!�Q5�5~>�9���ݏԍ��A���8���l�Y2"8L��eK��N!~t
3;�KTC�U�of��քMN�l�
g]�"4}_z��t��Jg#3aIS�h AyBdg���7l)��;�$[|� B���=s�W���^9��K�ƒ�¼�ۥ&Me�T���I�_�d}���k��D=Y�#�1�˥��686	��TI���������N��p���q�ɽ�:i����e��UKu���Ƶ���)��hÄx�5�%^3=����||i�!�k�,?�Y3n84=!5G�k����x��{)*F��Dcb��U���g���j_+]9d0�9�CB9A1���ڶ�8Y�H2y5�h ]@�ZI����@@@�}m@*���v����稧�����E{❎��;:���w�8ʨ����lZ��&f�2F�uj	^є�;��x��Z6�ڕOn<�`����2=��$4�}1�b�����Z���P�������iQ+�����`�6��1!t�1m��髽�:A�T��=�S��$ ���6\�g��ùO�m1��z�	���@q�e��MK�KG�Ԥ�+G�]�=����bt���4׈c�q�)��'���x�/<U��k]������~k�a�񭼝�/�jtp�+O����_��C���
��>��-�D&˧���(X������#�j��S�s;]k��뼦h/�ܴde~u����!e�wPu��-$�j{~�=�o���)p'14g��Yf)\u��=OU�b�&��u���%/I���ٵ���;z��޾��s�i�wQNŰ/���c�ւ[���2�^ޤ�b�J3CE���:�/{�h�@�C�LP�����SA,-SU��E���Nq�E�s<򯳢U���J��	�>N!\����t�]U	����9gM�V�[ny�`�`<��֛bf��E�1B�_�����jo V�C:Vܡ��*d��G��"��}Y�s��u���q%�! �P�5�7��s�f����su�1��"F>���S�������Fs1���1�{!馜N��++��	�ָ�/�!Ѕ���:��A
� m�򦰵Cb4�>�� S����Ѥef�}�g �s��7�?�ӄ����#��-+]lՄ:t��b�*+.3��q.�� b�*ZڍN��k$�t��g`�+�����m�<���'L5�ӬH}
���+��������)�x! ���O�`µ�n8z���������󲱡�N��h6��Ǽ�Q�\	<9W������C���4���� z��a9ew6�mT���));�d��/|�0yU�������4���c� �� �tZ�f1����t-Y��+���L��!e��;�?�4c�w�h�;�T��n�&�ϭ�?1�-�_�� �S���N�Ʊ���տ^�:>0Hx� �o��JpVgK�{�>g��`�)N�����K �S��x�
����`�C:�;��oX9�0�t��J<��;0���ئ'���!FaH�C�x���ʋ E��R��dh2$�I��Kl�G�ld5�5kH��o����S����I���h�r�v�T���������lIb�y�O�#�gs�G�L;�
8��^�k��A�]�!������Ps��ƾ�lZc�C)���+	F'��y\�v�o�8�IP�֬w^Hn�͖=����΋�!�=���������cf3����5��z�[(��?+�:�~u� ����ԕw�E�%����� 9�b-~8���t��'|	@>8�h���6:S�T���t/⍆A¹�l|Fxk�NS1cL�<��s7�EX��8�k�x5<�w��r�s�I@�y� ԋ���;�?��A�\[j���&~y	� 2�H�9Vs6=znE�q�o(�p�fx�_��x3��(��K@q���ɑ>�,t1R$����񷘱� �l�
�m��iD�-3�9pt��L�-��:3��ϸ�>��E��$AD�@j4|�zn�B��]�q��hP�M�,��k�적\������F�UA!�#|t)�9eE��	8�O'�R�O�	��U������:5؟:��e��9R�6�P���+m�lM�F8�u~ю֒9���N&I<7R�p���?^�(cr�!E�__f2�	�xz0*�7u�v�8��5���l��M��v8��W�P�ŉ=`�Dp^����Jh��X�%�gXHd��JE�x�f"�5���4#����ޥ���Xﰾ���e���;޸��6A=��%!yD$Zu�;���w������������b#?tr���'��	O3�r'7j7������*�%	���椢�]� ����gEFWN�ﶗ����O~�;����"�٪8�Z\�d����NAcݏ �K���9D���������mK�Ȑ���8��Yߊ�j���[��pm���2�2���H���,=s�sf�����J�iW~>Qg�P�f����f��R1ֳ~�*�q5'�)�U���9'�u(Ѻ#S���H��4H�Q��
� ���ZR�Niz8�Z��fޚmj���pm�v��s1zj��Om���7N�s1&���V�GS�:n�@�S=8�r٬�����Ύ���Pֱdx�^g*c�7嘡,�P�'o{��˴�l$�Eӕ-�����A"�O�ЈiW�k��WRbZݟo�����9��ؤ*�iW�2<�D �ފB�h`
[��Y�_\��.^XϘ,���+v�2&G��6(9�p$�u��Ͻ��͜o��-����da�ir+$[��|ȁ|6i-�"u}Q�(��8Q|ztm9Ȼ'�?�3O��a��N�n�ɲ�p�[̒ �j��8ѱ#�nz��������-���8c/AUη-��
�X�/_y��ݨ���5L*3�)z����L�n�U�b:�]���u���b������|B֘"bψN#342�eۼ�nG����B�{P
��.��xgG,�N��1�c��m1�[Ot�
��
w�-=:5}����q���ͤ��i/]�ݎy�y^Z�'P�b�֭�`�R�������i�?1�񠲭Z�$�|9J
]�A�&:�5�d�g���8�(/7�(�͛K
�DT[^����l���
ƎB�R�������,M�X�<!�I�'��y������������6�	�3*.F�O!�E�8�7"��Vu�B��J9�9�fm�B��1��g���9�7S��Ǥ�8IC��!�t
`/�H�NjhwvS���2s��M�S�����˒g������q߲��DF��{���,�ո<K�)D�w��'��֤^����`�����l9AM�o��Z���²�"�ʻ�0��ϐ�V�ښ��K�5\�:��K1�[p���z�h&�j��njYk�j��|�k�M� �$��W8n��4�>`	�{B��#�����<FmhB�8@'��E�"e_"����O���M��Sx+�G�;>F�������>�V-}���l�iX���>�y�"�$�~(�c��O�[���"z1��A^���~3m��:�"�$�6d��`�����.����-3�>2�����_�	3�"�ޣ�Ml=ԏ(,s0&���KC��$|#�J���'�Tf��◿P���3��]��Jj�^R6���Q��{'&1�>��:^�a�dֲc[�ژ� �5 <�&����Qe��Z����-'6+p�;~S���M# ���բ?m7J����5��m�"�a�R�lI{!e<��؟T6�~��<�{�¨H��DL��d����Qt�3�Z���E��`q4�i�}5���.V�<���L@��gf�C �B�+�j�AI�� GK@M$��gg��f���-H�\�t&�
z��E+L�r =F��@4U��N�g��h�E�g�4/\j0�:>{�2��4ԕF��x�&�DT�ާs!�$)V�#i6;��Ө���Iek`�`Ps���.ߟ��g����)8��agp�ܭ�޺�E��[e�!�Y� ���u�xZY"�Ӣ�����61�Thi�mǄNu����(�R�A86���V�&��l��+��8�E�~��!I֜]eK��E�f�����F����:@��B����<�g�/5}�kψ�/Wنʈ��r�2`��~0���� �Ӛ+� �{ٻ]�� ��P��!����?穲�ϒ��n˕e
f3��q��{�	�-��ҵ�ԛǩ`L��c�� W�4��_��1.}*2c�<Vȑ��#��rw�ݍ�(���H�W2���z�F�ߚ浐m3$s�6v��%,��;xIvb[aڙ0i�g�M:��[=G�[	��
}_2!.���"�W�bF�I�E�l�)�w�fD8߀Y�\:��kD��i�a7�))�/�3xD+~�_�i�� ��7�Oi)�]�T*4d��@ִK��@+��?'r�Q]�2pr�#?�P�گ��X��&+u���V����,/gY��u,Z1=�a�k��w`�''T@O��}�}6�*�^>��H��6�ʓ�F��:���풥���ᾜ��~�C{�R��l�)�ɦ;�Aw�*[c���4]��}��N���rw��0w�2�a� 5N��m,��6�1p$��9��쀈������>�e�PLHw"!���{�3�K8�v���6�����4��/��rWB%o��ce ���D?�/�hG/�/���8��7`S�g6�i��%i陰�������C�x�Զ��L[���XS1~_�E��R��p�[�͠�_&�Jc}.}o%�Ӯ��M1�Km{C�阷(R�|M�n�H�q������J3��f�N�-��_��!7�U+���S9'SЗ���6f#G��Ϗ<�mpܠ4�.,�7'��f�2�Og�������U.{C}{5�y��eM�C���M)�⧶��#b�v]j3C�������oIS�I��I��o�+Y �<��e�ؾ�(�|��d��UK��)�2�V���;�%��Wн'U/x�b"����я�>0��j�Ԏ��=�i������i��S0��i����}d����+;������#��@��	gv�Z�u}g��qC��G��=Ăc*��)7}( wLvX^R��i��l�k��������]�3�S4hf��U�M��,ت��=t`y�eA;�u����)�&�8�lAoZ�������jLd�Dc*�]I�t�m����W�PL��AL��5E��>�.���k���b<'���H�s�Ks"5nc�m���'0o�ܟ�|��R Fh�6�)�?76�A��?�	�%�2��?�0�q���rDF7�m��.c"
q�`+��*�������n~��!��f�a�,�4������*I����i��OJ�	�<��|B�+{*�7��
�t��rJr�����wh[+��_t���p�b��t?���P�zZ�M+����p^!R��P�`"3�?�C� �z��}`��d��O{���=?bo�����i�"+Y-����N�0rh%!B�[�*G��mǞx���a%>���i�@������n���i����z_�'M����*�4�r���X��탎@
:*�D�5	����uBc��k+�����W��;�)t�7�>�o#�"���gRqZ�#k��mm?��?}� �	&��&�4n`���IG�
}�������[�a6�NXa!�#��Y?F��8uN�[�*$�1��������=qw�6Glr'�˩��7�r�]Q�YM�����e�qh2�t����<<�WP�q�%W]�y�r���Sa|�@%����z��v�<�>e`���t&��s�c�07�?�/$�$�}�]�~>⣁�@!Y�,���Β��M��Y>�6SÔ`�4�p���>`
��G2��o�/�N��}#Y�n:/o��,��,�B�b�� j��[E��4I8���&��/)��'��h�.�9�u��������6�9l�j�4iD�f�X(<e%n��.�LjT�|/lU��Ӱ��Wk��a�͠�lz�3:7��\rs�S����q�z�柧����H;C������%aQ�TtxkH��J>�<���I:$p4h=�罈 &�d��?�O��*��҉��Zv
Q<�����+('T�A�D�~�ao��X$�9A/��w�x�xN��|d6���u���%�Dz{C��G������(�� �.`�o)���
��S�1]���P�o��������(Õ�K�G!�؍�;uI��!G�&_i�Q�ƴ"?3�k�A(a`F)����b/U�����S_�AU�$��f/�|�Г��+��z�ؓH8*����c�o Xƪ�׈�8��9��~{�<�X����?�ረ���M�zE9N����HB;6���ꔽD��E|5K��>o_P��v)�Y�E���s��DW{���	��n�6�R�������#���-4�R�8s��w�).���j0�\�6�S���u*_�a@9M���P�3-�0��J��V%	��eQ=b�����no3��)|�(Zb$o�P��E0�j#Dn/	����1�4�;���Lj�ĈY�!�N 9$�y��I���r�p�]m�6ǃT��K��T���Ύn*��$�l�q� ��^˒Y^A�
I��_�jN�(6���F��d)C�"K8�y�����o8���OU׺)���|�K�z��l�]������)C��rD'�[m�Z�t� Kgo(#�V䞿�H�F���'Zޖʤ� q�����FQ�3��*k�U� �]�����n���կ=���G{|=���{��mC�7U�c�}�AȽR����n�Z	�]8�H��\�0��^?�����"�b!}oE�(a��7�Ņ�$�Ii��Ę�ÆO���;Ҿ�'�l)�a��#�y�#?�yũi��C���N��]�O��Bݯ~���E�VcM����@�\�WܷRu4�k,b��V��n�0��)��{bY6�K��$��T�P��7{8^�RK#vNH�ʗ@r.�Ԛ#���cIwg��F��Ǡ
C�s�7r-���.��x' �q����#�˧Gʁ�P�{�	�.(ڂ?]��/t;Z�
ғ�.Cʂ匱�X��Uf��>ڰ-�^;uy�E\i��'��X���K��l�A��9�CA��԰�R]��U0����#�?揭ِ�m&�a��`}=G@R����Gؠt��x�)�Z�>�������S{OM��+��X<���V�7�>�w*q���	s�@6߿i�� �a�10h�oޑ�u-����r�+e}�)��F�Ad��O79�D���!�ye�@����)��?T,��$�7��H�����3�:��j"7��s���"���}υu<�B���!�&�$�'�^L2�~��Y/�~ ���!�P����������/�U�ҙ��f�e�a�#�����j���*�&ǧ���,�{w���.���`��Z7�
��������9'���);���֣4 ��&��/���>m����QC9F���<���"b�]���%��gp��9F�ꒇcI�-*�u#�x �LY=����}M.l)����z ^'^���r�� �v�j�Ox6��ټd�l��@�N�?�lH0j�|�#�Fw�>�h�a{���Pb4 &�.�y0m��@�o���hOt;��:���/ڸ�M��	g�YU��2*�����ލ�8�& .�H�}�Np`�5�p��2� �U����nד4r)�`:?�S�&'7V�
;�����̟�Q�;��f9\��R}Ne�<
�Zaa|k-D̜�ylAR�*�Q���8�k��;�L�2�S�r���C�;�U� ��^x�^��)o�C�c'�O}j���鲸O1|d��B�Ǌr��L7��v@+9��纗����62���k�v����J�&���8Li�yS��Ʈ���EybZ�	����F��u�L<���xP#x��Њ�sȱ�&��[ռ+P��n�J������	�9T~M����=*��]���C�{>�J�A
��F��XF�.+"+3򃤮ã�A�ء�������z�M�+��ID<לн�驜A�#�G�G�҅�69�U��*��ߌ��o^�>X�ev-]��I��ԕ���Г��:���%9<d2O�[�yf���| P�����T�zO��_��E�&晷�Ȏ
�:�N�a"L��ג����Z^[*G'��+��R�c$�8��>����\ =�	<13H������g����(&W��e!��]��p\>����3�kʻ���/$���ΑR�&�
 <�~�����Awy�-g�13* ��mv���n�Dz{.f֝�b���!b�OT��ʙ�\������*%���q��M�V_v\5�@n�1�0��=�=��Ni��&:#v1�1�!�TݛO���������KP/U�!�z�%�D$����m��MN-#Z�<e_Vw����E+(���(\�͓��4�ˮ�.2d�{����_uz�3��t��*�FLϽ�!��eu�K�qc�����k�;�w��e_�	�o~��Vn8Y��0I`�ca��m���U�x<��8t<���rN�|0��E>�FC�A?�E���(���S�e�L6��'�����9��ʳc\�%����f&B��}h��=��듨K����6����%ϦɅ�Й���E0��ml���[��+�?)XQ�n��N+�9�l�$;:��y�^z{�.��룢�㇪B�� �2��=Y�S����}r.2*7�po)���*!�.�i�^uF�[
���ш㾹)c|��4=�i����H��&6t�lJ�+&ܪ��]m؁S7�Db�2�q(8��t��+P�9IGK�o�n=C�z�}&֥�g�.���W��K-]e�,����i�3
R-:0�-TW� �l�Fu�r�~E�E��d(U%Ė��
������[|��:^��1�G�K�PP�+J�R*��EhLo��A����k���_��v�A�.�wGs���s %��y��9�}TH|R�Ss�����Nx�_��LK��}���r7Z�_bA�y���	@���n-L@��hݏ�ǻ-�f�a_��SD��ԗ�M�_@���L�M��l1U�����]��KksU�R��
��g䢼K[Z��v&/�¯�5�bu�_���/����K���S�:����V�����7�\:ﱋ	�"��5?Nҙ����-]�~����/�Z٬5*\e ��Y�"�1v�Xq�3���S�z�n�˽���ә!����`(��/�q�h�ҿ���6��&�<q{�Ϛ>:�H��D�϶�j��%9Da�K�I;�y~�ӷ�R�_������������;l�,��vz��7ɂ/Z��\g0����f�7�HI�U=�z��v;X���a�Xg=�*���D�h�n�u��q;��1g���\�o��.�9̢U�-��ÎJj��b�m;j�wJм�>k�p�WL������k��f���0�X��3���2����	4+��1_>)��:��'ډ�?���fX��\�Y�EV�<M�ԧ�P��=�C�2W��G�;xJ׋ijJ�ԍ���X�rM\��	�]a��]#�܎
~m��J���D�+�N���0c���Lp�ME@�n*sEZԴ��b��#�wߟ�ȯ9܎�����#����߉U��Uk�h��@�r����;p�z�Ft��RVWk"���-8�q�͚a=e��<�E��73nw�&���d�p�6�H_���ho[T�e����3Y�&�][��<��r�R)�������סr3�Cb[���ԖdnY�����k5r�e:M�Z�}����hq- \m)���n��΀1�=��hŁ��[���:R��p�T��,���*#��;�
\`w��c6�2�'�>��i��?���<��	y.���ێ'�)Nr�rZ�k��-�D{�i��=M\�as�J�Jz�0�e8Й�/�Q�瞁�^��������<�E��j�(�^c4=��.��MC�"|n7ag������܄���(��_ڱ�W�Q�~�j�����gاpz���S�~��V��[����kY�ɽ��r_�ϻݘ��SFCFSذ�,>�eo�*vqWqh.���k�@��1�l�������(�$�9�{����t��Z�)ai���2�ꚱ�\��ۂbIDR��ϙh(�hM�������^��0�Mu*�pFP�t:�7��<�8 $��ȕc��@M��TA&���ud:P�E?a���7*x�iNIj
�-,�f�>����*Dl�@W������J7\ә`�|��B:�|�y\Ofk"� ��Ay+<,��+`}�ި� �R(�˄b�<�!�y���1f62x��C9� 0t�_��A���Mר�Ee�EWw&Iy�O0��	0�}�c��9aC e���'y�|4�R����}1Y�3*�xP�Ԛ�� �Nh�4�	*K�m�*1_�M����$��L�֑t���nt�0lx���l���G6���_�Q���r��9�����򭦙M3Z����B��Ǥf�K�i�8ڀ�kp�������[�p���<G���Rh�2+����o�׏�n�4z�b���k<�(���r^������7���Z3�{-�;���#�1���,��qr	���0kȇ{�������)L!1�<nd���!g���}Wb�b��\���m|�Wq�Z����4A@��cMis�_KC�#�Yc���-�~	�X3� 4"�NT-�p�09W�;Rz<S��,(U�~���Y��p/'e�=~� �Eˇ������v�lF��,k.Br.OJ���I趜�Y��Z�A!�4�\�}cB���bwN9�E\�I뎘d����t�@!_3Ć��ԌB0VG�n�():k�X�������@�Pp�f�=X� �i�x@��/!�Mmc#�C�z����Ջ�H�$�F�g��;��T�{G�luK�'h� �p~���,A+YY�cv 5�|-�V����B`�"I�T��^ǡi�����+��h��I����ͤh��ؿ_e_Ȣ	�K�^�^������
�B��
�'}���?�$����k5/�k��QmSI��zq|R�t�{�`0m,�L���8�H%������&�x���y����J䩦���\��[�ٿqZ���N�9Co����"���x�w8�s��>�wCD�Z��pJ ��0��~�Gn5}������yͳ���i�^CNy�.�p���q�/z���Tbn��x]<��R�g�Ak�r� �+j�i@��@c)���+m�}���e���X0�_�?aBL�B"=[�G����{l5�*({��\��X|��t�S��v����{��=|N69�e}��Q��nX���&����@�y����AcwL�3����N1�y�}T���?���4�l���fD(!?ˤ\x�G�(��M�6����mps��:��2Fz��5���E��\h���x�����}J�:��;�!�"�:ћE����h�"�X\s2��^����xV�S��Q�%�4?*ԥ�gZ�I���H;�$�]��A�r���i�2@@���g6���,�Ss+9-�j�Xן�𨁬C��c���$��-R�"{7��h<���
]5��<��c|w`�`�N�Q^#��{e̖1�e.�ʁj����-�ot��R*潖�^g�c�o�!��[��S��&';��#![،��bV���h�	���/��'�(�!���L��:���~����Ԣiఝ�ģfHn�%�w����7xkP���:�^ـ�S�G���
��6�w��yuQuB��j��W�&�@��Q�}x�[͚���}�:������r�#__���|2e���XM�);E�Ρ�1W�X�cg���o�h-q��'=����^Pн疾F7���mƧ����x�*��`�C��/�~re_�y������ �d�����KrRPB5N��%�nG�\;?I�z1#��'�?7�R��¨~�/��<+7�A"���=T8-uJg��=��٦�N���u��Q�(L�{� 6�Wu����/�X��H�F��W!	�۹.��y��::�O�]o(�Nϫ
b[�m�]v����l�H�R�*�����@7���h��� 2�-�����{�/�өLOI��j���|_(���?T����g&�]���ck f�S�@�T�zy3��^�
���V�k�pN����Q��g�2�?�l���j�,/�(�k��d���/�)���}���=n{�Q�O��L�蹷�^D�R��)<�/�>,6��S��z�
����s=�l@�Z�]���/Qo ȗ��W��v��?���-���c��
��ȴ����E�+��Fu8��&�aa�¸f�����=D��R�)��	�:О���tk_4�)�%��=��X����n�[ĝ��L}#��K�n�D���ѵFm	Z��y��a�����X��	û�mwN,9�J�,`�3�Q;�I��e�57������q��5��ڞ��.�m#�-�������r�2��ye6��	��
+�ܷ�	E5�e(�pG��;�1$\�GW%��M��U�~�=������<`i�Q����iҧ�S̗�:;�� ��V]郍1g&�ʤ�\kE�c����㶏�������rh�:���Fx�,�L��9�r�ǵaW������m�� y�P?S�鸾9h�"�Iڇ��*�W���:_�������|;)<��?�䧜Hx\Pp�	|[��x�0s��=�1�EI��'�xw�O�+/Z,��[o2��DY��� [0M�� ��K.��nµ��h
�.�dG�uQ�ħ�Ykm��mt,$B�5��^2,d��G)���Z_�Q�v���$X���2K�TZ��s��)��Y.{+A>���;`����8����t��c(eJ� l���0�a����Hq�y�'Z�8OJ����>"w�5�UFC�!����"�Е"`�\�>�����󿥄]u7����!b#�|׿���W��'�(PP��K^��q���-�J�=N��%�><����pw� 63�.h�ݫ0��L7+3��m�u��'�4�@�B��Zm���Y�&fSC��K2�F<}�t���m�"'��i������g�v�{�o,��<Eq�˸ѻr�L|��C����&�o�L����/Ą{#Z��(�`}��\�Ԯ�����tr)iչ٥��Ɛi�S&����y���[�'X*�-��)�XiEН�����T�w���긃Ч�S�� L��_�O5�$@T9E���NF�6��O��|�sw���N��,&�������f��6��о��s�v�\d�ut^��>q7F�;�J�lq�xnh`�8�2H���x���`�/:�~��_�Y�[H�pO�X����x��8$����Ps{�hh�&>aj�3�<RKҡ�t9��Na������ V�q�u@��|�ƌ
?M�b`��._
E�0��)�?[���M��������A��H�W����Rp��(�w��k����I-ǉ�u{alb� �b��m#q�b�ݲ<���Ǟ.>�(o�c��պ��`0�E�>�g�jg,�8�EBKI��`��#�]�<#ĖߝQˈ(�S��`Ķ`^>�Q��B��tqZ]#����f�D���Y_���w���x�c��SGxB3�(UA9g�f�N�=�o��y7�F}ϰ���=�{�,L׵`�H���찗���1�Q\H:1h��Nͣ4'��6hX?�UC
O��6�9��~a%��r�H7[O�o>j)�k�W
$�W��OҰ�uU�����7�����a/�%RK�r���]�;+�:���f�<'���T�EW9�(�E�!����a��0�N�i���G��F�P���Ⱥ��Q1��?�ܸ���@TN#�[Ǔ�yů�n��Abz�չ��nT�;�ń^���	��Am�m/kQ{٭�U�/����El����+����d��&��k5W�Ƽ[��q������iG)���y���i��_֮�DT�?��p��kq�/�X�#UT�o�L��E�ۼa����	�����m�h;	���#��c��?�$���b�W�H:,|�����7��Òl0�� &+Q�~Js���׎&�w�E�XEh��lq��4I����-�ib\R�%�z�L̇B1� ��yPr�L-�!ڿ�_Ts2�N�յ�rbd�>a�4�U3w��.1)s��=�o|�խ�x����?VY_6�=h��G�ן^��4��s[��,̏*����ž�N�=>_����vTZ?6y���T���u��������Ĭ�js�1����{8�Yx�����}P`��\>%��7A'xȡ�*�Ѕ����m씌6���q���̖4�G����so�>9�?��z!��YA�d1A&/X��D���<��"ڐ���	�n��m���)�}�	�CJ����dRg�0��GT`����o5�`��O����L�^�Qԃ��c�Izm��:c�g��&p�!u,��1�Ü�����ދ�f3���r��h�̿e�Sc. Y���X@��=�y�" �'�T���_���/w3�kFQ��
��<
�}�D��c���@.��H���׾�{9�ܠ��n��S˵����/��F�G���=�=�-INY}Z�X�b�D��7Bߥ�;ڐǂ��j ����|��g�T*?�IJ0sbִ��m����������J_h�7�9i~m��v�4�S���BH�hR���V���IF���r(�{)��'&O۲����K�߈`��B�lIyJgZص�̐�h�!�Q�O��ru +5�:��4�Hf���"!T��!ʖ4k@8��f���c-���Ʒ����e~�αh��iE�"��T�ɬ���5�(�X���rkw�/^@�l/�� ⵀ��2��	\'���`?� �v_ٮ]�Z��ɗ�9.<ט����G��Ġʩ�|�ӆ�!\��9G�mw���8I��z�� �A���o46z���0����r�	��f֕��-h�}� W��8i }��ml���y���>HQ<8c���LҤO�A�3e�����;D�.�V��i��c
lb:Ih������	���'�@3F�5���p'pϝ�e�%[�{��^ם�_s��" �����v)4!�sQO��Ib���)[m-�L�魹��҃��l���^�3�s|v9��i�5�2�$�C>a���*'�=,h����gu�0��w�L_�"��'n�B[=��7;�eKH̵�;+4�U����緌�yu1o�,!hڰ[�uà�Q��6�˺g�J @�~ Y6���_�%5uŐ���+Y���.�yk-�Wd�pf�k����eD�[-�*�+1���Ved���U��1`"),��w!�����n1��G�"�`���\\//$�G����=� �8HJnw�X�MV,��P	xLMD�F�K~���]���)�H �:��Ē.(�:��'{��1l�+� ��� T9�*s�W������ܫ��#�q||���X��i����{oYΨ�\:������S�zu�k������x��UL��?��5CV���ёu^qoV�5�2W����%�!��C{}���w�t����W�)UA�c\�)�N2�l2���R���
 �|�)���������?��]H5
�WJ�(��Ξު# r^�(ۥz�G�amvwM�o���K���.���C�͠j�A� �Ed� |�ȥ�7#%E\F��_�w}`��-u�S����q�|�z:�jâ�����&i�=_�E��dT-i/�b�9t	&*��Ӟ|!_�u�F%�}}yeY�]�gaܖ� F?�p�~��qO��lc��z����o�7%����u��~�K6<�����F�=���ܳB[��<�cr2<�����_:��-�!�E�W�q���L�";�#;�:���~
�D� ��e1�9����B5e`�O��a�Q1 ���+�����;�cV=��a.�A��'�8������*{*��£q�*"�8p�/�F����>Ϝ�,��|���@��k�l%�aZ�����g����`Xh3b�_�Mb�1�b�����Q��卻�M=��g t~��?���З�5w�|�]H�Q4^vI�
�K�bXj�Ă�t�d׀�ny���6"�SH׎��=�lp��?s	�q��=��ߌ�\@
����]�\ɚcD9��@C����q�ؗ��`���9��R챯T���Y��o�t�:t/�U�
]GT�^[q�����4�	J�5��=�I`x\���~�`�V[	�ν�Q������b���G��R	dI�1X����s����JZU�s0�9��8_]&R�m����3��>�A�ܱz�Z�ҿKZ�m
��O�V�AT��_��T���%�)�����ğ�rB#K�L�/���C�QP�[r+����L�:|�8�wl���$��"�B��շ4��&38|�I�1#v����>�{������6T�u�!����A���CϷ�	�{e���j]e�*�ό��$VT��#�	�C�_�w��οP8i�`���ш2��N��\�a1���9��.��7G;d��i��c*!F��0}���u7�|�-E'1$U
IH��.�EcL��v2	��ȨK����Zx{��IyAzV<��W���[$��UÉ"����p��%?7]��5a�]`�2���Uu�M��/s�r�/=��Q˒ױ[W�޺�t&��뭸��#c�㣥gA0rs˿	�zo_��xCd(��%��Ά�~O��c 9: �{�۸��fv���wA=�%&~�+[ �c���`��:�jP�Q�1�Q]��fv��ǥQI-0Q	�ŖG� L�VH��;w8�٫��PD��'�ƴ�{�G�6���>�Y�_�'p��s$��d�2�1����"Rֿ�4�A�6t�Q��	���q��x�L����0o����6`�* ����8�b������6�`�U&]>+\��'g��_�HHH�g��)\:�D���6#�.�~F�c0S���7©.�U�ڛrğ�4�&���Kud��Ir�s&ecT�U; ��Bj|����`��g����4�����b�6�)ulN|4}�D� ��^qb�7
�~�`�U�C7ۖ�a����g�9�,ia"U_�cO�F��*8m�	�����8'�=b����Žy�-��#��  ��T����y�ΐ��[Xƈ�jqC�9{��;��F&X"y3)E���-���͋�4�kؚ���6ǪK?<\��A��
t����L+-mBǻ ��fy׎�sTt%���T�{|�_^KmU�z�<>�؄b&Q�D��\�'�Q��v��ݵ�۩ ��w�R�p��@��+���̎�� ���F�ܾ�Y���$cU6ݺ+L��F�d�����ޝȽ�K�����d��+�J�Zc���־o�$�U�J9[����5Ga�	}h��l·�����f���6i�\��MMÍ
��������2�l�9�K�:@�9`�C_qዢ��d*ӯz�R"���`au���6�i�˙f:��2�9_%����%c̣l�|ٌY��V̄���3 �c�$�Dn�xѱ&Q�؍�1�.#^���1gլJU���u=�/������%6岠�gM9�	F��X��T����������%��>�j�t�`��IEyf-໫
��9k�Jq���cQ�J���Q�F߽8�r�s��,@��ٛ���	4�C��R-�X����	L��!#=��}$���rn+�8���廚�-��įS桭�/6衊�@���R|"Hn��y�ˈ��)�\�{p����p.�ϡT���p0���.I�0�k�hH�ꋜ֗ި�<���BĬ����&�A�}���H��_\�^AB��:��=�'� #���H�ou��=�q7�#L#k�[�^L���?2<�ne��:xMhn��� 0���J���A��6V��2��Uqa����3H��V:��y�5�`Xɉ����(�?������\ 0ǩb�8�5�3)���so]���<���5��̌!a�\���;Kю:-mH�j�������	%]x<bDy��X�+���M�����ɲ[��6(&D5��k9���>�q="K�6];w#�]1�輴���~��"t�F1��Elt�	�g/Ƃ)�T|��.v��g�F(�Ƞk4T�s�.���m�@���s�6:'lJT�2��-$rmJ^�X�܄�ܳ�e �-X�����
��}���� �6_���mk��}��R�� O!��!M�fqE������F��}A՝*����xP&5S΄ܬv�k�Y!��kٚ(���jXZ�)�Vfo��̊�W��l�K�w����W�Y�7��s�2�����N\�0z�p�q�@����;�aQ��s�<!��p��Z�>*0J�{�`H�O;����ݒ�䤃�Z �'�^DsK�M�h\EA��'�%;]�,�E�� i?6i�~�i|Qt���|^4n�c��f��N��Aҥv���3�,��-З}��yr����� �f��z]nӧX�3�Q+���W }�K���`��Z����$�=;
?G�����mF���n;�)y�B�� ��;����WI|~=2B����x�$`w�7���J���-"�a�������ң"Q��i�b:��;��
J�@�۵�E<ȝ$�rK���p�:-�L� �`a���������ܮ�j=ٮ�'�Vi��0���&� 5w3�������v=��^��|��d{}{1�T	�x�@Llr2]\"�7�Y�(�p�'�XU1(�vE�_C�����+����Zxyҭ=r��3b���Q�͌�]��6�C�� ��&}�|_�v{�V�ǡG����h�WiX�����=o�[Q��!���QB5sy��tS��,���	�v���T�Uh;�w#�T�C�e3xϺs����ǿ��g
-��*f�UD��j��޳ �DK�w�jX�7S��֬/ ��i^��2��G�����1���^9���7ct
�c��]	E��Q�Iw-�j�"˜!����L�Ij*�@H����^Sc楦��'����P���>4_�Cs�װ�q�˓9n��F��H��q<����Y��XD���M�n��ތ�]�M#��,�)��!��M
�C��)+��@��y[�t���y���ʜ�ǱDv�]���o�����޶�>���]t�������&����)X�n{vX�웷�K�B��k�DJJ���������eoj�p���>����i�"/S��q�[���S�v��\�u��סpW+Ӝ�=���c^PCI�xo,_qǂOJr�e���\�t\�ō��~�!g;C�C��}1�����*Z����]��m�|a����"�We?0���Xl^y�61&�&�q�z�ɉ=�td�"�R�1�||���f��\&�#�6�|��{7���l/�K`��[�x� �yt��u�Q�s�q�x�l�+S�`�uEM��b6n�.�;��<�~�gކ��Bn�Ƙ�F�f0E}����h������Z-��2���j�8H�!;�Ύ�퐎f���ﾚu�$��?x�;Ud���yp>Q�<SEם��md��2	|��(wK�������e���hg�[��*��#�_bp<<���l�"&�aɶn���ar�}��G4�3���4=���[��ZA�d��4G��4�\rS73�8}�}��u7chK��LO1t�ۍ��ԺOnN�O�0��5:�s8�Sc9>0�d��dt3��s�E���ua��q
����:�z��?�qq*��z�f���(� '`;\*�Nt� Y{V)�!&X�2	9��P{ʵ����H���"H/x���
����.1����n��BJ޷,�N�Ϭ���	n6F�P���+��>f 0������ÎL��xٙgD���VM��E|[r�H��`��E3�#�ՠ���@
z�k����S+yzt֑�m+E߽B/g�R/�Еq)�wP
�� Xi�F�'A>]��k�����,T6�n��D�`_����(��E@�����_��ω@]�M�?���7��p����}Q�ػ�/�O�[�!��3�C�JY`�NV��Q&�o�~w���$��N~��;��K��� �j'U�|��9:�w��J�5��]�&@r��#H��~�dY�ڤ�W��i!*c�0&������>O���#�a����]3y;��rY�u;��2�c�hs���,U�46%���0�=0t|�Se�2{�MEυ�?M�.��屼Xp�8�Mx+��f��\}��z�v`��4��IU�;�[y��t���j�Fyr��j�9K��#(�����T�qJ!��hJ�� �hobw�GγHX�#0',4�B~V3���M���ooLs���A-��L�!��ʧ�{��:���Ƀ�2 ����	�s��AF6�*���0{�0u[��7��a�U��	P��/LD@��W_`�.�V���&y�2�V��ETt%��*��&���\h�P|Q�ǰ,,�`#�ϟJcm�o���U�㼑dϝL���ʦ���{��\�Qz�m�À�^a%G|4��=E14��;�л�̪J��>T�<���&U�5l��#'���2�7ds��)[���o.b�þT��Ky�����+L�#d���,uꊻ�9���<SQ=�X�RZ��"����E���X#�s�;R��g$p8+��]{.�FR��p����X݈U�������{@��(B���v��.TJ�I�;4�n�C�Ń6�er��������jgjZO<� _�D�˛���,ne�#5e�43�@����~1_oELck"|+!tV0��M��N��UF����j,�
zո�\S�nS�d�ţ��9)�G�\���[.�mzڒ7�������vl��=�"X���Jo=j�jb�i�Y�C�Gwh�/ĤL��� �hL�����0�ׁ��=8H�|a���:�y����O-m81gu�%XdBDM�,���öM.�݆���@����_\L�2������L9�69xtc� W^�9�SrbO]B��q�5�Q�v��Pvwq@����bp�aY��Z�S��;�e�Pڗ�`s�	"����W���L����9�qN����	�H�s\��݌;PH5A5���B���'܏�\�T4����#V	|�xE�^ICXm�M�N��W[��[V���N"�$$��6:�C��hT����q�֖��=\�6��ǡ���)%���w����t=���!�,3E�_9>���BK����Gr���C;ˏ�a3սA�O����(VOJ�z���}�3�aZī��e����Z�6�Uy��k��f5P�ru�:�T��񈤨����&$@JО�F:���K��a.�m^7a�p��m��0�e}8t�c��OP����.�#��r�^x����(�?�;ӏ hJ��aA�Ε��4��%S�C�(��i�#���4(�7S���d���* �@�`���l�
����\�,@�Ԋ�Yz��!tzz$�E�0��'�mj�-*����6ʉ��:v�`{+NO�S�#�K�h�u��Ylߞr(���3�_�a�M��ުQ`>`a�;!hR~�a�BvW����Q<P$@ā�<�9<E����ZG��B�œ�r���s@���z����"8� 
ݍ��!�	8o�v�0����-:j�
��=���M���- 7������I��q��-�_X��v͜*��^\����
u��_#��Z赲�ПcR�HE�$��~d8�,{�^�,�\o1��{���
O���W�Α�=��g{2Ҏ�1[�\vNv�O)���>'�"��US�=�̨�!��?��s�����ѯ�$p�����%J;vO&~)ޤ�ۖߌJ�Z#^�(�wLT�lzuZ"; ��:;uh ��5��(N���ܰ.V���¨�?"a0V%;�=�Y���IS	/���ܔH~�3��t���jz��?��9�4Ζ�ַ�ȭ��>�ܞ���hUֵ����E���	�]8��)�O�l]`�?1Xyn&�[�=�${J����F��)�l;�鐁9T��*$�.l���*�<����"����;�@2u�ƭ܉�*�fu�חQ�C�)>1}G�q���M���czA��m���v[�j�RS�N4�#��q�ǘ ��cܙI�B�a����m(�����z���bǣ�����l����U��g$�c�l/�u�K��_O�.H���KZ[g���'�<9�ڷfY�A�TFX����_�����]ukL�[����t��W� v�d�*ci+>�,^�3X�s5�dx:�(��a1vc�|8A1HE8>g�%Ɨ�k���Uq��9�u��6wlL$F�$�u[U�MPO`v�1��K*�FW����E)"���- ��i���y��q��-�d�*��F�dB5�Ǩ6�B�j�%��Ǳ$b�;���Hl��.l�h���#0C�0���#�ҫ�cR�\��)x��WB[�\�(��Ɣu)�������Y��qA���咐�t�ӱT��t�3���b��M: @h�#a!�
@�-90��Q���"��a��zYo6WR�c�p���W����=VPO����&`'x�D����i�5~��tj� `�40A�4��t�����sZ��!�u��Qp%X^|�G),V|ܜr�/�Ћ��jخ��l�b�5���E�SBwV	(���G�7���\�}F2k�7c-�W�,�3|��H�Ο���#$���>~�=H�m˒�fYh:(��i[)�J}�|?>w�Ț�[�x�t;VD!>Q�krܸ���I�q����o_�i+�᪍�M
��.��O�%�6�.3�`#h��Q�Kf�%��V��R݆r��j�vN��ty i
L��[ۈ��'_/���_�/���a~: �-I��,)Z�OW�_�E%��zŜ��A���!���%T]��Pd�	�h���z'�L��܄9�u��&��ږEQC�uW�a��1Zh�[�xl�J����X4���UI�gk�*�,��QJP����5��y��$I/�V���h��b����L�91���9��w/W������sJr< 򌏞�9n�7��}���/��ꬲ+em�3�p�c�T��j�З���!;��:��`�i�|	�nYY��RSn��ڝ,B�e�DY(�C�	G	8F(-(��"HvF��<L�g����:��T҄���^m@9��K	��B����%F\��W�R G��Ɇ��e$ ��L뀮o�*�\O��pp�9��o��Y�SE�W��焬ښC���W��7��sJ͈�+���yJ�^|D�f��7�#8�ވ߮��hR��X*�}Z��ʃ8A�D�&C���Mǰo������hǺb�U�S륹j�Z��8�|�yZ�[�ݎ�=�>Hq�_�B��ꯉ8VGz��M�Xd<S������2q�l�ݳ�)q)�]M��4`�i}�|9q��
�!C�..�������&��j�T���0oB�vb�)�	ᶷzʋ�EQ3᱄eB��l�ʜ��V�\�8�W��06��`����n���N/n����][�L�ez�W�1����n����"�\��Y�8�:�+�=���瞴�M�N7���
�˱�[J*�Ep�l�D��^���^��Tz�F<��̗�X�"�M,���08��!�X��O��ߓ��>f��]"M徑xZ�⒪Ϲ�ׄ�ޝ����|~j)s�	��x.��Q��S�'��u� M���"SX�*{Z��Vܿ@�΁�r)��t������u��E��Yw���yx^�[�Q	����MaU��o\h;�sNĥ�X�1�e��Id�s����V��	cn{���1���y_4��r�mǢ���>cB�)UӉ�
�J��犯��T	�~���9��M��:
@�j�!���ABt�!�rY$[�l���]_tx�j�H��&��d��;��M�YH#㴜�/�F��$�cu��\�Q	�͆-�D�!5��E��|j��"1R�׀+}^���� ��G @��]@k�Z[SO�p����fG��j�dV��}����k���~bK�C��XgW�I����Xm�䉎>ST��4��OgaC#�Ñ`�.�-�\L�#��9��U2��8�K2c���c�������g� ~χ������0o����y4��)���~R��Lq��Mb�p�}�`��\b��}�+Cl1�+:�1�\]2Cg��ϼ����o�aQ�vyRv�nD٧����H�l+��&�[�4p�����󞇌���i��MR�#��2�赉*��Vq��~��u��5�n��4;��C/�{����B��(��� �]zcK��lI�|����_ۭw�
�X����~���dn��Y���M�vn��b���c"�0Wk��XQ�՚ �U���	}���`+�`��r��&�nUfX���ѓ��S;t=������Rr�<#y���A�s������5x�4(�X�Z�<�bS?�&g[���|�!��� }-"~	�?¦W���Z����~��"��)����h�&���&���Ԫ��b���+�M��RG���iK;�wL֗���r��
f;���ϓ<5�X��mZ��-?�ǝ��@����d}����LZ�7�g?`շ����������e���v�R�։`eC�;bDn���hQ&�b-����:����}#�S8�n����D�R��}~�ST���ͽ�O�D�;�J���(C���-�$ґP�,[�fX���y+�� ����h��QRo����[9��)�@)}�t-d��f���V�f��@hk9XL�`��&��o#I���k�B/y�L���ׄ�W0�iK'��9J����Q�����g�'.R��߷_G�T�/�fn�i�ꟷ�?_
W���x��r�0'lCnL@���[��`|t�D+���S���5w��Hwy64��m~��co�X�{gd��0;�Lϰ��g3 o�hc/���� �G�ܕ͒�� �y����1�)@�5��2�h�Z��3I�B �8vŶ��G��MD�ϵL��x��1�,����.���$��P ���'�V��*'m�{�G�0��!��^`Z1�M]��Yh1_^��D,���S=�o�y�K�ޒ�v��~cQ�5���ݵc���Xͤ�xq���sQ��U��Z��p`��T�L�ΰ�� ԿU�_cE���n{�kRD��L<D� ��=v�d���<���R�{���[d�u0}��6ƫPh����B,7B�;�E	��u�Ȟ�`% 8�/�������Z��No���L�*$`7�!�ܘi0h�6�Z�&��Z*
"ƨ�$(o�x���}���ɗ%`���S��Ӵ�"�c��͑�֘ޙ��Nu�:���M���u�$sMA~}���m��{�����"6iЋ��?�a��WCU�*��G��@�_.�(�ⱥ%�>w���EYƮc 9h��<88��,C�A�
9�y7(b�'E{�����~�q`�����)j�\����2��>��+'@A�Y�5/����Y+��`u�Fv�4	�?�!(���A'�B����*J`j.e�;0��e����SZ�NK��O��
�o�	Ǚ�8�T��ؗRCn_xE��*�n,��������ȗDD��(��`��+���{�SH�2Z|���>����)t��k��s�����l+a�­�ͅ.�UQ��Қ���� ˨��f�N��ق%�tr��TLڔž�A�߰	JA�4��L�`�?���oo^�m��k����m�����u@��p�����W���e5��ï��F]N��p�\���O�?��u�2v<����ꟽ�y;�{�+x��*�6k�K�zŢ6��(�t8K����z�^pE��EzJ�ܻ�S퓅-��	�������ʨ��	A� 4f�:A�q+� V4�!i\鱰8}n~[�����|A!H��`����]e�=�ǭcK҂Cֆb��ܵX0#J�� y9�8�����M�,�S1T�rT��a���u2����)�i.�k5��Q`(ې4���+=
�t���! ���#H�F���Щ`���^�z7��-6=��uU[�؝8�^�3�h6�{�����Pwkx���z�TU�?�G~�]����3���}(UG�ʎ
�<tw�m$"t���0��^����ɑ�Q:���60�J50���A6��r�J�!E����t-����+���Φ���0��9�<�UX�I%��&j�;���]/}��!D2P�
)�/G0>�I���cR�tok���v��Ss�0"�µ��x�pJ'�(/)���z�v!��rԬ�Ҋ̠s���`;�f�����5@R����?*W�r���jp�,���O�=�^_<�o�V)
�����t.� �����W�|�}#��:���_����C�؆`���pM v�I������q�X˭��n�*�k�ȧ�����5�G�[�-V%%a�+���&��m)HF�`.���p�������^:C9[.%gFL\��s��4a�9��zk����2�H!)ӌ�w����ՐG��4˦����/Ӎ��<�H��0�o�[��0�L�5�8s,��+����7�W����3���`�A�M��{�`wt��2�U��B�{�Ƹ��D�2=�>J:=�4�[k�K�WM҉ �#�5,�~[>�W`Ϊ<9�Y}_%a��5��ń��09��:3X>bן�t���w0�����x�����W�Ô����(��.@��~���i�ε�Ja�>���J����Z�<Y�uD�C�)i�N�{��8 ����	ؖI�0!F���������.N.m�� ���9��Ql@��i��(�U g_�X���_ ��~Vjd�ۦ���"gᣭ	/+²�Y�
����%d{"��7D��5Ϣ�D�U�J��@7����h靋I��Kt�[���h�W�]�kG�Ż.m�N�R=��]�f�OS�ߵ�-V����7ֈ��(l��n�)�,͂�čŌ�}���Sԡ�3]���v ��7J�����~�!���<Sd���]��-A*�o.�H�ZUS*�r.ܨ�23�7�	�e�a�9���=�����U�'�S�1+:�(en����Z��)2�_־ch(Yp��^����&��������9:�//&�2������ƍ�����g�X�QA��|��a��?�l,h����7d����<��KXZ�K��������jY��;m$�-=�c��;�i=�/!&�*%-����Èt[�yi����P�و���J�2��/���+�̫��g"N�]ϯmKʞ@�J;~2�0Q�@���ANh���>=�N��a2�ě�_�h���Ҋ¢��>��r������G��� 6�.6��a.�L�͇�3��|�~����麪�3JD��\S�@]xQWx��a���t������D�o"5��2n�K�|@���K�B�Zi���1[��79sc�6Ѣ��senQ+C�y�Ž݀hͿ{e_E{NsE�Ԍk��5�&2WL���'��울DS2�vE�#v?,�;�M C�m�߮�6,��W���x�cV��OA�ս�G=���>�,
�?Y�����:���S�ӡݜ�>���`\<��hg6��|����)$��i٥f��e+Y�'��� �冪#�eE0ڠ9bϐ��?�vB��s���<����	��~p���H҉�<�h��r�'��8��W���YR�Ю��4U�.˕��}cy�y�������Ȋ�-��;�EO=��s)rѭ�ɵ)A��2��5ÄAzbfqHo�z;j������s���̙��d�;��S�F�.*���VL�l�O�E��� �I�?���EQ�]�� kd�w�梆�ƚ���a�"�d��{$Y8i�	e�6_M��N�B1ot�|e�k�n�+ݠ���,eN�	J�`��9QOU:r�'���������Ơ�����<E�_��?a��^���9�]�`l,u3%���|X)ҲۃV�� r�����&}�3��|��m�/fB�N)��A �(�Гu���z)�#�n�'�U@���ϧ��e��b�_E���(�8��49�ٴ������f��u���Kq��͟�e�O�!𢚸�s ���y��p<hJ��s��e�J��l���1�s�5��O�5��uI�H�'=41�nd{�H����=�ahvJf������["ʛ_�t���q�pJ8�L��	��P$�F�� ��VX��D7V�˾�sf[�g��ǩ.ն;C/�g��_8f��M��t����:^%�(��%�_�@�tN�L��f��m������CJ"�b��R�]-ʽ�yQ|>�t�hEMTO
�Vf����|:�R^�EQ�b!P%�<���u4��F%��S�%��4������p�IA�i��:)��}��N���L�,2��~�5u�.	���¯�Ȑ���	���lRKj��/V|�H�Y�j���j�'�ߌ��ի۽�\h$���bZ �2�u�M.�p{�kAҰɹgF}R0o`Q782�?@�|����u&dj,!��20{�<3%	�o���X��Aӹ�$yPC���]%��Ή�Ο:��� b�����d�\�Q�SD�cv�%ԣ��IC$�����FAo�oy�)�@�x���7�3@�h,׹$����5K�6?�G����A��&A{VWUJ2wY��嬍r"�%f�B���<қ�?bhU��
ѵ�~�T���n�~�+\S�vax;h�-37�!��gIg'�>�-5(��+U��joL�*�����$͔���~[��\9SF�鵎�����`�'�ױȴ�=:�I��7�XK@�9{8b����W�V$�Ǿ��]L���ήΚ8�.~��Q-`�#�Jx��aj�Æ�4�=�� B.�'�,N�Ϳ�پ��rd���PJ �K�:���M�p����#k�R���֏h����@ ��Rֽ>f��)���)$ښ�ћ/m�z��(V~1�[�d�;��e�SZ��w�M��H��3���
hv�o�N>lY����\����b1�1��M�'aW${O��Q�K�����?���N��8E�,I쓑V�נN_��*[�¹�W�|���F�y�N~�j��ET�PJ̽���}預�t��wmaG�ev�� V ���	�ˉ�&���v�3�)1R�MzS��kʗ�B�ޟ�E6��R�Ű��E�	Q���"�S��G��ڡ�M.�Y$�g��V���v��\� aI���Z���C�vb:��!�{�w�Y�=���^"e��4�X�.+��e��:Clߡ�+pD�_৘q�nVrB�=�R�מp� �/P�a�8u��9�U(u$qlsZ��D���Kk�.�B䣦Ps{v(���v"�|��bxn�A�X;�yЁ�ɐ�u��i�/p���wT���p�E�y��C��oq�޺�]a�.��Kl�w��=<�=��
b{>�MD4�Сׅ����?0���)?6�I�V��4M�.fl��;�s��"�R�<�ɴ����f!�C���"���o�ٖA�D@���̸έ��Z���}��$�'����%�bP�����کK34���s��r~e*PaS�'X�οs�M�VBB9�Q��RO݇�A��?c[Bs����o�
�]���:L�'��婿aU��"_����	�CBT�������m�"0	TԠJ0O<��}�����\]�\]� ��]�����WΟb��b�=�2O�F�WT�C�}ĉ֌c�@��C�y���j��8z�� ~��ͮoY؍|^�����iI�VU�- ��P��u#&s%���|E�;ݞk�hq�|Y��
��-��A�\��	B�yw�F;���>��#fYj%t�ꄏx� �^��WP *�Z6�%EUDղrsنO���{��8���-r-���Wn/�)U���
��ɕ8�~�d���p?3��ND����7g�q�w"�*�6�+�q<�����5\�QETH3�,�����*��mʫ)�X��-�ʽ'R���Yߩ�~�}��W���(�)���$���&�-�W�Q��GJ��8O�q?���#�9>��ؠgz��S���E�����o��B�le�U&/���/m}�xɰy��;�� `���T)n0]�Qg���{���:C��c�������-On ��ݧp��)����k`/^���	e��?�ŹK��){�̻x�B�5�u�ԥ�d��f�i��%����HO7Ҩ�c})S�DlT��#�x���o�оNL]Kg�N�,?��	���}z��Iw���3V	�Y�����3�0I,IB�Wp���x*:�seo�* v��C.�yr��]���V���~G���$��I�أ�����������L/K0o�z@.���ּ��^e�4� \��/�V�����+�د�$;t{;��~D;6	��Ш�_���zjl�?��v���00��>�b�T�A}�K'��b�X>�Ă���eChg^~��1���&V�	�^��=��ud���M���Z����Q��0��z�:�8=����������`�J�g<P��H*��+i@ҽ��E������V�ż��%�K�=��-g��աcǓX���;���g
*�r�2��jh1�I]�̶=��@͗��hh�[�h�q/"l�BE�	v�2N'ier��݊��������jr��I��ooSS{�� ����쭵(���\���`;��L�2*��A�'��)}_��2ax�A-��J��O�?��o�P1�!�@��0�#Q]��Kr�F�$\�q������5s�G���+J���%X�^.{|Qd���ڬ���F֨'B�WVZ�:�Y����k���K�Y��N�2�ӰԨY�xV|��o�|��n�\$\�������VL���c7�Fc���t��n��N�!1G���߼�|)�nm[��c���rMK��&���ڬ�I��fD�A���(����s�L����������1ԓY��Ъ1�&�����#ZgzRI�G�PU��e�yߒz�-|⒮�c����?�� ����5 �����yK�Aj֎`����
��j����N���>4�
qd����l�ٯ��r��.0�H��j�Mb�����Q\�a��;��7>��׮VÝ�zE}Ȳu�w�6Z��[+��\��R������-3
�ʼWΎ���8���N��Spgv�I�(��M�#d�h��Pe�!����pi# ʷ�R(�p<6�P�Ni���H��)��Cu¾�|���q��p�/N��>h9w�?�C���	K�^�Wb9g��
��a%5mS8@�muщ}#t�#�e�x�0�3�	�b�4��������Ȕe����Dg������/s*��<�XwѢx�{X}�bjr�h>���
ѽ��T�I�$��5<�i6e��{Kx����8���]��+�F� &�jl�L����k0d������k�)����*/aS=�?����@Lf�j'��z(��i��Y4��>���z�Y �(���Y�ۣ�h7�HǊ�*�ZViwCR���E��{Iq厳(r�Z{MWĚ���\�2� �O��@�ZR/��_*z��[SЈSُْ��w���'3q��)
i|\ʆ���z5��M�1���5n���T��z�fD��7E�^zP#���P�7DW�����$q�u�q�v�&���K����&�	��~�8�x��>���\!����H���qT��fy�o�4���݁[|h���礴7"��۷P����Ym�O�t-X�-��g���U��	Tז��Da^��h�%�:]q���P��lT�Kt����MQ�M���vd�j�&���~e�/.-xŃ�.�q7��8���0����z^/�o18G�LK�w6���MIƠ�Tn��)*�<6֏�����W.�^�v��B4$�bB��]U�mq�	�"��[�����'��Ϸ�ؚ�օ�KZ�`xJn��ɸ)��+��_�+A/�@�>�]CMO�%��o�+��,�4h����a9����5o��%���8b96�O��p#t&Rr?�1�YJ�E6�R�!�'na���"�(�5Λ�Tk�k~r��W��/-�Zc��փCv�C?���F-��\4g< ��Z��%�ۓ��9�G�Y�@�AxN��O���'�^}����U�~�e�TU��M��ɼ9��9�Hn�{T�^�{�ߏ��[`��M�51Ib������d�C�d�~��ݺOx<u��X�ꕮd�����"90 ��p�E��t�i����.�� {�K.�5J�����2�T�ɞ��!�4��UQ[%��Y���d��O23�����XEY�	�Ȁ�z�w�����ƚ[��/A�E��[��GW��R��g�����SE�_-Y|7�Q����(o6W��ʦI��iC�������@=)��BX�3?[&��ׅ�m�o���� ̌���ˬ�����<~%�[����m��р@@G���@(J]��m�����y@Wx��Z�>g��&���9�p�B�ٚ�6h�M�"1��t�e���A)�)8�l;�v�1IRCI֩@<�KE�?����>K?�t#�`"���4�V;�j��^knOg�xT�3
«c�����g��.|� �T��W���s�JߪEE�9����
�b���e�=.�x�l3
�dU��Yw�.�ٻ6�>�v�V˛��NJ�=�15���5�AL~P���E]�B��aʾ����'�^�5KU�T��:φ�\�_R)�Z�6$iwp|׫���]��b���ƞ�3� IE[�Ϩ�&r3��o�^��d:�pR�]�x�%�ι�PI+$9��EQ�s�#�����. ���Q�I�,��Fl��*�y��V��~�H&�t=�Ī��Pu���˟P"���e�`b�m\�}o���+���l�7�b��܈���HY~���ێ|bs;��u�6?���(i-/0B�k��G'����� �X>�ݐ80�@��d��Kd.��vɧw/�N������%?X�a�Ζ'B�Q��X�fѯ=t^�F�)�V��i����ۥL�{7Y��맩_.��U�wG�j9�k��<���l2V��S�l�B=�d��?�����zkJ���x��P�{ϼ}��P_���.��\�������}�K�����t�x��=#�p�1jOO��"�q���
�m���A������#u�$n��KEh��`��PZ�`帢*��/� #O13|�Q�L��Ѡ����Gr�C_{����2�vg7��)��Hd3�)�0�:5U.�вm�x��e�C�T�&�ݕ�������$�íj�"��� �8w�W���� ��B��n+,����U�2��?�ģ�*��<_�� �+)Lr�,�A@-��������K䭮���c"as%��0����y�����N���6���O�V3	�gg҄U) 9!�8$�=H�?�[[Q�;AZf*s�0FF��Eq�3�ա�9��!��d/�a ג=�e�@�[���o����9F��b^`�s�]D���Pt�ڇ�i�p/ߣ�T(�� R	q���Y6�Hs�$T�Lg�}w�f�E�E[�?S� i؁r8q�^�7ߠJ4Au��o�9�M����T&���\��[qc�	����5���G8�pm���47	+˴$��j5~�J_n�1�ۄs�$�*v����l�,�#R�?�3��i��W��G�٥O�5)x��<��yF1���+��U��+<�^k碒��!Q\
����*��������O|�Ѧ��y��>l�~�S�Ð?�M	ҧ�o�IJ�Ӱ$޹Zz����:x�?kR5��(H��Z��li���;��d"��X�e�Ν\��VP�9s�|QPb������c�|�s�?4N:mb���]k>I+��9Tc �3j=\�0/A�(<��_J�W� i���ۀ��K����Kll�O��Ä���m�\n�^���"޾�ޯ�Q�+.}������=Q$&JJ������#Y}![��v�t���?˫5�R�}�_|�B�9�c����q�ѡ2�3���$(���2:~5l4�NѪ�c/�n��Y^�.�5��B�0L���{ﭽW���Q͆,����lI��k紲�W���ĺ2�X�c�������@�;�X@�Җ�Lt3�ȯ"x^V���������)�D��i�ak����J�hwɚ�P�ځ�s��YH�S`z�
G,�5=��!���3�<���(�ۨ��`�"�ݍ۱V��h�0J��k�W�h��C'���,kO�Bum��7�x޺�B��Cu�"*<�����eß����9�/�A\�	[�	,1�0���ro&e��H��Y�_���-���U�J�3[�	(��ǎŝ�n�}x@t�	�"����1��G����&���nD,��4Z�owlc�T�,|��tҌFV��l������ay�# 7�<�Jt=m�t���5�~�{')�p7s,(�:��s�K	�TS�x"�o��'lh���!!>f���?�>��Ch�I3�c�n�P�.29WH:py^��h1�k��[WI�?��zg21�E
�I��H+�\(���[�L��;coJ~5�c��Z�Y�+����ӏyCz�Ʀ�@�|�x�M3Nĵ���tʎ�%���<= ��i�bg�.:�BIL���3
�h&&�g��ǟ�(����L��>p �}p�����-L�>f��cD���RZe�#�I�'6HE�tt�`��>E ��M�ݴ��?!��n�0��
��W��Zi���̊T
��<�E ��� V��J����[�Dwc�=�$i����fK���8��(�M��]\���� D|cXj ���u���� cC��K£��nd��
\�)n�2,8�S�5R�Q�o+Dp���lpi���q���(Ep"Tk��R���M�`�9�dQ����W��[$ؐ������6آ�@��V�)Ah�����Ľ-�����K����6
�5��;\��\#Y�+�k��
�͔/�����=���R8tkӝ"��5;�YPČ���(�E��`���n�vwn�aվ;oYe�kdK�B�W�z�W0���v�y�{�:�[������]p �}�[!�kJ�)�<�.��--a^K/��^�r�E.4��c=��p�"�GD?>S�Ph�0�7���A���Y3��[���n�P��FծVE�~���׃�[}Mk#O�M	�9q�9�0�0��A���D縦�W�$��S�+����>��18/�f�uT7,7Sl�K������~f������h��u�l_�"ag�T���LR�U��؞Hwp�[s���A�W��Ci��(ع����b�ʋ�w} -cA� E��ϥs:s|����,V/:��^�3��ٙ�0��� �Q��Ř��C!��'	��aAJdqŦ��ǀ�W���G�8&ۼM�yP�ܕ���!Yƣ?�_�̤(G	���>xߕ���b+D���4VC��˙��tN�TVG�N�	F��������=�l&"�be}���GD3/� x���9j+/9<H� 	�E�}Ź���ڹ�tM!�]/�\,��c�����^а�TU��]T}t_�k�6d�Zq<��]�j 4�9t��R���Z���
w��Ƿz�=
W�#� �#���b��X���ث��-�-;��v���ftuTd&`���h���W��� �)��t��q�WsᲅQ7���Nl�`�ثi0�'|Evdܝ4s��Z츉����TZ�lp=M%��j�[�.�7}��.P��a��O��(|]y����IB�aE���m���0�%K��s*���X��Э�%vG���nRM�7Q�.���TM������pd�xEd	��2/<	%,҃|�B2=�sL�˟;��;@'3̨�H�)5m��FPBv�>/Uv�������}���J�ѽ9<��'�Z	P,����O;xϕ,�:s]�2��::)r�X�����X��#��w!���KUDL��
f�V�� �i�m�f}��Lb����7�>A�ܧ~A:�?{�:���A�+I��国�
���q��C��.��� �-�(��!�lV�)�8��Н���n���iJ	�I�z��%,KoW�\�uj�}�l@P�<����%��Atg��-]��v'�W�˾��=��1yq���z�s�����e�����=Ḛ���=�㎠�&�Cj�����hM��QDC��.��d���A&O���nx��+i�� �i��At!ZA��b��;W��L�I>�$3�w_�k�|��2Bw����R��D�gw��1�������(�!�/�7u�i|0��<-��t#Je���-��]�wu�|OPN��$ugP����Z�f��r����0
 R�r:߳���m��n���́D�%\=�"o����4��%���ܼ�Qe	�Kn����-�ڭ��KW� ���_��3sd�{+L�D��Hp�!����C�p�?�x�J6	�^��t0��Eiu���ƺ���"u,�Ip�w\]��fɖI��V������������YM{W�Je�9��_'��0�d�#WA4��l�#�j`֭D
1@/*.
��Flش\"���~�)��I��随�8�h�q+�ǯ�=۪E$f}�!��i�w�(s0���}.��r�G�G��TC0��<d�`M ��k@G@�/i�{�V��?˓XK�|��`+k�� ���u��	�X��J�y���C`�d��� ���!��(� 5a8-����v̰��?vk7�a;:p�
��l>B�<�Ww&�i[1�־���-	��j�4�i>�oS�~U�ܰ$N֭��[3�v�,�jb�8����/���:"C��9�Ay�܉��1���<�#Y�6�ݝ���4��ċC�Q��޵JJ1䬯���Np�3E��J Q��3������zya�KU-O��_Gi�;�&�`B�|��̷�z�D�Р�-��7tS��ȏ�w���=Xb��2��Ls�a��	о��qY��+YSm�~�9e�
m\A��#���b�����Y�\oN(WӼ*�J8�t�k�r�du�a�v�����-�u�c>e]Ի��(���C�����uN��s�wAcUz���>�k|������ɩ������V��g�J�'bD�[�Ĝ�['޺�Z5Nc�k\+ɑ}�f��TKW��Kg�X@i	��x�0�q���c�A�7>[����#Um�����R�w_pk�=R���<η��QMŨAC�]Oٸ��_���j�J/P�q����BV�B��� �Intl����f$�%{#�~B���Zt����ө]h5v:J�v8,o�����(߾�;�ŏ���{�"��4�MIL�fJ�Ʈ?�~�h�Ҩv�9��l��:(uh�ሓN�6G%�O��"�P��mzPzz�9���<�o�*�[���?����G�s3d#ZX�ޥ��3���f��8Aw�Q�tG)�ʢ�g�c!Sg�i)	�6l"MjCy��yc;Ҹ�E��U�W<7q@oA��xZP�D�����qJ�H6JIݓ�GR{�/* t9g�?C{āv<�E���}=����ArnәcHR���T�'\� ���`ή��)<�����;���6�-���{�'�+Қ6U��|��ɵf�u�p�O��Ⱦt�^���y%��hЭP23�#r���$�<-ۗ�h��|��F�余d�mf�6��!�����3(�zg��*�^���n��]\_qA>�H�I3�� ��Q�ba_z�ˇ����C���c��OAɌ��|F���r:���(6����j�[h%q��<����d�2����c�V�<1��Ý!昍�4�(>�鑋;�R�h�(������O%_iY5�z�3�o{�u%#T�n�Pe�'�XF�V�b�=����.O`8�`�4;��S�;�_��8_��q���D��&���e���B�N�J��G'��U���=�V~b�S,L]���{����ngG`;.����:� .��ha�c�ݭ��= ����)ώ�#�{���^��ށ[���W��\L̋��A���j�)G�E}g6��{�`|�����E��2��o�s,!;L�BͶAk��KU�0���̓�n8z����NF�n��6�S�G �"�S5�i� 6̷~6vy��3k��`T��|uh1�q�ƪ{m�X�"ѳ/^,/Z����;���+%�����ɨ�)��=ӱ���<~k�_:�`sM�5���]M� Ӂk��N�"EV�2
9�c��L/���E_w�w�G	uw*������`F�����C�9=E�@G%�z��+�p���I�O�!6b��w���bz�7T�-JW1Kn �x�buP�W>%�1�j�����v�Ӭ�b����D�;�'X7%��O�|hP�ǆ�$�qH��Y�����&T�K��𙜝�!�Oz��]��.O�s�1��d.Ї*W�1{;=�AI�mZUA�
A������a3� �n���b�o�m��ňS��!ĳS��&y�)n�4���4N��DמU=�bk�r�����-�D�����Ý�D����s	?�O�W��ϙ��s�z��>�	A��^)V+]_Y+pxje�����ޣP�r��%�2-׃�����O"���U������'�9Ct�I ｳ���ە<����OfM
�Ig���%�'x����A��������8���S������W�7�^��5�C�>�ϻ�o]e�_��H�c%;���I^SD�;�er�YjN�O�k|�>���2G�V�Eݸp��Ƞ8E:�[��:2)��/�rMa��vszhD�(�V���:��4P3/���8����uB���|ؿ�bw��.�)\p�|���>����M��h��/�եVo��mM�1�:%3H���xuxc��J"Ҭ�kWkp�V����Jtx�����I�鈞�Wa�h�����\����������
a�@�gK�W��6�»:�`�����5ĳ�8�/�-��.K�٫��n�H����m���q��p: ��X�śfV���3��PΏq�Ρ�qnך����rh���ח��E��v�!��> ��xk�v@��e�S�u�9�g����u�&%8<����qޯ[]�h���V7��|\@�Xe�/��7;"h4���h:h����٥"���H}"��֬�Wր.�`��R�4�{����cRL��>π��q�9Z�?�}���&���R�4��673�4�z-�E�?�?����?H\�ˬJ�x,�w��Ă��z��#�����V,��")ſ}�+�>u���	 [���4�$y�r����О�]qpt��^B8�_�M$�_�<�I.�~�iY���n=*��|��no�U���-G�_�K*�0V:A����T1u�� �<2��yo�)J��p�"�ç�A�Ր��U��m��NqT�0�a����{1՛�6"�@��ހKx4������h�ў������髻�x�7/�I�nߊ��(����AY��CV�u6� 3��S�CK�ސ,�Oc��L��lA����}Mz�D��7+>��`�襤�eU���l��߲1 �;{2<�,@�^6V�]6~x7c$���QJ"���#�Sa��.YB�P��cd�����غu8Rf�Vq��D���x6:x����hqz6Z^�ZG+�0�ƭ��T<t��58����La���Ϸ:]��_s��I⩸�cA�V�7��7Fb2Z��5B$>��Hj���5�i��#N�H��5xZcڦ��&`D��5�K���R���w,u2Y���2����!m|^��z��oWEO}�����<�T���$�����׃�Hm���dHo�D>V5�7�M�١��E�>��ף���[�y�IV/ �כ$����|r��ɝ(g�*8 �{�txBPQ+N a���_\6�|�Z���d̼U�;?	+]H��:B���-+l�-�zVMh���t��wEI38���^/�ft���@*�ګoO�U�n�ګ��TMA6�j��(.�����m��M^�8�/?�G[��*N����S�~��}-��GK*��z�o�\���Ϭ-���uX�su�3g�Ço����e�>r�qU��&'?eҴ�����XW��O�N�mG%Jn�4�&��=�C�uC���B��A�{.����נW.*O5�Dd;=�r�d�yM���=�L��9!�곛�5�6�'��C��W#M2�t�:��B�Ţ��mgz-͖�%\�A��?�����*�\��% }R���t��[�{��Gm[�@�ڂ	�Zf%z�R��<r���K{r�Y}�s��?")�B�5��J�^���G�uo� ݊�J*A_�"E��z>.�;N�&v�J���
�-:T�i�t�I7}糭����L���[�Dă�
g�߽���ʛ�7t?�5X�!��~Vh6�F�` O`�B(֖�?^������Kd��yJ~��y�����ϔ�14��~{��ȼ;���4Z4<z3L|z0n10����_��J��F+�B�A}6m,���"�y�MH,ܾ�"cD�`7dA�^4cQ'��a��%����L��y�WVB���x3�����}3���׺��l(|�.�H��07cOpu[�iW�:;�PR2�n�}\���AS�e�X&�1@�<?JcǇ���QP��3�ܚ�Vw8E���.��k�#����k����#�w�j�z��ԗ�����۞
I��^����V�D�=e3u�+"T��Vô��c׃�j��^�xF��j ��zn+!{�J��~�S��h����V=��5x�̆O_P��i3\�ˆ"�9��00��_+��M1��i@t?T��������~��?���
���/��^	���}w}䲬*AkTA�3ܺ�!�8���.��$m��.s.P�b�ۤ�[�djZ�t���<bK9�ً�ۄ��A��}PI����w�lf7�l_Y���.x�׃��@�;y-9(�USJ�T��C������&����;�$^�^{��-�)�`����~-�!g��-��J�1e���S�]w!@t����Y�B�ɜ0w��v!<��nm����2I���4��,´M�Wԝ8^�3*ͤi�zɿ�Ü5�h@k�L_Y��F�j_�:~A8��~��͡ 3vk�yl=����܇&������)n1Οt��Y]\W�yN�^��Ɩ(�F2e;w�uj��|����xs���.%��U�s.)�g}h���[3�WjN���֞���.:�V����<�ey%	9���&�E�W���5G��-3G�g�C�)]��+��A�P�oc`HD���y@�Jn����k�V�����>����(֭���~�G�F�h��h"s�tk���Q���i9<�<��<8�:�Ȳ�W1͟�D��D#�9�#��]��F!7�)�G�)���Du!��0��:�	P��q�{U�i�|x��T���9%��4 g��8�V�n��ISDF~�Bk���:Ib_��w�l�7g�:v{�&���>���q�VU��:��Q�:�������-N����R������k����J�:C�^x��/OE,j�NSE?�J�C�u+��̟L�씈��j�:�D�/��e0!m8�Є��L5��&�yN��j�H�Y����fB�֢�@;z�IW��K+8���9-l��Of�j�.�GN�8���"bW$����(��t�s�3ɣ�ҙ�Y�uN��W�i�*�7��:��G��X��;Ev�lYV�W8�U�0�Z�:�}w���~:f���"',"{J�d�~��E�/�w�;�ч�mRR��VXjNc���"����u�Z[ʋU$�������s�o��O,�j,�Pi!?�Wdh`�m\)�P�_�m�]�;܏ݡ���6]��I�NE1��[R*mC�8Qh�����If�8��Ũr9���;Z5�����{�Bf��c��\[�:ԧ!�غ5e�"/����^�G��LR������"�J�CO�c���8'5�Yr��"��Rk�<�*�.�b��\LYS�p�a�Kv*���/HT7J��?���ua��i����4x��n<f�fi�[%� ӍV�E�!�����@{�(�1�����Oi�Z��82�u�u�Ϯuqh���A�`"@�<�m�x\2�'�<ͿՂI��O:&-C��d���t�Bv��%��	I��^+:��[\ʉ۲��\�� o{z7���;����22F6EfEנ��/}b�lMw~Oj\�v��J���
�߭d]�2J�I�3�H��'��ªT��G;�j%�z.�9D?sL_S�e���wv��"\噫!h��K��$y���)��ԙ��/%����a6�2f�ޜ%8&�	�^팱`�ow����#�`F��ؕu�Kx��'�T~P2Й�	��j���'�5�a�{�: ;)6�+��6C-
��=��{�3H�u�O��P3W:�b{��1��L���
:9��hB(Rӂ�ڿ�9�6`jb�!��V�r�����id7lJ�W-�]lc5�hמ��3bdK�6&j�[A��UVC-���a3im�a��_<gi��>,�F�@z9���==M�,��a
Q%�k�-�f��/���%� x\p�e�k���D��z��A4��T	 S�BQ8�T��Ke��.,&��n/$����}'�Ŏ��)���[Ь�[rb��Ж�o,�5�ƈx|�M|H�����WX	ژ�#3����o��N;#kl�w�l�ݻ�;eUB�3o^�T��&�f�UH�[�?s�<?���E��z�&|W�i�����\l�8��,g;-�7���K�i���_G�1�����+W�}r���*�>g�/�!i*�f�˺ՙ����<�TD��6�~q��7��?{앀G���%�����N�vQW߾l8�3�iW�"����kivS�D���qe�4���pv,��u�ha��U�-��&m�z=G���r���"�OU�����*�(�)�����ї!��S�%HP��
5�_���xf�å��b�b
Bm�{`]r���߲��kB�_wխ�N�V �$n�W�
K�XҏwR�'T�2y͈Bo`�)6�K���>�_����JH���eu��_�_�?V?��
~����X3*LN���j�|	j6�l��;�ɒB��6���괱E����r�d�"�ԋn�9�V�����u@pP��m�%���窼FZ~!J����L��i���(�j�b��TPR��J�k)1t��`P�����K��I!���Qlx�7�E�9�Mge��n	�C>�,e�U�Di"��0��$,Hs���-f�=��A���v\H$yrRAXWF��^�`�K���L���ӭ�*?u����u�*S�1��C{3�q'o�i��g'b�hʟ2�F�H�m�6�<�t[���ǁdb N��:~�z���&��:"mUR	\g�ْ�W�z�c��o'���+C�l�P)]92�Ը����jCW�G幣�C�P�XD.�/�T�~朗H ��^S"��Y�M#���	��zxu�Tl��K�dH������dwI��}��vvts���� �X���m#��H����1�Gu}�/��f�:ޢQ�-2���\'�#S˨�#��JEtJ��HK���E�j~�
�
�[�_K-$��	��9��0]h=�������gK�!��h;�	~�-}������@�5biVgVd!*P���#ZC�	���,��T�Gƹu\�x�/>���,M}2�P�, ��a¡H�������\y�Y>V
χb��(��������������V7,{�	��C�a�|79:���&C��KH�$=���Y�Օ[[�%�zPenr�2�'�*�w�8� �+h�^��?���z�<�Ã�|� �D��Ve���3�cV�Q֣��KA@إ�;ęVRB�1�Jn�3aM��4���B����z�&�U&�柂� �4 �㓋sl��p�6R :�>My��#/�q �z^	��v\GO�U�������3�]���b5�hQ^��6R9]A����=����B��hqn��\��*�gam��i䭏�"��1�z�*���Cq-��Z��;ԛ�]O��3���:������]yLN��8��DHؒ)�1��B�l���`�]�o8�[#@�e������jW�W]�]�۹��B�B'����!d;���q���m�m�«p��ާ��,��fo��׿�ձ<�HIP%�0���)0�g�=M�
GXg,��u��/6�D�\�tJ������S�g�%��e���oyss��ŏ`Y����^�@<�d_лW���]]�t�{=�]Y(p���C�\��cAl��	l�7��>�S��N|�H��!/S��>YɆ�q�w�&~��������*�}/v ,��/��S� /�V�Q��4{���A��غ�z�_/��az݆�9�T���a�$}�P��q���a�D�����o����*\SD� nr�茡�0-�!���C\S�b�	�Y=y���I�O��94LAR�Gd�4\���nz:h���{�7PI�aS�B4X����s�|�A���ڣ�<����,+N>DPH���#��=G��� �B��r��Ŗ�B���x$SN~����5�|
1��Q���*�<Į�3�J#ݯ�I�nOC!��K��D�TW�,}��v,W��5��#��/�t��~$�z�O�J�'ۏٖ��s�93Rd8���h>��n���S���E��Z%*m����)oڐ�-\.�e|/��1p�As(Z��u�ٝ��x`���������]���oZY���j�k�[ K ϋ���n[����6�<�gN�ꣽ�6��XW r��]Y�
ܿ�`�zsϮȔ�$ݿlv1�Ȼ���� �T�H�e�xە��������8E
�h�j)�Wy�6Z��}��f���g�v����('���B�uȎ�~�(o��F'�� ��@��#�-�|ZQT�X�!������X�1���\R(~°c5����e�Z���K�~,O��{}��U�yb�Z��٣��eÏ�nZ���`+����Z�.�'�r ��B2&i��#wk0
9�H��asN��)����/U2T�m#A��BMgɗ>Sn��R�U.޹�\ߋ72
v������G$(%�O��AN�A{(����6x,�l�#i=��c"�$�B8rT�wb��l��~��ƪ��M��HQK�F�i� ���^W��,�sl�#i�~B'nm���pϜ<<�}�8\�����!r��Ϩ}Q]D)�#�������-��V�v26�D�t8B Skv��n.�z�[��˨��C(G�eMq��X%���\Қ�%P7�;�� m�6$�ыV���H�������3P��9j�/�K)xp�ЄΙ��<���7�U[����)�T����r�]0s��B��ܸ�D#*�A!�f�1n�1H�J� S�/u`�n��ku�&���d��kk�bX��kO)&9��?�=J�;�:���}с�
�ݸ�5�@=:���L~|���.G @�J˨�-.�*��uG�_�$�i�T� ��l5�� ��(���H� �?�+(�V/�~L���ɱ�PPmF}V�嶋$�94>&��S$�u]-��]�YD�l��	�'��_9�+�`�)�9��*�`Z?nKg��\��-�b����&��������8�QyD[`�$m�žw��F�ŨU�3:�����2ĉl�u��aŰ��4k��t<Y!�S׶6��)�sK�c��g�O2w�b" w=�"�jrcȟ�u��D���"�v��7R��䠷���ga�VsY6~�T�|:j���K()}S�AE�SL�~��Z�r�g{֧������d"� ��x��������M�^8`H
Kŀ�7��!�;[��ph[J��k[J�J	��|��'k���9:�+ƅy
O��*l�S����d��R�����d�L@3�Y�_-yƞb�ڨ�mbAQmMg�; �H�DCϽ�ߋ�ҐD$��[��"�Dokj�]��i����J��xԖ��;Z.�˔W9�����=��@G@�K������AӴ�6�X`�J�L�R�%ߕ�]�d5�p�{PK?h9���v6��r2������,�f��+�m��hU�w^���v��ꉑҠ��q<���LX��Eu
��"8P	$si���c�ÄY��F&�ŏ�>f���y~�ƨ�uG�y��1�ݜ�N�!p=8�AXY���vXL�)��u�S�FR�|6�u'1��L���7�0~��N��#uƒCW!�G�i?,j(D���[Fiΐ�ͻ��w���h��f▞�M����oC���2���ɝ��:)	�k��f�A��9\i"�j�-K�,Q��\B����.�EyE� �?�Y�o7b���Ry% �Kp�ܶ�� :a��`G��-j�U,zmu�7-�x}�_È��i�P�8�V���$�̥�ݚy��|�
�oF*.���.�O3l&SŌU��A1��OlDv��0�.m��k+��l���n�7F�zD��w`Jߵ��gƳ�[l��hf�odl���K�*ؙ�O�)RA�
O��V� �I���pO� �ѐA��گw4m�vX]�;���|$��LjzO��vD$ء��H���Y�a#c��cRߗ��i�G�@�$�!�o;�/U�� Í����O{��ʞ�*����o /����Ea0d�5v��rԓ���! `���hWގ��a�[J�� kw�ð��XU펷H�˰|!cb�%ӵ~�R�7ϓP�tI.ϓ/�&����z(q��-��V���rsS��v�G��M����(P'=ž��`�x����4��Zm!�w\���T�]�TŊp�{��v��8��y��W�1�
f�����\�0���`�)D�pn�l�S���y����x��G0�|��C�6�z��
A���k�Fࣂ`#	]^��|;��)1;�߼�J9��T�` Z�
t ꞺQ~
��
�S2�w"A�GC?|I���nu�^�e�X��^�K�Y���>��eB
D�0��l��G�B����
�a&r�ж�}���%�9*KL��(s�+�|P������j"al���Q�G��E<�V@7�9Z"�o�Ԁտo�ݚ$���/<z���p��)��7���Py�����C�ؙ�
��I��V�y�� �Mz5Z:�ڐj�W��l�3ĳ7��
`����K��"5�H��B@����O����/����d�G��cMl�$0Q#��������������
2!���m��𣠋vl�.-%��B{4(��'ġ{؅��2�T�5	I����RC�[�n�	�"��4;�\z	M�D�f�9 u�c��B��db�5��}j"�g����{TT��Q�x&��
�>�~该�<[�)ʴ{R�Нq��9�X�r��v�*b�\-k�X����@�4�wlfm}J�#�K��9�t�b]����O��]�qS�r�Ju��;緻�E�3��b�S��̛a)E�b@���k���r��&d5T�%�;`�thM�$�[��7�2�+�����g���D� �_G��w ֎F*����S
�C�vY�v���r����]ъ��ʳ^�W8�A�Xb���K"��ૡp�`�fY$�F	L�m�(���#�AJ 9S��[c8!n-ԕG� ׈yq�o��r�l�I�H��^B<������!,�y�)#Y���»�`�W�v2�����9;'k����� r}�J}���g���`��C_X1^�FO��Fe��q�~8	�q��7�(v����oc���܊���Z]�f�oW��Tk������p6;�d���-����f��x�;������#��I���<.�m�|j��-�W@���/6��O�׏]��<(���0e����$&� �1��a�5�������h����L�]�����m���f��{+��?$
����d�g�gs��Ï�)�ӥ�_~i��[R�Wsح��C2�5ʼ��n��k������Se`@���ڑ�a��h5ޜl\	�&b ��/x��e/hG7��v�$k�9
�;3��3[��Lz=��^��ii��@o��Z}��>�W�TԖ� ,����g�@�{Xw��p���[	Oy������1*���ɒ��m��C���t�.&����t�>���J J	���i="5��I'Uz��[���$��m�2h���̀�\������=���!AI?�sAX���my�l-0���f2Ya=�!��5���
�L���GH-���~ \��
���J6��i��L`�&N���E�В��%1�̖��й���8j|Sn_yz�1ī�O̖�B�tc�M�iz��b}��d�؈(���f4���b$-�d���/� QR9`�LBSlӼ+3�m�Th�#|,�f��ɾK`�s�ֆK݆���.�.d!v"��<^�����EQ4�F�.����ɀ2�9��
h��A\Mx��P{�����(:`g���|]�pxV~ ��d����� �w��q�
�h��j�R�Kq�a�~����C��qd��ň�>�/�b�������q	d��wr*��C������O_Kh'
�4��Ҏ���Tք��^��f�d��x�✏��;��9RXSOe�L55�>J�_
�5���amo������z#�R/1u�~�̅f��D���Ϗ����q�a�q�(bb�����j��,\̇}h�O:>�@�P��6~�X\R�h�?b"���h�{�"��(o�♃���M{_�n�]�؀�F��j}�*��Q(��7����#�ʩ�g|�@��08g(��YS�(*}'��]J��k�e�_����]e�X)�-��z.'J����`NMyRC�a+�y�\B;��a5��3Rw�3I�\��t翫al�S�c��B�)�~]m��GO��dU2���9�j�`�u�Ew!V�B�� �c�,�����v��y8d��q\
�}q�]�vp�d${iqEL�2(�}��Maҏ�S�ϯ�&smz����<��N��9�_��a���t�m%ݽ#�X�����7��m�r���X�f �n��=7|����� ��E~�.:��"%��U��Ϟ��������3 �z�ULm+��s� �,J���x�ֿqw�"�ܯ�_é4�JKn��ilC������JI��t�,֤m.7�]ʬ����T�Zo�$cn�7Hх���7�L8���TY�W�:B`�Y!o��Ƹ�Co���h�9:�{"�«�:�����մӰ�����c�0�]Z��鿇E$�L](�2X�l�F0��Q��>���._�.iAz-��+�h�L�{�_�s�Ud��U;řA�O�����?׃��{ ��$:^������?��/L"���J����./Fx�ta����Լ�D�������J��ӎ�9g�f���� 6"!Gn/����쏢u�HȚ8!�^��|>(@��B�x������uj~S8#�I
��t0ƞ��X��v�������Q=>�a�;���b�{)�����6$�A!v^C�
�!��%	�/�%m��Sʸڛ�1>�^�鴷8ps���1����\v������K�闳,{tG�zx�q�G�=ɑ��c��cvXH˨Q`��p�o|x�TeY"��z�;��|1�2[�n��@*>�0�"�s� x:�D�������Х��9z��.�������N X����/�n܄����C���Y/��-<���kᐢ5����
11��1r"e��K�{��f����/�US]��6�dnP3�\��y	ST~�<�39�;�^q#^`�Y���2��H gG�xQ-�>@���a�ً+d���ʰ"k�T'vQ���kjq̵N�����7 ��n�V^�L��F��˵�#�:�'��TLF�FG��V(s<WpS��Ёq9r!�M�q�K���`�/^L`��w��-g��F�a�Q+(�a��*^m8��\�n�G�����Ù���	��U^R��%?��� 5%[M��S�f>��N�q�j�\Z�!~�˻�����N�ga��7܎
�X�_�Ǉ��6<�y��T̿���$���R�{�[oLl��:A��u�>s-f�:p2��D|$���L��A�P$Ued�ꖖ�И���0�l���冖-YU+G(eQ_v�wȬY��|��O���Jx���L�U�;s���b�ҭʞɾSL�mR�ʗ���=}B��F!9��t1�~�w��� ��C%4�^sٝK��� �:���_�{4���o)ɑP�jrd�͎oyn��6���iN�{��z��c,D�Ǩ1Gn�x�Q����@G�׫���m5�'xg&L�'�}��{]�L�U��a���Ȫnơx�xc�ǎe�o���ZY}�s�ɣ<H�]",�(x["����
Q��<FleA}�-:+���qu��6�Btw�pL�q���2�������{����
��&H*��E�s�kھ-D�ޛ)h���W���:�#�B�q&s�{G��ެ����T�]w��$A�H�D.�$�TQ�M�o�����+�����q�����ei����AoŐ�S�7�l�l�	�_��L:�C>e��l��;�L����ۂjb�~�/6I�u��4��aJ2$�v[
��v�磓k)o8ܐ�I{�W�pe�-�l?���!l\�XD�e�&NB	�V�=���,Mo��P�/��!E�(AP2��Цkb�	CIX��D�Y�V5����0y|Çt�2�=�i`�B�PqZR�_j�YW?ɍ8� ($	^@B ܳ���IE��X��s[>~Ob������kLf���5gt�*m�Wr�0@|���� ou��bzA؁B�& �JyV��4D�Пe���;�1��R����R�̉�<�"3�{�d����71��G�>G��<<�@�Y9Gۛ��/^���ܟ�ڵ&����'UՖ���_	h�Z#}]3G&e3'�F��a !^�Q�fP�����
��R|�e��Nz)�nƣv�:_\�p#�� ��c�����Zv�}�i6E�0$R�јL�vh��n�����^Ӂ���+�׆+"?a�p�5(�oL��
Z��g�g֑�D���O�,U�zy�;Wg%R�����tvow���ش���)s6�]��2@�%=bk��*0��Ɉ|XA���^�J������&��m�Y�fMU_F�3���o;�pL[���ab���y��<3��C����ꖟ*H�*�Q�Im ��'�K?��@:� {)�P}�{�K�fR�R�4Ƿَ�C�e;3��۶"µ�O�:П>�e����M��A��JL��_�)�r���)��e�:�N&�҄R����h���SӅ�K�y�3Y��
�H�8Ȕ�vaB,e��fݡu=1XC����H�ÕW�CJ�#8?p#Xp#h]&�><J��<s���<J2Mϡ%9�������{�ʘ�[9��/�g��N�N�yoܪ6~�t� �E&H�*!�8����{ʝ��j&��G��K����G�_��:�:O;ڳ�m����a_h�E�z={kޓ�7��z�b�Fz��zB�/�8N�yg�-���A�a��(�0�#�]���w1�j�cٺvVs��#��.1;4�(;j��qoy�<-���_�09�׷g[(KAZs��&�?�����
����[��pSW7=�m���Bx���`�H��r[���<p�7��E�=�"�k��s�Ic��`�/8�����:��5_H�Ɨ��J�p����������#`_��}�~T��s���s��7���w����x};�{�f���͵J{���Xs��r]T0(��w��i�*1�%h�{N���%:c�׽p�6R�]^�9�zNQm���u�'�EP>�6��.�	��I.��7�AR�Y^B%������}�J��Nv����́���I`W��V�/GJ��_��e}�_�wq�i��}"\�<�@K<��4G��A��� �]E����N���"�h�,@ q�{ 3����A�aY��/��d���҇5bbgȹ�a���:,褶���a
��R<�dG�G 'J%�NX�6�Αx^�I�Z�=���L��t��?�^�t�#LbQ�j�(<鰞��R�"K�ņ��f��f�I���Ğ�il�.�Ap;��Ef d�\�k�A  ���\}�)��|���,[M�8�.�In}�ǒ����`���m���9�v�
�C> ��(- <��$���s�,_�	�p{?��%�t/5�4z/������wJ	u~P��(�2ۮ��vu���#60��C
�Ȳk��~uNhT��҂,0�}�N�λ2�K����.��O��pIT<V~���
b������q� I�p�<��	g���͒�I��]�8��f��$��7!0�mΜ7�׫Th�˾pWM�ΥA��z*��%�c��#�w��� ��W��Y�l�[���5�SE��%�~����Ǒ��O&.���-4]2M� D=�^zH3~K��ߐ����#M�E%5R�n�;���=����0t�8�g�i0$9,�5��;bD�X-��zZ3L�����sF��?@�@�$Y+`t��P����E�܂ʯ����!���ګ��/����u;�xP���@Ɖ�����'OtK��}�T�{~����Ói҄G�,?��W.�τ��돸��r��$�#���1[tU��@�b�w#��
9H�F�\����v��oL�q���h�C���^�o�1H�s(o<3�&��8P@<(�Ə`�X�t�3)���F`Yh��J�H�u�}��H�\�c��`��� [Zf��ׇ�w2L��\��e�� ��s����07������;��ۊ��V���^ld�zZ����&)�/�T����[30��@��i���ݾ:SF��W�Ac*F�z��}ڌ���ǘ��N�;�gl�k7`�h�T=����c���%���XHpS`w��+_e�[񪗵B��_;hY��h/�H�&\�oێ:u�:��;d�poI�hP[:��w�������#ɀ��,R�)9�O���[���H�ƭ�>�O�g|��/PÉ�[C�A��)���lb��߆�N���ī��}���m���;v�_��l��n�S�[�H�%$��N���%���n6%���࣎T�@g6������B�+�	��^���E}(��s�qI��u�Mx�z�h�t.��^���W�?�f�vg�1��,��颋x�j���ؾ%=�&�C&CPI�v�cQhH�]-�<R��^�dG���i&�Z�/�>�,���࣢2��j�����`7�����N�WR���L��(.m� �z�p=S�)�(6$���n*�7�����0i�o�8�j�_��g�3�ZԴ�!+��ɧj9*Q�5�Ln�<�b�W������5��Ð�`�Z񵚌A�TF��Kt�G��e�ȁ��Q�/(xB����?|��ţ�}��Th!W���T�˘.�U�Ic�@G1��=�tr��<@z9�������	T>^N���`�'�|��JG����>P�8�Ȥ�zskμn��ǰsNe�p�A|�yRYg��W�|�(:A^pFzhՋ�q�`�_�j�2�m��m����a ��"��q]\���[,���L�#�KYU&`]�
Hտ�j�$�[yY�եɇ��N,��b�@�w�!�����v�CHj�˻Z�.��f=Rq���˴��燊&4����T�#�b�y�ϲ���U�B����1�4R�Ix͙�?!���"�3��B){s���&�9��:�*7����,,rV�n�	�h�PɈb~	�p�,zC�&���R@�^;�NՓ&y���"JV�s�tD�i%- .#��&��B�n���Iw{
�(Χ++�Z?������� ��������-Ca��j! <{ml�	�I9��3�XA�H?w4}��Z<T85�Rx-���b��%��1!��NF�`�&#ģ�tR�_�I�]���u�� ={w�v��o�}O~�z١5\����:1�;w��(�gP;�����~����>͌yJ!�� ���������2�E+�Q��Ŗ̧/U�{G~�����������=k�ե����:_�e��H�͡ۛ^��f�0��E�d�3�)�T��Nd�E�8�gi6|f�z��+�.^}�Ol�5�{yh�4a`Ũ��s�+Eo�)p!x�����1w�n�+}7�����쾋�?�{�F$�<kz����HB:f���asdB\�]��l��n�9a��Ƀ;�O]���PM�����	FoG��}��2I��A�B�>��q�	��-m�<��Y>�m���-+���虱�C�Pq_�����h��;F�,��Omҿ�M��6�a$՚^u�_莖�I��@.|b��ܺ�?�T�p�3L�	�1<�'0���x1r�
#�9c��O��܏M�i�֋�C�n�Za�W�:�#�rB�Y��C1�Fok�5�H�	��E�,�����G���^C��H�P�$� �-��n�I���B��aX�H���ߥ鳲njL�����쟝�hD��dN�^pљ&�	��5ǣ�d��!e\G�_�[7��r��㛅���-��ޞԍ�@�'�$�l�s�j�G���Ȭ�/�j��j ���G��-.�.4��0��m��+�B��M��W,s��!0�{�{��p�-�]�{ۓ��
|c�q�Ol�R�����ߢ"w��b��&-����)�4�?���9d��&�hR��d�hV��?���=8�LE|��}��ŀiqq�J^��r�a �����*M��k�c����� ���,��
z�bb��0�]^�� ���d_Y�."�����0����۽/�������uHG��~���u�ɚ��p�t=P�m}�p�A Q�f���LS��VʀO*�_R���K�񿎧I�#y�K�kY�w}�kUb��,:T�X�:Օч�Uw���u����j8Z�o�60G<ͣ��c��W�˗dG�_�����7�����`*�� �
<����0�1Rvp��}��'��R�F�#���t���cI�/9�2���1�g�?c%Շ��N���v��*��_5Ѫ�����E�9��?̶��l�2�4�Ny�tr�5��+G} "�&�@��<�d����ih�yj�n��]�*�@'&�]R�	�uI/�4@�Vǡ����+KN���	/Ǘ�w�V�/O�:?O�g�k#OUF{-��mLO����8�q1���}pΑJ$����b���]B�*���ֳ�`��30i��Y�i��(��"/���ﭻ�P�����\L{�_o��6�#�������,N�\��ܺP��|�SA���V��'�Ga���i�7��-�lo.|F	�iwTIw���<�'jpȝ�8w^x�Eu�gǉ�.�`���l`,]
1iP�|p�I��oL�i��XZw"t�)z�Ø6��,���A^Ƈv��߽�Mϗ��=�7j�Y�A�>�t/�R*Zaƃ�J&����I�2%��co���s��8z/�W�OD}��5\���<�n��<\��_e���a~y��8p��?z�6��Q'&�6����%�hyZi4�U��w暆��K�i�I��)�U��� �B�W
]������nOX�_���0&�]	L��Pw����U\Eo���T���y��'�I�8��-��|�<��'�N�bS~�:������4)�|	��]/W/|X��[��u�&�f.�E�4J6x�x6d�ȋ��wY��W=���ٓ�[m��Ǻ�/���Pa��~�U+�vW_q7z����<�:�e
F���Dس����
-�4kF����R�8��p~��L�7t�ҕv[�#-өVRר��uY��f��W�a��#�Fl!��;h�3������}~�����;��=W���^T���U��1 4,zzJ,�\%鼵�=N &*�ܚ&DO�T%�!��?�}5����"���}��mj���G{UD�I��ErSTAĢ2D"�1�9}�����V�+�x��"��+�U��J,�`�}����l�M��з~�w	I@w�8M�S�+'������u���f��yg������"��i^��!K�C�'��M�{��"B?Ȯ)JO��K��7�X c=R�練����������3g�<_g{���i�OC���6;3��w���Q��&[��x
�]+�|��d�GR�6i��i��F.U0#1�!)1�����M��/��Hk�_g�~�IF���#�H:���9���mU)��l�ƑV����FkX=�(߇�u�Z[0XT�Wc���9OHpeGS&A�RO>*���6J@�D��I�^�T�~�O�F�7��s��[���������:����s�!���D�B�L���scBD^�ah��j�]���������܅�(8$���9>�\�ĺ��4���A������'���ޝ�G����d*��tq��nІ�(X���d�u��d�	df��l�Oe�/�{+��ҹF�(A�\��06�	d��"#Ø[n���Q�����d@�*���<$?�H�	(@t���@/����@��
�o�U�X��z��h��:%PrN�kX�}��L��:Q
G"�f�Y�L� W&m0��Τ��8���|g�2\Ŗ���>1U}\D���O�w�
�m�q�O�|�C�ۆ/�����Q�
����ssR9�S���s�`�IHM�2i{N��L�薫�V2�,�'�vz��v�S��)izi�	��L�oj��%l	|�DR��[��*�!�5=�h�vk��љ�!�w��$�i��+�����b�d�.QM��ߗ؆����WpCݜ������)��WL~�i�r}	ͲȌM>My�����hD�A�/�?M����D�.)�&/բف���\*߻fY�.�XI�A���е�(J�b�k��#�Q�R휹�K#g�8��}6F�X�	V��s+q�z�di�|��F�,���-�w����l\h�P`q*F�B�*-���y\֪�!v^"�;u
�ĩ�aK	)if�����z%�bQ?I3X2.`I�l�l��v�n�V6�y���E��mM��:,�R�ܵ��F�=O����>g����Zb�7GHn����!�j�����ן��.�ø�h�b�ψȯ������ӕe�K �Y�1�}eSxCb<9��K��j�C��LM������2�ȯ�����r��Nh��-(N�������ޗ�Ǐ�H�w����A֌�cb:��u˔���	U��9�2 �����4a����ЙXʦ��[D3W_"�<�*�At���
`X�"���$o�����3��#�.ę)�ǡ�a�Zmt�&��h�����Lm7�=à�@6��ͫ��E"Ƒ��Q�
dB�"�YNՕQ��0�.�s��X��D���x�����Zop5�n,D�,>o5���a)��Z}a����&	�=�l��_O��w��d��s����{JO�VY��'��:�JI�B7s�E_��)F4�j�����Y��G/�^wR�y�e(�Ty�/���ǡ�j5��6�^��(�u�;��[Zp�(��L�&�x��׼�_$EXH�m\����`�a�U�͔nlE9p�x�C�n�t�`���!�L1����T}u�9����(��l,�3�VnY<����h����A׮lX����N��]
�s�E,��R��a����:�ŦQ)�<@�L �6����H��8[��G�ge��A�l��QyY��o)�N��U-i�sS,8,�jz�����S`g��ًJ�eA�Dc�	6�T�D��6P�],��p9������mi�yQk�YvV�}qʳ�W)e@	󝜶�,�����6���O�Ņ������a�:~�ێ��s	Q�]PQ�o��(��f�+��A{68Z�_�4@���u����+A��e�B�~p4�^���N�4k̀��u`�se� �Å���X@�A7��i1"�fÆJ��뷃�]�������:0o/���klU]-W�R�Yi�����?����4��\�b�r�k{�zm�{A�3�'6��8�p֫�7E�7ǹ���bM+-=�hX�>u��cъ0gĝE�¡,UK%��a�/�6Ӣr��Xݵ�F>����|����)�ӑU=uM�X�<_c�Jl�0'*���$��m���R�.3��qY��¬ʰ��?�`	�9��J;A?h�[x4�Y]�[).}
 �ݧ��o��R��5=�z��<.���P��7��E�϶e<'�~�'Š���}���߄]~p�#w"n�=�B	�c0a��Y��+H�B��f��\�$�#q�>�;��|5�u��ӥ�:��q��n��϶^�(9u?u*�J��6e� 9Q�x�v,6�އ|�|�p �nvB�(��(\P���s�RvOD�h�JJ�/��E�S���L�p�i�W�Kz��l?���(&[E��?�ȫ[�������4�}ѻ$|en?�<�]��f7]W�M��V&�4��D��Rn_Ow����޳Z�gY+n��Y�F��\�x̅g���8�d��N:���~xn*,���H����*0dy���A�F3O�I�����qo����x:O�BS��5�� o�3�n~����Ԁa��Iw�R�Ny�:9ʪ�Kr_N�{*O��:'�SX�:ߡ��4�q_�G�ϫ��ݗʘ� 80g����J#�VS��L�X�wScR�i�W��L�bl�Q��&�ꩽ��qY$�Zl
pP��N2��y�L���V���*�'�}���ѱ�	%�����Z>�Q+/���S�0�� }5/5� ���1T��9�5�j����p�p�:�%Qk�+�3ܔ}ڰp?�7l¬�,x��p�n�;X�{h��_^m_����e�����\�O#��z��lb�D:�y��㜥��$�h��"�]��>��z��?�l�G�0���V���ٹ����τ���Z�����Zk�A�Ub5p�P3�8?Ȋ{O����O, ��|"�C��,O��S�)��$�|q#�����8�&�&R��=g��7kץ���&�ۚ� �+�Pe�3��p���h'�O�m�[��'�����z�[}�g�S7a���>��ǃ�P�R�Rt�	g?"�ۂβ��-7W��X�V4>��0��
����P z�i�g��NC� [/0 ��~�?�s�4�s�	L0��K��(E)���	��1���}����K�P�u:��#s�r���U���|�JE��C�5�5�p0�I�s�l�'�uƟ���u�@W �6�Qi���8GP1�0&�93c/�pZ�ͮP�g�)ꕮ�w�n��^�-�-i�Қ��@��^���әc\
 �.aF�,�5����6��c,$�C+vF����wu�~��j	D��oN��]3Xs?A�[�:s#��~����r�������o��c{^K��h$L��� ����y@��3�X�PM�jݎ�;�+Ԡ(�W���@�0�x�P6Z�L�A�/C��L�r���a�%��v!�%�t�"�D�VLXE�o��rr%dz��s�"Ig�ۤ�H�mT��# ͧ2M�,�z��
��A���ؾ�&ݬPg�w��mP�v�g7'av�W��noͽ����$��C�u��Y3����wu�:5&|� ��]�b7on׊)��%��-e/�y��T��P�΅�fڒ��=4ݽ�z��]#����(��pB!�Z!/>d�I�b�xG�<� �
C]���X�;�����`nc�{	X�V� ��f�}mr#c�ؒ��0��{�
K�׆���8&p��f�@���z7w6���"�t|,��h���. ���_Pea����=̯1���T� ��mdL��H�:/�(C�`�>�|>#��=�#�Q�6�bQSW|�$d9��xpԺ�0��2<���P,��Ƣ��H��������eR(0a��_��60�\ԋ�m�([HNm��S�9�ü�0m���󶇳� ����vC|P�*p�]��H-�7��Kezy}� �ҳ�P��9_�O���ŋH3���JII�����@�0�12�����jx���_�<�!>��t�u��^��ׇ�%���E�DĮ�,��5�2����M#�M�B�����/�x�$���00M�:𮁀7�'Q����
���W
r���5C�W�:/�P�E>��!�}׃���$�xn�x������*Q�텟x+�P����7���ʡ�5�>{Jkΐ�_ݜbC�NB�eiP@��-X^d����d���Ͽ� �yN=�CB6�Ө�.�=����$C?E!�F��O�ט��_���X���;����"4	��
�H�0���Qk0Ͱ�=��N
�.R�
l��8����q��b�1�
w��p��`o;$m���yyc�L<N��c�E��Zf>8@D���mO����6kCI![hS<y�^u�����d<Τ/ΰ�h��9̞*�?]��c�Q�/���m)@"�l��@�����������fY�`�'!y#i����m�h��:��6�Vn؅`��
%��I�U��
|ebۀ��̶�'������3���JN���6��}�'�O)�??�lq�3��E����Gu6�-��Da��}K߃�ҽ,�T�"l�M�y�'Đ�jmSV�5���t��������\�E�1킂�L�u�]��G�C#d�EW�:�\
�s��ӌ��	:�X�UZht�R�{�3=ڻ�p�#�;�hG�=�@�Лy?�H�]1Oxˠ�|���@��Ck�x����?_4	��2~s�s�^��C�"첪G�A��Х/)mJn�LS���d赻���U�z���Z���lk	e�kۿD iTf�E���h?��'j���ϥ��o.7:T������⣄����DM�u�:> �ط��%Jg�8v�ƫ}�Ţ=s�e ��ڒt̉Uב���5��A]����U����U;�3���՗��2D��R��X��y����F>zLq�(K}��d���@�|���%B��,2���V�+���'�mY(�����c ��,�]P(�74@�~(_��;���.8!���G~Ku�dWh��H���Edה�k6-�@�g���m��*�l��Si�4�R*k����s�iQ�sV �%�ŔDJL��{^0�?r��r���"�1(%�����߻������kxy��ĉ�}ReC�z�.-c�-��bF�o
�૰.M�#���������ɣ��>~-R���C��':9J*������q1ƽQ!zw*�r.rXʈ�VSK�+�Ju�v�:����]�HX�`% ��o��#��e�Ac���ǚ�*�W�mXǎ���"L�:���?�I8:����3�Op���E���k�3A��'����W��R f���mHj3 
-zg�m����E}��ɟ��[8��4��M_z*i(�]��f<qʦP���	�S�(d���?k
~c�X�wa��Eup��t����_�ҋ����D�e9-�rX:=�t�A��r��1�'��'���]a4�
ڱd��Zf׭�Ͻ���>8���Y����	��u܅�=�uw��qb׀wڛ�ٟ	�m�@]���jjWv6�D2����Y(?kh����jl�?��x8��վ��z8ʷu�\�s��Gt��d�4|��	!���HrTX�g�{S��ͭ�UxpڰӢH�fFM ���t��KO=,G�����5"�Azx����Li(���Bg��9�:s賊��n�)N�lp)�PUK��"������'�ي>�àɽ���ܮ�<��m�X�e6f]}�3�����G��o��hR)*��ViCHU�B�����b�=�՗U|��йC���O��s|�\$��+!��t��#�}��`�ǡ@��57��K�ϭ���[S��_�t�9�O��&�����
���U�p�O/O�5+�K�ʢ���%���q�՛�3�!ae�;��@@���˦�/�P	{�OWx�Q�@�sE�"[��A�������0h�~�%�ȈDw�L�T�L��Y4g.�,��*.;6)	~����Z�Y�R���8�u��/��b�۔kY���=�*q��&Y��Y���I���(��oϣb�h%�	a�C�g���{ʢ���ߧ�0y洼����AP��=��"'���w6�}��U�z��_����/p�?*X��*F��P�â����1c��[�%��fb�B�r�>�ܶ\��46p�u�"&f)K�{��J��� �L��%�5xb%�Hυ0�}��t���6����(i�ꈵ�b��I�2��2�OtCyc�^�t֏�N!��Z��!7��-S�.B�O��U����h��
?�T�)u�KEK�A���W`�M��kc��c E��2R��c�W@���ג-ʗ/��)NeĂ*�̽���Z��>Q��H�"���qO��q��8��e�R��4�v����v{Jw�$���)%a���������)� ����4��A.���ؿ#��t:VI@R��#��<Px��0�8��#��!OM�5��w��G �69n˦5��#�M��� (aՖ"�mM��О	�SCa�X� �&~������x�h��@��ڠl.U`��	&�YyM�G8�V�r?	�R�#L�Q
��m,���-܎�'ݚ�^�+�T�"j�D4ͦU�x�KyI��՝�{�DnT����޹�dW�PC�Iib����������Z:b�Tyh�u�_U�%�.�k�T�:�V:��=�p@�v1y�GS�z�����%l�2�+[;��j��1J�>��&s�k�x&�}E�ɽD�?oxX~����5L�7�!Þ9p���i~���D�p���"S�5�1l�������GH���K-Z/��,'��������Y�\��e;�UR:��z2o�-,<�A�E�S�\���ݐ�<����xsaŝ��"Y��;�"��8��������j#.`l��S8B���X% 4�>-wBZ/�W'4!k�r[�/��%��8�$����
;ע~,��#�(
	:�z�-���k�	�b���[�I��-.,�W�L�0⒐�{/��$-k(k��J��"��i$�C��B���`J\��@PJ�Rhi���>���*ms���0P^�"�+s*ǩ��R�:(�+e�c0�t��)�t$�E������sK>�ׄ��N�2�mC�͝��f�go�>?
Ol�I�2+�������rj���nj]QǲE����[	�v-M�N��>�a�v�T�_Ou�� +e����3Pٵ�0�����l����u@	���O7-��]�}c�i���ysU����"�-��Ssd^�Uڙ� �&px��E�1��U٣#�A��I����sѣ������v�7-�� &��gZΘg�H��U�s��/O�cu���_(^�J����տZ�VhV��j��	��g(A��k��ڛ(׼���DQ"wSH�R/Zf�����8��X��+����?H�r��������<OC���1Z��ɏ��=4.�]�,Z�Z�	]��y&�(#"Bcu$�L�L�6X`�#�H(%�2��n�n�aua�">��$��4[�$���![�`�`\싒Y�E��3������:�$k����Qn�2��$�n�^U >��"��ZW��0C�n�k3�?]�Ԩ��m*	1�]y�q5��VГړ����)d��T����V.��tIG [�:���bb�m"��X�{��I�d�IX�R���:e��_�mjo&���]�^o)�[�����B����@v�IHOȵ��GJ���u�Dkٲ�h������:`��Q@�T��x��
>��̘>�H!��NIn"̧�\���h�|@f�" {';�}�0����B\��4� k��iUS`��+S#�\)����^�B��?��U��D� ���Ja��o���,�Aï�Һ��#���'�m}F������ٽ�1�
�=�F�L���'2��[�$>E�=�fŇ]�3\��P8ӄW)���2������C�����a��},���rD��F$��E�'(�d�B#���l�!�Z���p�2J?�e[��ӠDm�	��9Qk��Q�S'eʖ�=*�ȫB黋���x�y�%���,h#�����rʸ�����v�^sH9@�(+lٌ��VB}eƲc��]�)������Gؼ����gs�zDc�N}�k����"���?A��BA���;���PQU4k/����$|M�9`zOE2����l��0̝�ֹ��Ѣ��,%E'p��;&��e�Q�hd	�bzb0�W�%^5��z�醮Z^k��~SZU���RQX�])��9l�[��L�S�~AT�r�n���=¾o�843��������rr�t�n�t.-ڞ>��g4���λ��-����P��g�ҹ��J�Z�܊ZM9�!}���~�l`D�_��͒�����:��d|b;&��9ir��x�=�R$�{P�E|�!�	��C�� 1F�����~���>��>��,BF�.�Nm��*!��U�%���Q�R��[���*�~��-�5�<�� [���U���Ś�$t���T�'���x���sf7qƲ��@�g�6���*DyA�MN�I�3bn�i"�^R�ߌ� � �;�s	�n��s\=C��n��(�`Gq	���k]+Iߙ�Q��;���N<�Ex�����(F��v̛���*��1�b�~[�=���)���,��g���_dghX�Q��0U������>���#�?����&iVt|�v���l:�U?�6�^�sKh�����PA[�u�nr�4Y�M���=� '�����2�,/���g�+5H��Cɫ��7D�fZ2�]�i���$6�X�"����g�+� ��S�z�y��v����Eo��.�t`�h���0�;݌�D(�tȸ��tb�w�Vy���*� ��m!��u���x���/�0.�#�h��^�~N
�؋E�x����{q��0X�»�?0C�3�u��^�ݘ��R��)r�ϥj ��;>��?#�8*���.��Q��_���nZ�)4t�A]�~Zn�n�b���Z�x��q��
)C.H�]�O(��Yl(�8�h���)�6���efv�X T�p�/��O������y�@�]Kfb������f��٢���������8���LlT��e������T��! n�@��w���Ҽ�Z��۞�zyE@p��K6N) �N�b=��3J۵��릢�Q�m��Y.��+�
3K�豿1oN�[�M"]���τ���8Z��-^K�2�}Oo�$��&��w���~M��֫ Yr�kU�`�~Cd��"�Q�J�O᪊���_3���JY$@#�S���=+�BĦ Y�n�Z��4�\��<l�7E�Z� u?�+pT��*9��oKj�%��4�YHf��-/w�m�V��Om$��|�4J�K`����3��W�#�ȳ����>���\,9��&!����*x~�Ki�Tڣ�t�?y��0G(��khZ}��o�s�l#[Z$���9�G?`#��T܍ޢq������xg����DMCY�``聁����V �8����m�&:�߯뭪X2�������]k�D ��{P�3�{�? �
���Ĭ�B����>��8r�E��F�C+qt��}ņ�1K_����%J�9��t�*@͊G��
�y���\�M�����C����A�N��4q^��6�#���J�V�.��H]��D�l�Z��眑.[����C�d�/f��б{�6m�����1�!�����e�U��sz�	��"ܚgx?��F엂�|��#�,S���ql��鯵#DMC"a�G�DK�f 4���8ޱޅ�w�|�����{�����'$��]�=��~��<b��
't;ZɈ��^�������X���+���g`�5��N�2�����4��pj�-�{Ќ�쑎�o]��kQ-�qz�[��.�� �C1�]�PPGq�Mt,F�#�5��/�L�r +�ڏm�e�~������ ���ɐ@������n��ek<Ѿ˅�gsYn�ED!0lS]��Jc���ﳖ8�P����ٟ�tZ�ٝ�h��|n���<���Z���O��x֥KFE��v�t4s�CDєN0�S
���[�����Nf�A3�<Gh�㩹�U.)�j��V�U�C��QZ0��ֿ�n�}M)���_���r#��!<�2n���{�uz��'��zڐ���'px���A�1�O�C�9�=@o�<ػ�>Ά�$'p,?�<V�W��_u�(�n�}�� �}��R>J�����R�!9�����b��ր�f� ��>�t�[�o[����>�0��]&���H$�&����_<V�ʼ���W;�Ȭ	�_^����Ў��k�4k��Ce�V�t�����a�t3����_| ��n�`���4�TȂH�J@J��ބ��ig�0�|����wk�u��8���XH
��z�Q/��fV�ܙKS��d����OxdhxHlO�zL(���*(�w��͛����A {�t'�������W�D���ߴ�CC��q��q�Pd
un�3��Ry8�#jڈy��
��G�R>��G�o���z� �u�؞��#��-�3#�^�n��"����r1Ƚ�zv��C�T��]y���ڽb,#���C�E���D6�0��KJ*^��J��מ��A
,�w����w����B�e��ZEW� y&��⺰$a�a�#��*���$ތD���(�K�T*C���q�#�0#�ZK�D*�Tl8l?$θZ����O��=���EY��f*�h�7�0r�Ԏ>�s�I���a���U T"��{���$�������֣*CUd"��l�s	���,�,N+y���N ��x�G��7b>G�4��g��y�2ѩQ�ͫm����K�< aP-���%M�}�֚�����=ؼߌ_�(��K���:�t+	�P̚����]#�6s�W��	���hH��~AU� �����z�����XS��˙L��B*�䈱��p\i�t���|w���`�5����
�������>��U�2�|�[��r�iS��u|jG%�U�<`#B2�h;�ty�[���Py��27{�d��te� bpl\�m.�n��܍��,8!��_A��{鐘�	>�f���|!J}6xdZ<�x.SOp���AL�`:z=�CX8���#o��y��~�4+�zB�	�X��P;��Ϊ�Tex���e��Х��r�P���?���w1�Ns�� 9��peH㲼v+�s_�f�S�}R��w�t���\ �9Ax1�V�?܄���c�p\	=��5�k*�-�Xq�(��8�)�
Ky�#����8�s W�4����A�
Q̲��
�]�>�E�r���:��٣Kf�\��[�o����"6��׶E2��ǋ��o�磌5	 �RP��IUퟛ���|�lTw`_���kd}X�U���k /r:�|��6��
9݊`�d�irIM�����uw�/�:�������ö�����l�ڙʞ��T�A�}���Da����8�1�LE��H��b:%y,�b�G���"ds�M��N�=�\�^;�D����
c݁TDGoٷݕ�Cg�%�Q��b�O�����ݼ�٤�������)���-�Je�`[#�4�$T�����������{��)-�
����g����f��~v���Y���Y�U�]J��Cn��ǩS?-�����,e�(b��;����H9 ��[��yW�lLڠ gs%EȤ��k\T׶�qc����Bd��I�#�g�NJ��Is7�I�k��d�U�%�`gJ��}�� ���)�WIF�⻂���M)Ɛ����r��r6����#�,`hI%N�x�h4��?��D���PG	4M9ʓ���8�@و��1�����̓�ļa̐�Pf�zw��	)��tĔv3�f'���\x0�LdN�OK��	��j�=�9�&���13B�|��@���X~S�a<�ht®ǻ]_��x<�/5߆�J׮l�Pz���N/��oZA�k�A����/�n>C�r������j�Z�g={���r�,��E'����+Z�>�.C�Aq�r�>;�1��89��\�ОJ��Am�3xv�!��a�)m�k2����<�N��|a�? ��䰑|�������G��c/О���]Y�n��l��a��`����|�²\�uN�M�P�|Je��nWt���ݰ�o��nє8U �#sc<�B��������,zG��,��s��ד��Ζ�!ĺ������<��:���k�*^��]#�8�DK�Z��t���d�]���5$�1ůȓ��cdp���z�j�H��з��+_�9��۟��&��&�Y<�[�M߶o�Fa��7�`Cy��,(�I��aT;�M����Γ
������E��_�%2jK�4]Y��Y���`���j�L���yRwF՗��S7MY�I��c���Y&�Tԗ�w�S=���y����!��:[K�h����7R��Ԋ��k�������c��t�o�擜�Z���Y�IץڴI����WҀu�Ve�!�V��Bۡ��K���쬸Q1KYml��*=�):֊^ �=H�.�����j�,7S;��K,���(��M%�E�_0�8Tr3$���6�;o3ݯ擊9�2��bɏ�a������������]pG������O����Q�;��@}��v��x�B<	VB%�˚?~o��an]x	��=qV���&���'�0!7� M�*�4@1����RwS}����{�rSg� �1k�t(o����sݒl��B_,��X`KG�h�U@�i���8����麣Xzu�i0�eD��^�";��*��_�X��g'����gX��q.8���^HV����:�wc�F���`�YZj|�W�\�¾�����c~)D@�2J�A�c�g�^C��p��H�����8��#R9HJ�Ge�������MsJj\Y.��~<d���<�>;�����F��/��Tŝt ���Ծ�;��0��a�.M�am7�������~�I�y󚕑�9�)�V�|��D��)�9�1���|N��	��|'-f���#"����S�7���
)���凣���G�s�e����Cп��ր�O̘�ܛ��D$Gc�8qaйz�Ab����8Ob���O���W}�삇��l�����}7~�*��Qϖ�<�G�5j˅�/��}��]T��vm� -�Ot��L�1K�}�[�J���QxD0�x7�]%���X�Q��gߥg�Oe�so�7p05�XB^��^�)â��)F3-͋�y,����H᝭nͽ��9(��.U�ˈ�dq����&9H����^}��$NѲ������'�U!L��D�v�[�	�~�*��3sa�@��HS�7��5�;*d1F[�,O�t����(�ɵ�/U0F�����'�;o�r�Z���'�����2����f���yU~|%#���D�Zdp�9n2v4���	_���ʹ�2����k��s�R/��_he��T���s�Q,���m���a��+�ռ;�p�B^I	r��E���@=�����G�p4u)^��O�T�Noq<&!���]�ik3v�w�u�ؠ2|��K�EY'�x�d�1e�ް�N+CS��TH�J4?:�O��l����L��0�+�\�9	�S^%ą�B�H�K/op��w��k�q�v_K��yt�fq�1�6��PV+�kHH�y@7����]���Q�.R�V����������4Rb�$�����{�U��%0@)7��+��
�������i�ǁ��ԥ�2x�[S-��<�[ H'ߗ�ɧ�!x*��GX:�P����eG��X���d��Ҧ�`�#R��������w�t��_|E9'*$���u��z��W�WA�����U�'�I*��%ԕ���c�������0��SΈ����]��È��ݺ���3浦Z�l@�o-�C�U7g�@��Yf0�r���()�-v#�:?�l,5�S�W��ܑ�֕w�'�
g��
X
_���\��=��D�ۈ6_��؍� �eQ���s�@#ƬQ�P�a���o^��e� �+���@��>/J36�$h���f:�6�o9R+�޲�-��xE&4�2OKё���Yh���`l� �}�W��WWy�?Y�fM�Nq�C��d@�v5��e�F5+���J�=�/�k�t$�<�C�Q^����x�|p_��׉��'��#���Ƒ8d��IT�3c�*CJ�-�MXeZ�b��ɏ��@���ƫ:�����YƂ}/b�aL��ay�qjn��1$���f�}f7-� ��}�癨>z��<pbn-��9l�:�)m�B�X�ir�q!u��'���*�,9,{H��5��2��o�[��]�2	$^�rmG�O��@I�A�,_��p@P�-����.�j��|����6�{�
�����Pݎ��ѣ��˻`3t
�C7:��t2}ݢn��F�=����z+c���ěuN$�U����K'���3,��UT�V�<.N_�&���B���dC60ڏJ(��퀄&���W_91pW���� ��E�~d�h/���Ϙ���ݭ���n��V]Μp���Z�`����	�B'f���g�����f7� �y��9vx�W\AA�`<���@��˼,Z�4�����{��a�m�A�t�A����u�F���v�{m��I
2'SG2���C�t�$�O��e?I`�ay�S�]���Aϒ䅀[m�<q�]���|22YRR)"���%
�$9��&^�CU�+S�稼K����]��_��>o����Mp�������v����Q<^�2����R�����5A��s��J��,�T[�����cN��,���e๟Axo����x~�����Қ�6|>U�����H��-jTS5a��5��k����k+�ƨ�W�|�񄉓GT
ADt����F�F{o[�	%Č��%Sޫ���]�+���[������_O�O������w�m�U7�׀rjs�#����7!�m����LO����U����v>e
#�i��=s�O︹��b2l���?�¤<̉A�>�Ps��I��|4KJb	��ѓ���q���q�+���A�h���N[�\�ٻ�Ĉ����
o/����O�{`��U<C
ޛ���"�٢�lt��^�..�[�u���WD���U�oR���ӊ���8?�}��ٛ��"�<��h�	őkst����D��^~;���C���.����
�9�5ŕ� ԁ񩟍J;�I::�݊×�I�Ƽr��7e'�ϼ�5��l�����x�\�z_{3ò�b�P���(Z0��1��a�#Y��7�O{�ſ<�-� ������i��6��� C���w��l��7N����ۙ�&5/��UG��_E�-����9�2��o_	&�nl��o�=n�G? �k��&��U
��ѣW�=U�n�AJ��u����Z��D��L�q�2����\�?R $9��g��Ke��_���.���ǷCG�?�B��YsO����ﾲph6��β}|���A�>f3��o��(so�:ʎG��b�[?!ؠY��")S0~s\6۷�>��=�\¦�X��p͙�Z��t��{�.4	jXga��ߐj�k(���OѿV�y��1T�&��[z�E��@L�	(�
�O/#'x}���b�������^?S���PM��?���R�Xm!�XV���-���]�ea����냐�Ӝ��ʶ�[��%Y�1��-f0�E� ��׀0Y.l�"�U=��h�(�ņ�qa�7@w��x���rIDO{�!��
 %�J�?�z�ϴX,A s��bi��0���(	�V�=R�U#^�S�C^m��
�>\�	33
pn����?�cZo\�e�Bz�r~	�*CU#�=��>�X����2_�Y	U�{�y�~�.��}H�0h�@�R�,����jT���('�I���(�M�/���uY���~��
�S�J�q]�Րp�#�Ϋ�d�wk��n��2s!n\g�y{G	�5a�^#�|��9��I}W�pJETu���!�.�hY�g�fg�J�BA���;�އ A΄H=8w��ȒV�����\�z9����|�E�V�1�}�B?gQ����(��,�;-�MW���������aL����<��,�K]X��1�KH1�U���L7�Ǘ������w�!dG"�{J��mH�֛T_`p/��D��}NrĽ�ˉ���d6��v�Q�jұ3���b�%�q��[kCp5$��_v2�>�\�Z��ѐ��q����RTT
���ھ�hZ^�j���S�G�l��Qx�#��W���l�=r*f����8D��Z����6�<��9(�N��ѵ�w�\"�T��a�}ű�j��h�>
NB�S�*��U�★��x�^Cƕ�#�:��3;���V��J"�rx�_D?|0uvE��?nV@��r��e���8��y��?������Q+����:Ŕ��[�R���_����	з_��2��Pk�T�Qw�~	5����]m��^8G���|H�΍�hrO�HE��E7�/�\f����1H�ڇ2�^eRo�֮ θF����d��u���R����ߡ�!'��r��r�����]-��d�	���R'�C�?8�񼰢�{������^�|�)�E�G��!�ō��F�2����� �:/�q��n���K f�FwS�4�ŀ��=x�~�~Ѝ�pԫ��E�#Gф�q�juc��Qv��' �Ao�{ R_+K�K��)��O*b��s�1���L�ob�h$�W����`'U�A[�nܿ}�����x��t�V��g����J/OF����y�RA�'Br3�/��e|��Z�/>����dțD���괠9谴�mD���޳�%��1�d�P/A���'{jZ,}9��U�I������ߣ~��T��S�.�c5�~�[JR��n�)d�������C��`��[.�SK�Cű�Hu�
���� 3?d��NB��,gtP+E g._�*Hÿ$��e�&?O�Q2kU[��
w�W�"?P*�x�;u�
��
��O?كR�E(���.i�ҷ~��}����k:knjq�Y����*#���=�Kl������2#��q�^!P�I��[��GQ,�|l�^P���z�#P�˥qd��!��L��y�x�}<�;�����2�%����ji(ҷuA�=^$$!u{x�9��P�G}���!� ��P��A�gK�"y��E�ⅺ�隇y�K53�wN*f4�)2����ʧ2	�r��KI�k�.�>TA�jd�:m��"���ဂ�<q�l2��_���I�v�wO�M5���b��
��k��+��u�`�?,rn��G
@���(bR0\G�Ꭶ��dˢR�xD���"r�0�A�'S#��LT��m�[��g�O�w0d��RC����66���KS��֘D)�se���2 A���]Ӛ�^���.����o(�S�@>�(��C&��o�3�$o�%��?��M�3]Y�����?pZ��9+�u��k�?��_��x��!�X8��A��	���Z��x��e��c��7�f�"y���v����G��Z���tԟi�N>�W�\v�m����[����ܲu�4����
�?�������$�ñ��SG��8�5De��/<,�W.�y��Lq��v���2Z��������YxZaj�@܊��#����=%w�5�R�B����.�G��v���8�|��ه�(9�ޙ��(�>5G}���V ��i��𺥹y.8����*º��MM�֯.K������j�RG�ٜY����E��Ox��3ץ%4���:�%a� i���H��$<=��k3g�<�ßs�-o��m'n�=J<`^Q�y�x��	B3�s1��/��/BJ	oJӷ��
���I#6l�г}[E��oYY#fw���ז"o�0�֌,l�@F���!�� ����G�3�^��(�Jqn�s�
�Jy&}��6;�l�"�Aߎ�zz���qr�,5 Iُ��%;�<�U�\�)=}M�H��Uj�q�r������䓶o�nծo���2�����K`�~��)iC�?���#;��0'��L������>�Ѽ��R�����V�����4�+	D���xB���u���F�B�̃0ߝ�/���L���P/���T���XS綂'��|�ח���!x���y�uDB�a�gy��?���
�"�w��ߠJ~�7������/����lM��q�-J���C�d5�ǘ�PN�F�<tO�w^�K&h������W ������_P�sL}t�ط����s ��U�M����l���]�D;͍�E���G�jƷ�#�{w7g��n�8A�5�L����}����5�lR���7d�$hfi��	��.a6|´b�;��N� EI��x'fz�&���UE�Q��� �)!�&*6^E����M��0J�0��Àlj���m�k�)�~�~��߄^�W"��_���M��Qj`vϿ��4��m`�[!�j�e	�1�����k� �.��t��Q�B���`=!/�D��\���Д.�F.�cz8^�_�j 2��,7jTV���P��Ss�������It����~ܝ��%xM'-�[��j>gZd�a�R'1��v�O�yo'�3�~�_{��|-��W��`�t\�%i!��I��t�o��\ߠ0l�C�5M���t���#5S{�W,	�R�����m�`�ì-1�nCp�]�0�Kn���<�2�SN�}<<�Ϯ����Q�ÛȈd)�$3� M9�}t���S��qq&�Nr�&58�_�ä��6*��C�`��!ܐ�%b֠2`���
�]����s�����ښ��I�i!K%{�����{����.���P�	� �,�O��:�c�L�KL�]�@���\l���2�,��7eg�`��hn���OΈ�r�A����|���KOM�!�&!�3�
�.� C�{��ɀ]�V�I *�m���q���b�M�'�Tp_��N�;k�=2�O���G}�Ő-b��d��Ǥ	��q� %�F�4��*s>����G"��P�^��@'�;ݑ�� �����N<$x读R�c=!����$:�0!��PFv([(�O��"4p�c�!Yi�* F��$�.Ap�F��3�����r�dO=��fF��/)9%�JԻr��6��<3(ϖ��8�@��Ni��v�N����d@kh����,��-�{���:�3֞���R~{5��ӿXaJ����=�/�jXM ���U'�*C㨈��N��e	���s��\	��w!warA�CD��p��ֳ��s��2=�y�~�`s�зْiX�#��c������s���b&���d�/)$���3B(I'���d;�㕻���t�H�!q��ӐA��6	��H4K�ǃf����[׶��8��t��2x0��ʍ�pڞ��#�4p�S�!�Fw\�o}C�����/E���l���uu���n� �U����0�O��.����wR�1�i�0��a�!bN.X�g���7x��Y�;{��ʽA�[��E��p?���p���N��i�l�S@$I����K`��t�맗�܆��k����_�/��i�`A��g!y4�Eۨ���p$���D�$<�|Ox-l���I�˲�
����O����xG�򚅒�6���0N�|^ki�����	de�r��ebk�@�:eQ�P��`S��Ѓ��h��n�Mݳ�i{����k�}�~�y���!�ldb�O|(�([��hm��Vq%�a� ��ZP������)�V)G�<�),2	Y@x��p���|��̶�>�}%��3*=���
��h����L-�)��1H���ch 3D���~��&/~@� x����
J_u�_�>�w�v�a0G���1D�4O+y�d����"檑#���ע�FJ
� :��AI�0�t�{n[���}f���ud�s��h���@��ЭC�&�.�2i'{6��`DZ�y��&1EQ=//@�v�����n�p�Sw#U���g���g?���c��%��wM�6� l��Y�����莈���/]gL#��Q��16�+�\�g9�+� �f�o|#��t��	�L�&�&㼽C��Y���p�
S/�{Av{��zw�㲜v��ʶ�z��MP���
�r����<-} �����jdQ���r~�6��&��Xx���':�	�{Xqp��ΨZ!At�7��aE޾3_8��{�9-������[[�Yf���_W����L��=�'p�j�<��qhH�I�fAf���'�-¯~�&���z�S'���@���D��Cɖ&e��*U��~�l_����JΎ�W0�X�J�����1�5",lc}�
�����<Bv^Y/�?�=}�HTk:�y��J~�+�F3m)��!G�0�q�J�l��r�n�X�n��_��=����'����
'�3����XS����X��J��y-?�����+'oj�/0k����P*VR�ں�H��w&��Xp��%(eg\��Җ�]F��k��LgeO
���?���n�"�If)������l���0F��K8���N���.��XU(2H�zrz[c�5(��,�j8��l|�LYL�,�+�_��Bn"�Qr�෉,0��5J�ċ8���� ��r!1o���)���m,ȫ#7�!+,UT�G��,fӚ�X�-���[t����EC�RLcg�=Y���M��ȗW1��U� ���D�)Ъ~;#���<��eǈɉD�dJ��p.�h)�Q�q,�s�?b��}I�YWR�s2��Ќ&Z��h{Pښ��Q�2����.�=��j`��Y�D�9��(\�>7_Xo��~�A�l�W+*�K�,H[iz�0�-qw���퀕��^[�c�����{������n���w����Ә~E��r,�R��&c��!�*pf+��3%���`6W~���Y2%>��˞��#��&g�;�d�y{�}�\No����3O���z 3��l�R��к;	��{bl��Hv1e=DK��r��(#(���O!�N�-���ͣ_�&����\��G��i]�H��PơS�oH�N8��_�����h�}"�wX _��@�[��wf��m�A>A3e�1y<�90���H�|��̘�M�u��<�IF��Qo6�u��N__f0�r8������N��PPUP�y��y�a�Z��-�qڦ�1�4����l6g�Kf��5q��}޿`�x�1�d��LX�̩�� k�Or�����f~�uN��sx����[*�ߝ��7[��Ա�7<O�<t��������Kxo�+xSX��QS�i�b���d��*��Ї� ���zL�y�;�#��b�Jo3�!Y�����5����t���"����NұM�g�Ҵ.�C��������hB�:6U��P9,��ʲ:�q��J��p����%���tE�6qQ9�����C�kfY�LC���U�.wD�#R�Z�C��/i`�c���b����Q�����NP7F*RlL$��Er{�(iۓ�;�I�Q"}Q���)�d���+n6dl[~�KB1��L�8�(�z/@XP�_��1�*���΀��'6u�JK=�$
|@�
�-؉y}��yA^A��psbQ��g���cC��[�.�����j����	}���6 ~Z��X��]�ꪉ��"ە_�8ڈ�v�O�N��*vt�&Դkd~�^�]:��o�����n������"AN/��Z����(��[rS:dT펽��z׹��Z<��~��O˃���'t+�'���@I�B\J���(]���F/0�Mſ���ʉj��8���XB�,d��{�ة�r���H'h�˝���n;�-GV�q�ZHk¹��	9��3��F��R��^C�*��T�ʮv�!pOZ����b$������D�rS����.5ō�$zO�1<`��t�I9��
���.*�������:��QWc���W7c ]9��A/8���\u[�ڨd�����`�#�h�z/(��\�C�a�v�A��ʝ�?���#H��(��=I�OGb.��C��I��t�8xK���Q���`��(�W�Z�Ҥ��r�[�_z�`=���2���:�AZ�b	XJ3BL>fv\��yў�F��7���}�dɛ� ���L;�;�X��bٖ ^��y��}á��|.�g�J�ofRٻ�@[yu����`��Z��6
�GyT �u��ﯓ1�zQ�L˜�~Ch���r߷cIc�I^����MeI1�ʤBX1��L�iF�&RU��?(����ZȎ'�H����Ez�"�uTE�:h���s�Õna)%Rp'>��h�H_Hp�w�"�䷸��:���R}�z��Sm��I�]lƤPjc���;,$��@Vs�&Rq��9���b(��:�#�W���Ϡ���Y�n)�˂/�q�B,��u��R��1�ߔHF`��])#�)�@� lU7Ž;))�zlG3Fzuԃ���$؎�����I�U.�2I�Y*)��'� �I��I�-k�F��7���݈¾nt�%�	�_�/�2\��V�4H��P@���&�_| mv�I!\�>�7��10Z�k��5B���OpLKu��Q����Nra3|bx�C����=�N��$3�z�3���Icf*"�iC��s}�Xi�t`�Ͻ?��[����.���{�!zK}��;��n�f>�}�����D��&YJ�8�֑?d�$KW����:M�Aws�5�RxQ��[�i��_��QTV^�����x�d�� �8Z"�:0�r�l�Q�(��`�Zw�����5U|���+��pJ��1��,����ňuE}H��(��9XE��5l��5�a%��y��wU
����V?�f�,������H@.�^�ň�ǎ��U�j��r�Vh<�g��Ŋ��Aq�\
�)Q�&[�8�[2m�V~�#�.#�_�)4V��#�6�T���/�o�;�7ŏ3={CI�t�s��K��i�%� �t%�-}�%Ƚĺ�&C�=6�������:z�%�|7�S�~=k*"K�D c��d��oy�(����^�s�}�2)#�,����Q�]|g�C��]�|�w�������ΣNz[�K�h��CĈ����۩K���|IU�Zz$�C��/��K���"S;kk���Y���-H��dM9-�=A]��d�?35$�t�E4Q��_��2�#�,n+�v �1V�m&���=9�E~8o����9�xC�Y��3y����>�,.p�A#�R���7	�j-�����Uح����o�\��a
�59���j7��s�.����PG$?q���h�iY�_Zg!�S5S4*��P��Wqfo��BZ���=�A5�}f�"��@P=�{ro���+!߹�J�R_���g��MIGIƚd?���ӹR6�)M��� @9�j���x�B��{�`�����X�v[kFp~���2�����&/���U�L���h_<Of�����8Ѯ���Z��β��?���,�4j�3�OE�&��t�Y�Yچ�S�1�}:^�������	�R�_)YT�%*�i ����@nJ��8E���(*ȸ��#�;i�9Am����0�����(γxN���n'��{�������d�c�2��f�h�0�?�Ib�����O�l�ˡE�s�ح�*�Q��Yy�[j����1E4�3d���Q��'B>ϟ�땜�ñ^�\,�XV���諾�^��㲓0��`��w-�X*��]��l��1�ο�&i�������]�3�XS�Q�}�� 5�ȠR�+�kZ�){�<��(Ğ:*=�|O�d��)R��u�i��a�}{��x��tR�F�ܠM�6��nKPT�u�#J�ʫe��D��ݔf�F)X̖�H�%f���m�1)��DX &G��Ls�}U�|��`��p3�rGp�G �l�@�9�zP��� �C�-�� <��z�&+iKWTb�1�ƌ�`�!�1�i;N_㜟�0�5�W[�B�`2S�O�8�X����Dd�aЛ���d ��-����klF�!Z�2�aZ�x�v�@��n�=W�m�W2�3a�p:��K��e��@;P�m u���O�S�*�g�GfYM�����cV(�li��d���v�4TdǑ|��ߤ]+āDwS�`�и�����%��0o��USBk*r��Mvr�ٶ�$J����W.�y�A� Y햀�Hn������3.��u��Q���m�VXD�r�%Dt��N���'�.�beφ�4�}U�u7˞4�銱'�R�����}ĳ䩬��X�,��骒�H���F㑂%�1��u(2��IG��U�8mkPevN2+K�������Y@ީ�y��5��&jˣ�v h���Z�&	ZO�v�:�)p�nA�����?�Zh�����}����8���P
>o��V����F���a�/�OIA_ '�%p]�弅%]��D�h�d�*�	����S�hS&V��@�=jK���:�;�Gh?K�2-�
x���0���"u�'�sCX��h���2���9����ͣK,����r�o��/��J���B9����=6����!�PZ	�؉�������A1�(��^`�Y�VI�\"tgG�����Խ�n����-�M���^���n[�*=mk��-����ؾ�*����y�V�v���:U��W�o"X�z�j!����k�'H�zU�!Q�D���/Y�9�[�{�w�_�������!�����<��\�+��kVX�����5�$-e�d�n�J+�"=���:�\�;�#���C��H�Q���r%�ݍ�$�P��n�)� ��a����]������)�p^�m5���&H�@�C
s��pz$Ұo�X���m��|緕 �Pޕ� �z���]�7�ճf��bMG�{�t,BK5��I�*U��_��<�ܑ�%�O�;�[�z�J��.�=��H�𻜜�^HZ||�z��#8EѨ���Q[��}&� )g���(ڍ�!�0����Bw�#<Ҍ}~��'������K3s��1h�^�mv`j�u�����N#��w��/2K�d�g���$pQ�/P���}�	�xՓw���}�K�k'�CAA_T�h�L����[9n��e.�#�;I�M|�/��|��b�p��R�U�B��<̿j]:Wj�ȓ�o����-fQ@)�;DjwH#�$�ik�g�m\̴�ΧҢ��PC��<.���Pc��Z��u
�@�3���A�kR�������d��Mg�7�B����2�J���-*(0Udd����v}�>�7ڰ�VN_�qg�@|��b��)�����X'O���=�XE�����^Xxf �������E���G�O�fygL\ɷ|V�g�VH��S1�/�BM�|�O��#ﻆ*ɸS��j�_����P�����Xĝ��@6�Dy�f��������tˇ_N�XG��C#F>L*.��A2�P�|��05`�m5�ҡ�����c��$��9fp�G����Z�CI��6�9��CO�&����!�J="`b�k8�dzF"�2;m膝i�|�j��c�lµ&�Z�l����v� ��r�9�x7��Ӗ"��\I
d��F��pl
I��C�g��S����uX�z��q_���#��x��z�M5�KI������÷3��V�q��c}_{��R?p��]�w��HU����١������̼a�4R_.2��x�1{�0Z� ��g��jU�nl+&�_|U?�W0��"��������xJ����w؁@�����ZG��\���qR+O���,��K�1n��n!�WO;%����-Gb[�N6֔�a�� �4r��VdK�p,�ꅳlG�����T���9zO�l�ύ[��ح�e�O���Q�����z�V;W���JM[t��������<��� �
�d�Bd�ߣX�\�y���7VrN�������`�h`���:%��Fl@�v�w��	����;� � 3��0�	#��/&0g0%t�ja�p%���jR"�k[���q�!P�����35�+���=�2������c�l��_�ƀ!�{���+3Є���S���]�~�]��CW8���я��˟߬w\���z��Њ�B\�����1j������ G��h>��{r0�mU�må8�mmf�&�.;_Uu����h�5ћ�c'�Hx�T��N�o��r���zn��M�n��%u,�xM$����!�Z6�h�c�§,�� ���Y&��_��| RUl4�a�U3U�?2�7�~A[�W2�η9�B�W���ψ��������e$L|��_�G�2����`s��?�<�lta�����h��Il�Ə/��ʿ�{�@��k}���Q��먠p�棬�o��ez�D��]JK���)���8�)���V�\kl8���m.ѯ��];5����<a*���YP�B*vR=Е �Qr�Ή7��{p�2��U&2�fMk$ˇ�meB�@����	v��Z�Xh�X*<�%��}t?]��Y{͘�=pX�S��O�T��}�����ۂL�Ef��tՕɕ�:b�����#}j/EN&��h�w㼯�Tr�W��t����᥷��*)�"��*�f$�(�&֯�|�e>��~��L����_�0EH�d^�O��ۮB�'.��>�O��+_&����C@���L��|�/Q}�N���L3��̳J�
5��|���$�~��x��ؑD�k�{�]��,��fV��Z,�@v$b�G�cָ����'A'�D�r���٧��"W���� U�y%M/mJ�bi��<d��=�/�ER��$�#\�A.�2��ذ��[f=޵��V�1HM�����0~)��������O��%��hzm�WfM�R�u���P�9-J	'�~�������r{B�jΑ��$�x˱�\ꉢ΢8����L��ڵ��J����� ��Ku�U�e��W��nQ��P��v�Q���Ԏ��uf�N�|6{C	�X�)�k�4h��v���3�V��<p��g���6vF;E�o�P��}S!a�}-Q߲��Vl�B���x����r�r����s���B��f$�����Je��5����-J��ưr�B��a�͔�A
�zY��ô��81t��m���U���r[�I�q�i�\����(�I�� ��u �[�E<��;�t�Fs-.��{kBA�n܄�E�R�~(����V��g�$�F�z�mo��?�-������M�m�tD�7B�hf��8'A�c����yl��وP<�*���m�k����d/�j�<w��I�cݴ�kÁf'wvW8�z��n�l�1���1X}Z�L���x<Y@�1��&) ��K T�b�@K��6�Ƀ�r2�r�\��	�NtI�RJ(��'�p_̉=���ۧ�ݯc�ke�Y�9��2��̶:�=�f���&��D+	;w���d�I��E!
����r"�[K@8�-<7���vA*Be�N
@�'�q�p��U�d������㑆��ҜK�׾�#4'PJ�V��x���hJ��������T3A�CD��Mտޅ��u���EV�(0:Faw�+ [Ĵv�m�B���	?r2͇B&_�^/n%��^Ϊ3t|�%&B�x�Qy+hNҴ���V��� P�>͉\����$q^�*&�sk�+���@:M3���v��ûɛ��UD�?��<X���������D�)e�C���>�$�WH^�b���H � S�Iw�L�����]&��jq��,��H����C�����h�i��FGX���<>Ę��X5�-�2���m�e+��P��K ���<�,ak�kT��C!�x�����!�3䙦�4/-nN�l_lL�T���\Ir�@2W
n�$O��$�I��J�-�}�V�&}����]�dO:+�U�htgR����؏���Qb��7�Rc��U�FoP��Fȶ艓GD��a$ٱ�N����R:�i�ʘʼy�z�|ۻ�_�(J�a�������w���^x��]� ��!)�h#�\1H�S�v<]�fD�|	��֜����xЭ�f\F?nTN��{1S��1�9B�^�� �9<M�擰����*�>��?��Uc�Ae�znJ{�<�7�8-{�C�*+C! ������� ��������{vB��8<��f`�@��Z#`Qϋ��U��I�4oM�E�i��t:�E��Tǔ�H�.-]?>�������qW��w"���8�+���*GG ���1-�}w�m�:KgJK�i�+��?�_�5�w�EϷ����l�$Ӎ���n��=	���K���)Jl,��b�)�tFR���g61$�$l��Iǩ8,R�.��
�q$��v�不Ϧt�I��8�Z�SǑ7ע�iW�N��A�$�)$�\A� �ԭn7�)�K��b��\4u���=E�G����m�wꈾ����N�"1�t8ha��~_��W8����e�9n�s
�6��E�D��y�Ɣ��`d/�����O�H��p?2#\,�(��@�"�v�w��J�����]�e�Ћ����0f���@5�Mtu����~N�ڔ1��]qi� |��\� X�b�I��f�^�t���!͎�����F�uD)5����@�'y�L��(���G����ƃ�~��	j0!t� �k3a`����e=��T���llK�Ǜh�Di�̣J;A21���|:R�췘|��x���I��q#e�6��Ԭ�� o(�T�6�&X��*Rف���VJ��_k/x���Q��E���Th�]��k�6�>]K��k��A��#��_M�ܱ�f3P]��e�%��:B���ը7[ܵ\f3��7/���%���P� ��V�C'�C�R�vt�&w��<6ͽ}�у]�C�B_O�ozR���ml �R Zd& �P+ l���}r���U�`�q���cS�}�O�R���k�;/@z[�Fe�	����%�3�A�?�[8ୄdᆫg^���zOS@��N=��Y��&l1$����f���������!z�(��\�2y?�S�b��S�2�9{	C������Ytv_*��U�s^eGV��y԰	��1��a��k��c�S�v�q�'�Y?A�~�Z[���dG��2���E�����h^�!�"�_ZH�("Kv�R��#N�I�sА�N-�94�!.��I3o��,s�#��x���G���;�[��i;�=~#�i�,�U-�MA�2�5Bؾ���`N���%���%E�a&pK�*��R�&�)\�E$��-�Z�z�sb��4�p���@_Ba��ߵ��ag҂��e����f�#M����q�gƊax�4�z#���/t���(P	Zvf�+������	`�m6[��2���PKsڛ� �?o6Y�^�	��-&����(��wIno�2�>��l�)N&8�( 5�Z?����}}u�6�V&�)ž�ϟ�h�Acm�[����>%��vfԦy::|��F�#ߜ��
�4��,X�qpX%.'k�6��ie��r�T�t����8Hiܲ���Aղl%��y�lRIC%⠻h�1h�kB`}K/�l �)�_��i���t�A��pY'����*��l��9 /C���ʢM���
c�Fĺ��'T����݋q�.:������MW��:��G	!�^�#a�����Q)��B��c�)"�_�kƶ��P�=]�#��ޒ.?�47��J�X�mIW��wB����-����N��,j�!M5�̓-�)8Uc�p^�V�%(H��f���8������9,c{�me���7�Z����(˕��+������"3`^4c��e�)^��i��KY:�9�\|�iP�,�:����7z|� G�侌>ԄUԺ0�AD�%v�4m�5�-��3=sժ�k^�����5~�(�iT����[�W��s�~�T!���U%�0�g��[�s4+��Lg�鈚��K�jT5V�Đ�;��u�I�٤RA�B.d`^F��W�D�S5�j*[٪z���cO�mU�¡������G��v����N�����lY�����u�Ŗ������Z�MWz��>�0�F���y���]~�����r�ꏃ��6n�qq����¹��p����\*�i�pJ|	j|�α�������+���n���@3��*�������f:lX�/�h�W�#�1���wI��/ly�jq�*��֫T�>`�/�������܉ۆ�ַy#!?5l��C	�K�V��Ϸrn��A4��S�tB�BBbw-�!<W�N}EmI1�{�(vxL���6�Hg�l-��d��̫�ډ+'=�uPi�I�N��ˡ�6�2K�����	Nh*�ҷ/�3"7�8����8���i���m�E�d��>������#ζ7�L~�n����WN��$��j����T~#p�ם[/��G�
'15Q��c�T�2��5`�=���; (լҕ)�uO��Jp�^r�q{�K]tƴH엙����R[re��-'I�s�>1j���Y��L$�*�Cq]o�K�1(˰S�����:���P�����C��MD缰����|�����!� ���a���ʰB��VE�Ml+H�z\(7���ʒ!������,����Ls��7V
g�����vf\��+Bq��,������{E���Q�*�y7��{�����x���fw��(�C��Wۿ �(�ȕdǾt���f$O�� xt4���x[�$��HW�y 8L�\E.�W��N��$��L����Z�?v^;Jq�:��	����������9�JcW�W�L�%�Έ����H0�Q{h�Ux/���T��Y����+�9����:jD}��q����Q��E'+	�T��ome�D��i�1Ԕ���%�_GPy��M��!�D9���<���!�TyV��>�+k���M?:��Zp	n[����H�I?��G,����Z�kJ��o�e�*�+����E�d�Ŋ��ܓ�/�"���|n'�q�Zt�]ȾS�(�ρ����a(ag|���ˋAX�{������<"�H	����lOڞ�2F��������ؗ���f���5���gɔ1�[DU��M������c;��Bf3_�N���BEϗ��cT��<��^�6�6PƢaq�˵�(��jM&	�Y���!o�rz)ÝãH����4��K�ٞp��h�ޛr��]2 �V6�@E��IhҞ�<��y���i��B�	��*sQ0x^_c��*���I��"4��y�`*+B�*4i)^�Y +�è������D<�E/a|䖉�G�A2�5R�{M�ũW���!�V�`qlw�x\@����=��b�g�p��7P6�Y��r^b@{}��0l���.�g���I���'yB��~��oy
�?7��t�����eןh����7�x�K@��C2oD�I��A�$���7m^u�~��";��LV�7F�]��kV�a)J:�����D��ס,ג��gebx�k�ȣ/~W@aԽ{�=�l�#<l�cҿ�6�&꽅�ἝD�J6���L�̝�ӫ���l�vq;5�?�+���"��X�u�鋜+h��I�Mݏ� >��� �����=�F�6���ʊ���m��A�1��2��xo���*�?P�b�\4֎��^c���Oӭnj�J�5���Φnp8K�[�U��������Y�H'X��Ǳm-��1v=�ʄ�ڲ�>�mmOHDָ�R�a�.�u�I>El��@8]W��Wˏ#^�J�I~m����}��0&%&���:����r�$oƕ�6ͥ$
�UK�y������G�,�����[a���f3�� º������8U�s6}4�α1$��`!v�����'Y�і�&�����ёC�n*�~��c1�B��Y�ik\AZ��ElV�V���+�$y=i��]h�� �MH֦�e�gM\5	0�Zw��]�������x��
�x#�K�3>�Q��Q��N�9ԊuPh�=6���?1�4C4񧍢�֧�`)� 1��o%�Ƽkd&Dذ'�/P��?�T�ig��C��Q�qrt8�Dd�R�L���'n珴�`�Qt_.q.]�I!p��ؓNqi��+�>�2���(�	[��t��V�A�wJ'Oĺ�88;�׮_�u=!�Uxq�\��]�T'��\���.�X"E�$�ꕇF�J��X��@�\|q��"�p�e�s	����gC� X����bɐPp�����7v�9�� 蚎�=;k�\��r	L��u}4����Cd���)�V��'�q�R�
�Yh��U��i�,�WK�2�pS)�+F��
�?P������-�`�{�XX0����0�A 0��,T����54�oJ�-�e�'�*���k��`ϼƎ��]��n�8��}Gci�G�9�H.*�lr.�6�b�`�Q�_;D����{���f����T�fufM�e�<r���7��o8x����p�FY~���	�	]B�sVݮ.�_��ȓ$��B���OET��{BL��+!&/�I�ʆqUH�1���$�&P�9���'Գ)]����sb �/)ɳ�Qރ��d1VJ�%�>�^�T$E�a��%p��	a^�P�����;o(ur��Ef��-�X��#��fm#�F�˴�7I����&�Ƃ_�<|>D�-z�H�ܸM��@չ�`��/7W���1b�'dnr�������yO�����.'���~�ۿJ\]TO�j�+�����R� A���K�a��	�#�5U�(u��{�BR`�/C~�coC:8��b��_�.���*��	��v ���e��3�3K�ڬ.�z��lKx�T����:�f���7k�ἡuC����l��PĴe�B���1���qNNj��]h�BJ"��6D���']�3b�Z�
P���v.0�KE�cMg��W|~�:|��N�;4��G��^�,��tGyg�C��cť�~T?�[���u�	��(�%,�)���T�P)[R|�Y�"R���j�n����U��Ѩ���N�� ���x��2dm�][m3�@ Q=�?�5VD�Y���BoP������xy(��텸^k��`d�/��Y,&Hyf"�~�3V���u"������ٗCU��!��9w�N���n}��� �'��m���� ��-HY��5&��	�N��6����a��*�C|.�EI��#J�i�bn8��}�b��
�F�V)1�[O�͏�Z�m  �]�!O�`�E�K쨳x⁬�
��{,��N���ƭ/�^ �m�A�k
���}p��?��j��
%�Vw�ͤ
 �롮)����%�Q4X���'�%�D���t�㍎M�]�Uxe��w�u���C�6��Ğ��{>I	���Q�����"�{?�\�8j��nn̈/=G�krJ؆�6=�9�jĪ�C3������9s�3��L'�I��z�ʲ�E�rqL��������]ڕ\�47�o�$�[[�%��W��ӗ�|p+�j�Ψ�4��0l�h�f�dbPr�g��<H��ٻ&]�-$�a�6�
_w��H+2�ź�zMBk��]eV��,>����O1Y�`]U����c3墬�7
�ϰ���IH����]S�Ͼ�#��b"Pf$+�M!{��g�>�E�3�!V�-�!p�Q��D!jo���]�u������Y�$v]��q5C{��N�v�X\� m�{+$�b��Rdu��dĹT�����"Ҫ���WMl���%Z/�9�*2*6E��M8�Z�^�&�G3��;̙�1�0����A��$��f1��FHb��
�9�rB!��âfǡ�v�t��&̣��0���j@0ܰu�*�5��w��?��]af&��XP�lV�}��<�L"�4�	ݍZ�Ta�H�oq}q6�����o���~���[z/�
��*����wߋ/��V	�N��5��y���(�K	����輩+ Hr%��;�ep3_K_�v��,��wҰk�(�xbY$,&W$�����x����kz��a�����E�1�C����Ϸ2xMFX��X�/P�߅�9��52ʖ�P�D;֡�˸MJ���<%K�۟��_�E8m�f�Ǒ��ˁa!�0���%a1��d�ޝD�L� X?��q�\�E��zV���"���Ui��n�c�^Gm-�]�d�#")w|���?y(���*ʰ�q��'<ۮ�sF��"ɬ��H����5������eM��Z�+��d簈���Cc�EސCŧ ������(����NK���%��I�Z$�W�bJM�������c�jh̎��R�2�cI��%�[x�Dg����'/�$��A��SAW�{%�
,��;�!|]��uBi�b�X?ب��j�D�����Ý�y޹�/�7r����I���ކ3�=��nW���$9�	C҈�^٬#M�O�d�ST#�G\�~���b|QH�ύL�*_��s9[��R�P���a�:��=L�4��_�pb��kqt�/���q�t��#�S�:4�2s��%��;��x�w�k��jB�� ]�>b���7���	�i�"�=7KO�f6�F%Rg�`r<x�٫sेm�}�M-i����m�+u���þ�Rϒ�݅-�p�ޅ__e���uǂ�>$�ۗ˰�����"B�����]�RraXsc�\PP��YR���u�9�4H��Y��C�y�~!�C���@�������Sb[�2�A��1Jcε�5�n������ݩJř�Y���[�o4!�J�O�Q۰R"�p���u����=�P�6ӃE���(d�^N �J��w6{7�<�/��?b�1_���}D�e�x5���-$Qi[�Y�m"Ћ�(�B�k��D(e��͍h�裪42��pT���a-M�,��q톍S18t������Y���4ܞ&�j��[��8.������f����wfm��穕Zg�]�9U��u�J��b���7kq��3M\�Dn!6�V��^�M������?�z-1�k����\�ZD��|�y�5L��z�&M��ʺ
��b���g��.�§��o�Lr%�U a�����&kD�ߡ^��B�I��E�lM�UH�"��������Nw����'��=+�x�'���]���&�?�.�x(�OA}h�tYK\tV�%-X�\b1�A��l)"�m-X�H)%A,Ab�1�	�ƌ� 7"�O��K>X�2����	]74���-��e����B���PVl��8IB�&�M}$��>e��"�h��X-H���U���h��H�N=��D���[�<;W�ဎ�;��v妀��ro�QF�|�W��mJ){v��bK�9g{��� �bJ��z����l5B�D��E�� z��
$����� �^}�	��k@U����F����:0�0*3^�g(�t������uV�ҿ6�k�8��Q1k�z^3��
�W��:��4#��i��cbк���ε�/w��V"f��v�md��-"w>u�X��Q����t�ě�!��B��tVvB"�������Nh�T���M�z����E̓���@��� H��yB�NS �2f�P.-��^�)hS}Bf\�B��|�#&Ѕ��=��^��G�߶
U���f��+ʖc�H����:��)ѹ�$�RyA�Q6J�#"G��J42)�e9��d����Q�Ҩ�A�"�g �f���y��,��v4z�w�JX�9U�T�Ռ�މ�3]�.�FY�\�k<��x"G�͐����l!����ن8�XH[\�gw��9ŪN���1�����Q�e!f�~}DvI���Ǥw�q���o���ȟP(�ۚ�x\�����~�/�i�F_%��'�]�-�VE�5�������,�rӈ����{ z���p�ۺr����<ug�Mb�j�4oN!m(g���~s�xQ.�B2�}yP˸�|��64:����7��W*$(��D膎���㤪��NWX��i�L�"n�ՙ�/������Z�o ��ꭣ�6�'�4�'Sc��{Oy^A8"衊��Xt�r�[�}Th�6�\_^Fƕ�F9R�*�M�5��䜝uԁ����i�����v�J���k�q����~[��>n~�G�g���w��x��2ii!Ku�ę�&J���bSgs�/�4J	����@��g�O�a慅ܤ�Tf�_ˈ�:�]��f�?��~�r����]�DY>���a�:(�3��P��VU��tK�ښ�0�acp&r{�`~up/�:��T���գw�%��4�2�%Í_f��Q7<j2����焩q��@�M���D)��ńA�7o�z���0IuCBU��IG~`e��J��W$�;�����k0��!�o���<ޘ$H6J��h<�Zp|&��p�e,va�x
�wI�y/T�l.�4���|� �c!+�>�W�QVaȰ�.!�����J�Z��bs!=�5د�d �0k���+���4�Wr�Y���C�1o,7�J��U(�%�>C��)[_��G�dYk�̡�DteX��aT�$K�m�Rk�t�'�^�Rrͥ@��	�*/�t#� �Q�քγ�
�o۫#� ]=�TKx��h\�\���%w�A?Ψ͐�||$ݯ�E�S�kߗ+��tg2��j�l1����bHO����D�2�J8����yF��x�0���= �:�Yc�&�`�6it��
��5��w�s'��O耩���Y$K|��(n��*��y���CLi��
�-<YDu�a�W��K�t|�`�x�U�� QӮw�w���]b�D}�=����%���ce2�ϵWD��t�aBܾEJ��	�7����5��n��E�߲������#����8� b�R�&m��<����π�Խ�n���-�n����g|{��Nt�9���h4"�,����'�o#�H�v��鋯�pl��X�m�6^�����f��f#}��K��ř�g%�{�H���j��Qr��H'��p����Կ�~��$Ń'=rI��mU����Z5�ػ����&n��8�ª�
V��߬ Ӣ3���7zN�fS]�G�jWa"��SKʯ����"��0���� �(�����������e�C:��Krԕa*y\�N�b�NDA8��S�ʵ��n!v����.z�G��k��A[�a��cm/S�n�B�^	�.�mQVM�}��P3͚϶��ު
�a9������u�>*d
����|�U~I��F-5w���0}"+3Q���B�'�e�$0���0��Z����Q�MR�9��97D�<����*�LVz�G�Q	�t�kSR��3h�SX��p���ύ}�����{���4�If�=i2�n�c�ՏT�!����1(��b���!���)/�mqv�i���&=װ~2�t��z~.�d�c�/Ȏ�v�|b`r��;@��厥Gs�x��y����Z�o�K�:����3{l��
�pf�n��C�n�I�P��0�w�lc�I$�������S��<���J������<pQG��'�M'�=��_��\DU؊iN',��E@�	ˠp�k���<�6�k����ê��U��f2�콜E��m��U*���VÅZ�/SF�8��Č������}���s��w��D?������̈́�˶�'aq��N�~��ީ�S�S��~F��s&������69�7�o$����P����D!��κ�k�¨��p���o�`O�R��WO���ϬIݗ���Y޲C=D\;J�[	��w�R�Dؚ_ڧx��֢�m���]`�K���kA,WA��V�����p�^��#�6@�Fb���1~��l�X̙j��?���9���Mn�	}���s�c�=��4�W����֑#>�f��6����A��t*m�f�k�>A���T�0�2�Go��q�C��m��C�A0n���R�S����#���z}sH~�k�ߣ�])�i��w�+�6U�:aS���+���l��d=i�E���5	@���_����=�Լd1$b��q��`�*�#�u`$8�LL�):�%s��I+~/X�����7��}�~�";�in:���A�݄�WVc%��ǌ6�2�"��7J�� ��h�d߅�!+�r����5����FŴ��Rʋ���6f�f�a@_���,�B���h��(�1��+��I�i�1����
�x�%�������UВI�뢀���)�ʷ����?L
��u&�y��~$g��uNEo���^����
'(9L<�����~�J>F�]�b���ްk��g�z��o[\�F0�;���#" �=&��
Ԍ�Z���_�šĈ�臭���GYV���:/��,ޚ� x� ��ͦ���a`��K�[mР�����yZ����gi:ZʻW2r���r|�U�D�� e���>Ia4H �6$���q �n�^����f
��[}��uU�hb� �e
�Z�C��B�&=�� �\����?��9V��J�J�����p��U,y��b��xL�sK���V-u �Ĳ	̻�ݥ����j4_f!�G���myg���a�j�yO���^E���a�ԬN��.�Uq�-�����߄��<��p*��L���*&���(.�`\ol�e̥�A]뀇�U�w�\���7\�Jf1��1�w>|����z8���
� �V.}�X��j�-���`La�������M��f��j�^ ���!�f�y�<m�ҳ;�;5Ů��v����흊�Z'X"��9��QZ��	93�s�%���GZ庙�|ޘ;RTXV0��O�B:l�豹	�:�O�%�^h���C�*z�0�-`��G�bY�-y�d����h��
;Hb9�yOP�!�_n\���eg#��� Ψ�%�zwC�Aנ��,ݮۺ���"�:A�5�]��[5�E�p���3[3��@�����ȸ�ܴo5��7t��?��Ic�`���.u�U�NI�'`���چ��{ NJ�L�--�5��ߗ��������
��<}q	CyO�++�j��-���.@�3W'��[ӻ�(�>" X\�9>���g�ME�G�#���-�)ʼ��0��(y�2|}���	pI}k/R��qSC{H�B	p:H�%��h�~��X�uBu������ �%� �Z�E�Ú�>PD�`s�ަ01��Ñ�ә�<)�9sYQ-Dzk���j-�����5	q�[�ʞ�v�͢���L~�/����;�o�t�����рh�2\e"���ŵFsb���r
p%�a�<Tm,N�R��Y���2a@��aMڥ�<�
6��z䬦 ]�'� �3��ʂ�x�_�����d�=9�y���7ץ�;=oH�%�/e��5�NY�7
)o�~F��=5��^9�ŉf��E�-NМ�y�e<�e\��~ʲ�!R�Q��Y��aU *7��h������y���j�&f"����s��Z��������;�:����/�Ӓ� (\ZqO�/��c�J�b+�w�հ�Y�P��[����[��i�j���3�bٰ�e�wb<��&�Q#�t��+�2�,��	�)����+��p�����q� FXf�}; �3�p1(Q֌;�82�8�-�5IT��P����`�%'�gt��ZYrk�׬#��U�8��X+.�����ֻYС�mG����_�[�!��=� ��Gk�E�Fc��\U4����W��Dj���g�%�f�E� M� ���},�'>�0�^?^W�x��K��r��]*�O��LC,c�+C��n��3�}OX����$(~�˕�F�܉j7N#��'�?��P�E>�Ca�Q�Q{ne��|8=�{83=��T��r#�=(*	Wk}�Jv�!BҪG'\����I��~��Z D�z�u�^�6�I)좴�S�b��;�J��u�����N7}�/~�=%5�ay~����a�ADԾ��Ҕ�j9�5�+��(a���X�F���|Vظ��`�9S��{�v���⬬h#�B��9�6��������&RXx�i�X��\=�гA�c=/�]�}a��1�#,�S�����-cm�I�0�����:ކ�#Y�_��Y\V�a��!C��%7u&�
���U�B�Ҁô;��u��:���/x���j��V�!ov.��;'�I�1녜�z�����/�j�Υ������B�n�Mcd��y>�&?��2"DP�
�!�th��u�3߉�Ic�jt�>��S�=�(J���؎p�)�g�O�v�l�X��Ǐ�fB^:^���0h�v��% �d��&��q�dP�p�@T�t�n����vΝ�qz�
r��0#W�(, �h�(GA4� ��	��G]aĤ�2�t(��x0�	��ze���`L�r0kMّ����W8-	��Op��_ׅ�K�h�d�z�"㞬x���`/��*�[������*aφY�ćV���=���]����xxԞ�'2V�^�j\�b��6nY&�@�3���%���|,~��<�5�ٷ!���9�I*o7�>�(����Zc�NߘAmԼe���"�"���E]�50_���Pt	��;/B���X�(�^H���>`�EU��� ����O���OP�̈�J���|=��R�������z��BZ����X �>}Y�'X�!4�c�c�9���{�^����2���}�Q��hHq�Nkd����ѐZ�׎b���������u��Y�p��߄��ץ�w�X���ی�,�i��4�Fʨ�5��m�5O���<����Q���
��^�U��]��u�,�o��BD�E��z�|3��g�g����ʋZ�K`n�i��+5}G���;r�u�.�6����$��ɼʫԈ�����5� �J�H���`c^|�����YE��J� �1�<瑸YY��?`Gi�E�%inv3`i���HTC�X_��%ǈ{>�V�_�F0����n*��ݺj6	�7i����Y���\P����i
��Xy�F K�T/��ZM�)Fh�EA₴�HNFMR%6�.6��/��5�'A���u<Y/��Z�^�Sm��A_ʧ.!+І9���w6��@�>�3�Q#��n	@;�}����&x�����I�,��tk�Ї��蕼sD�w�e��gg9Xs��o�z�{�!�6�Z-�y��R)=����u��Y�����[��<����^�M/P��,P�u
� ���G֮�@K��A.N�.�FM})	d/A� 9���G�usB�w7�0a6���+�$C�
��I跻A��n(;�U�,���YH�&W���@��}Ƶ'�oe~~9�b�ʤh��L��۫l���dNTQ�:��v\��ѧ�ϱ��(������9e�g�a~]V���D���S�>�]NH%C�3�z��ׁ�d��E�o7��VsQ +�u+MD��bꢓ���>Z���e&�-[UӦJZu�<#B�O�juL(�k� 69��� �� e�M���R7HрV3�o%4�d�993Ә�z�Q� �%�ߕb�W�*��v���`P�	Gӭ�~JP�&�Moj�J��pmm�N�l����-z��ǏO�X��E�T�h�.@:�F��!���X:�iga�+ht��W��l�G�a//���� ��s����M^lX{]�(�Fd�3qvr��Q"�d���4��>U�\~mw4*���G��)�m�FsJp�3W�/wĵ��+J�sTwq�q���E�rh�E���K���~�#�Q��E����ֲ��x���,���?�+��l�eKU�8����	�Prlf��G߳��m�~c����:;�2�>]3qN�rΜ]��C1q��}�� ��x�
c��� I�S�E��G~�mN�`�^A��YD�1��{����0��ct��޿q{�Y!�W����Xx�sA��
��"�h6#j2� s��N>~��?�E���N�t�k+L$D�PQ�Z���=�AG�E	��ꮬV9`�?9�������������}"��-���nfL�P����Ԃ|L����<�j�OI���(�<�MZ�8$��N"��������wC��^r4� �Gfu� y�}3Ǔ@�}�)����Q��>�r�|;4ͺ�g>~^�{�*ՇE����}��\������%�u��?��Md��Y�ep��ks�
ѩ ~�hT��^G�s�ʸ��(�~��]t��DY4����T�Bd�U�3��M/��I�����snsԗB�`2�7��m��\ �\�ﺪ�� ��Q��`���B����	�M�y٨vs��,5��z^6�3����)�o�'Y�ޟ���'��q��B�̰I���D��@���'���$�6�]�m�����lh@a2`��U���/W��bqb�j�ޗ^<[�\�)�5���,`�m�9%�_8��MaX>���ƒ:�%0��WRN�Ժ60^��x���DC�#U�A��Տ��yy�ڬz>	K&v�"�M��4�r��n�B8il����n���Q�����,���(���(�ف~r�u뽑�b��~8l闁�oG�w6�^��m��lƌ	� 
�0��D^G��[;�,d��亮A�A >{&����6�
��u�9�{ ��SI����[U!���2�uC0���m��F��C*1�6���%���w��۸M�X���Eo㰢8��L�u�c#�@��0di�;f�_�Լ��-F��y}V��D��!�3�����@���j��+ �Ά��Qc�}�w��\��3s�w��t�.�nO7
T�Խ�'����i�O*s�nJ�H�2��Z��-�u�;~��b��<�L]z�9-�7v ������Qj�A�Ǫ�Ҭ��yjz~��R�*4>C��?B�&n$��rf�@�;ph�<�ꋞy�#P��������hvb�D,��x>n���FC�<��y��e��C����O�oS��
�r�LC?����$�e�?v�1�,Q�b�5�ɠ`�m<?�~�zv^�.�
m����֕�fƂ��a���Ws�0U�$��]Y�E9 .���&bzA���m�w�W#���7v2m����I�Ѱf:Y�����v�~��Ջ�F��0 2�Ѐ��`̱'��˚| ^�<��u��6�����|��@��Ј��`�遅.Z�,Q�n�7�}��*�PM��X�A�$<���^�<���f��*�6$�����X��2"�t�A��O.p ���c�E��f���@I'ȿB?�b�y�ӻAб�oʴҮTp�:��j�:��Ϥ�a�H���נ��͚��G�p����I�N
I���?�mQ7ģ�{��3~Ac�)l�ef����'kg5��DA8qE&��he�Rѐ[�)���|�Ѐ႖�orw�J��5�������㓝Qhy��ӎ)֮��`��!F�����L]EIE�'/�H8�1��a���E��T����8%jQ��Q)�����<�(��j��`����	���6Z��B
%}���s'pri]��Eu�:��#̸��/��J�	��l �忤�ݞ�ݕ��ƪY���R+��(&|�]�x�q�����,��H�b�*-�P�0e��b5C��(�)ȇ�BH�\�|�����T1j�q+/�x㈑�|m�"�v���3�nY�7{멁4|X ���*}������ns�6�P6b'U�g,��T�,�QIw+d�o�m�*�e?hX�Cax�|;�D ~JH\��]!\�ݪ����*[��;�v�ֱ���~g!�dv֑���S�U.i[�h�%BF���V�%�8��7�3I�|���m���=�C�7��TV����Y�N\��"8���=gq����<W��� � ^����L�Sa�J	 8x#��E��R�sr��ShD��_|�e� �a�� �)���/8��П�����ڜ�d��1W	��}���X֞�[���<L3���C�n�B2Gx;<r��SHmHc�.nj�
�nS%�QDDv�����ψ/݋�t�̇��@6�"���C���s� �bb�"�;w������oM��U���S~�Z���F���k'�=��b�����D2��s�C��g���!U@k@�Yy�~Q�l�S�q�/��MK�8"��X:�xIJ�9oM�ƗP��K�D�]�Y� +�X�A�՚��W9��48Xn_4(w�Xw��]0��� `��[�/�b��I��fjo߷U\�-/�#D1�ަ��ቁ�N�'-�^�o9����Pa�5��S�R\���0����_�m��6�X8�@&�h^�[� �X�{���G�C��zv�t���Xm��ׄS��m�z�u���9z�c���1��\�ёڞ�I8� �[n��J���59S���������J����DL��}s3�o��D���m�F>q��rdtˢ���g\�pP@�h���HLK�������ٝ>�(�`%����Z��b��+��F�C���o��X�2Uo��l|޳��[��J���Q-�&Bv���qZc�0�>ZQ氞��n��rK"
��8:{��#���C��ͫ��\�~�QP��/M�02J�|�C�Nwh���]4L�m���	����΅N��N!$�yt�"&Bd�~!Y"y��{P/�MRo��ב+�8_C��^�a)���SN$��&RSh��5P@iڋ����1�U�n��i�(�w�?�(>�.\�VA�ҁ|�hP�-�&��Ȃ{X��B�Z�y$ZC�ǳ��^AB��1
Pn�Q�&��?��$�/���94���\|Z�)��H��ׁ�}��Z�J0��	�F#�K�l���p�m{D�H�6�\�k	�� 5�V( )�=�K.�oK�>!�)�;�mA|@���j���Um�f�E�׸��'�HY�<�n� ^�Ϡ|	�5ֻڷϐ{y��S�i�}����xI���[xd��}w�bMNv_��ZƦe04���J�?�UY[��7<�:�Kd��]��ύX�o`ڳ3"��,]{gy�v�e��PA�E�U���~�G�_���k������F�*�	��s��1��0�G;�d������t	p3���-�2Xo���zl�~�/S����F�$G��'�p�!�thoU�	�Y?�wcZ��i�P$<9m�o�W=!6K�X��or��D[_Ŧ!c^6��|��N�1���Y��'��$ٌj몾�?ץ��Ԫ�@��֎u 	P�6�:�A�q�Iu��z�Y�����3dM��'�A�7D�z���b�T3v��-5y%�i]���[F�|W7~:2h�k��`�&Y��~��rb�6����t*:RJ[7sOnS5⎣Na�[zHQG���L�/�&��ؓ$h��q]���U���
�8CB��r���i\���\�H�:��gY�SIƠ�� *�^����xl��(T��T�����Қ#ED�%YM����zN9��K��V���������(f�?��	�	�Tw��z`#�D��@7/������҃<����g�x��\�wh��G�p/�b�
c�?@G�Ar�M�5����|X͆��R)髬�:�uX�jY���@�����6����o�z�<7�{���>�* .��"L5����T��j�F.��`8�;۶i.-��U[�m|q.r�`0\�����	�E蓞�6���u���.�dDŮI�m:!�1��QHֱZy�?|Ao�߹�ߍQ�����:���J]����k��v 9�`������m;��N���\.jI�F���|'{�&P��aFM��	�<��h�=gYL��zc�4�{�z~�''U�]xT��À��<U����-��oqy�3��?�Mߔ�@#X�Q�JYl��&��]A�3�/T�0[edW@-�ڇB2�+vHȿ�{�b��p���pfz	�t'>*��/ZNS0�F+��Q�uMF_�t�$t��D�Gx�����W����C������U��}���1�1��S�Uՙ�~p�?����a`R蝲�`�=�jL{Cԫ�q�0��o���2�%0u���	c����ꢥ�D�a��5}?�)�h)��=�25���ơ��C�܃*�Z��4ϥ���|��6�@�LH�	Ht�my�븕�R[K*�3+�I9R��|L4���_ t����o
\�r��2.�E��G�%ϝ�&u�($��K�G8��]��mr�e����v[./������q���-�bg7�㼩f��tZ�h�<�����W�q���Łl^҃���[�['D'J
����M�cGp|ƣ�s[��v�S�Z�Ub	t��r.��Y��t�{����E�����"�����,�Ng%�[d�kP�n��~qB��AU���ԫ>��'U�m&֟�
5'�4ߙ�u�?e�ϐ5�]����f"�e�8�a��q��`�*i覘w�� S/�C�����f[�gA�L�G&Eo��Ϋ�&����ϔRp3t�a��SYD�p��$�	�cP�l5��>f%�����1v���`P��d5�6�=���K�����Xs�?��;����Ǉ����1A���=�w��d�B���dO�	���i��
�܂���stx��d
σ Q�N��4�)��"�TM�_�G3]՛A�����W��q��Ǧ8�����K��YV�ܭ��b���d��N��ݻ��YB��e�+r��}�wuc��E��>����o*��� r��m~h�'���mAӤ^����`�!��9���H��9Y���ue�$��톗���^��Sb�٬o)]��رc
���1\���f�?��,ei�H�Y#�9�~*�}�>�}#Ej�=P� 7a� ����S'w�ޛ�DL]�;�V+�d���&�A�!������T��i�hOr��V$��*U��j�6"��Ɖ���o�TPi[J����
�cε�
cb%]�1�DA"�䅮,͞�V2+i�)r͕�G��^$z6(�4�I�� ���lㆿk���\_�'j	Tne{΁�[W�1H���}�!�Ҝ_z���|��ޥ }�˲��aj�%�٥���N �d.e57CJ<�1���ኋ���-n�����S�{��i&>#�L�U���|H�U�o�����ti&dzrWҵ�[��� 5����J+h���}���m��9��-�`ҿ���âO�=P{��}\<Oi �X6!����Ęn�J�(�-��g��[Aar�Z�]������<S��Ր��ThJ�Â��]�7����~������H[א�9Z|�	�Dr[�D�1�qv��П���̵����+�S��X5��2E�<��#�����C,[�Ge:Y|0[EM|��J�!st�v��RS�돸Ncs�Se��Q j+�e�la�P#���\؆�% �x�l.B�@h�[M5���]��h�I��)�e��Ƚ?��4��(s�| L���ȳ�.��\�L��)d#$��[�*:7_y ���V~c�e c�Չ\E��	��,R�<�ح��\���|��`M1o>g�7��2�$I��?)sJ-\�4�>1�b)B:8iL�5���֢�:�F+j:|J�\��2n�B����3 ��_Z�>!$\) 0� ����H�r�֏c�W��4�[����5���w@5���\��0��I:j%h�'t��h��;���WPMA��f��!���t��j6��[�ˇ5bm2���8��2��d�/��xO#�����`�O��j)�]�^a��='���l�;|��a[˖ʅ�Ǝ��#����Kbs��`�{Ѷ�~e��+�#�W.�p�Jio�5s��c��ղt�!���a2��tKN���t�;AL�mG��=�g���{�%o<,u����7��K/��
��:�c��m	�g�b]��5�����a�e]Y�B`L���re���ų�H�U�\N�[̑�bP%&P�٤�r�Q8H�m�l���ߢEe3�F�l��4GAq�F|��
]Ē1J��ƭ����yZ��_S��uK-�xU�$���1>�4���-���U����W�L���졨+����y?i�H�b�n��P�ŔZ&�����+[��o�;�3k���&�۸��>"nA��gĒ��m]։A���n�����������As��'����4���e��>ɇ���$��x�9��0z'dӹ�M(��eg�׽u��-ƪʭsYd��@��=��O��9��MS/4H����O�)T*Fz��39-R��_]K��,��Ue�i��Z W�T�pzy�A�����"*�:�����g\u��+��W �v�?�ݳˎ�� �t�P؆�`�M��춥�|��;lIP!f�mK[	��p=��)�����
���0>���"}N��՗�gs�t0���I�h�׀Ï�~�0B~[�޽������s=��2Џ�g ���A�7�
�~
�Ѡ�q��q�+�2p�w߲%8����:�H9����*oG�)Vx,:Y>+uΗ�g��K��>�wI��U�F����ˀ�͒BlG\�W"�M�TK���G���G) �l�'@�x������,�Qf���ʾ�����3���q�(x�ɝ�֮�f�y��D>!��%�]Ÿ�Z\L֮�{��d;7�Ș\A¸OЍ��2[4w��#Ld {B���S�Z
��-WٙӒ��FVF����қ����n��ɾk�w�?��{���6��STgrB<W?(�@:&^��uZ;&	q��^0�����|I�Q|�fm�G�H�M�������]�[�qX"{H\	�wMM���8���$l{�h�������Ɛ�7��s���vh�`�#��j5p�$���[�ei Ŭ����%&�GK�[�܉]�u��h���&�}(k� ^�w? *藏lToh���7�p�����n��ZMN�8Z�G^��Δ���7�`�wu}#z�����;^ϼ�d��ގ�ʚ�U��^j��	k5-�rE�Xz#���-�s�6�e`NRH%��eP�Lox��CJ4 }[��殽�/tֵ��)b�]����0�����t�_޵�-Ǖ�\��ST)]��z��WdY���3.}-m�=ՐkҖg�<q�eJ�[�޸����h�5)�IM/<2����s�0#=Hé�7���v[
M�.%q]�u�7�@7�c�Ֆ_Ei�'%�^�#F��D�A�T��tc}FƸ���~�����y�YR+�w�Z��X� :X�Y�a�/M�*��)sb������dc`����[h�!�O烈����H>�:��]�_|$�hR�[;�]M_���Rԧ�x�H�&�yOy:�0I����҂���55Tȓe��>a�(s%���Èȩ~���v�|��oz�l��䎥��B�ʓ�Տ���Tz�����;���?Ͽ�zF-�&Q	�8���6�;�T��z����V�3�0���w(Jk攻� k��n�O�].9N�`�z��D��0�)H��T�p'��4��%�%�?:}����!��%g��~��I������("�M�@��fA'���~8�2a��lgx�q��w}���ٳ2��A��da2�0f|��Ӆ�y��HEb%�{�iJ�ս�/u�ќ��@v^�71BØ���ԗ"�h�
4�*Jd�����|!.H�n�G[XemV����qvݾ��_E��9�>�;n�)A~5�*V>���h��S�̶>���1(J��N�)�b\aU&s�|I"f&�����2?���y�po�v���ݲ�d��uM,6N9�}ǆ`XB�0����T�F�Piǅ )m�2k��j�eoNDH�;?�**�<�����I���
�̚Hh�8b;�*�W	EА����@�K(���%:��s�h�-T�x,��۞73�-o��w��@#;��J1e�Wk��qE�8j�όJEib�uh��B���2Ф�)�W@��H���=�~�Dc�jJ#�`|[���d�M�qI*�,u�7Ÿ��Q����z��%I��l�y=Z2��`�αċ��^��/�[�1w���#��k�x�߇^oo���k ��������U�]���ܻ�b!��vM�����A�uͲQ؂׸Q�{�yHu��F; �~+X,�SV��������ǀ�U�`�ˡXTv[����}��}�#�ID�M��$�!�:`n�d�"�Ñ[/%\�������6����Y��,�{<;K���N�c)7��������&�dl�/�"���Ji�~�1����\��r�0A՚_�O�$�&4s�����Q �����U~Y�@����r�;w�;F,��Ɂ���?gH;�=u� �R�f"�.�;�o��&K�"}�8]z��]7u4�NK[$+���]��]&9�3�au>,?J6p�����o�ȴ
�������KB�(Zd=!�=`@w�D���9�L�#��+�Y�5�n�1�,��Li.�0��oI(��U�G4���5_��q�_�j�^�M���8b��� q5K͢���p����Ɍ�}<��(l�6�����}��Gծ��d[ ��#ܷ˃u���|��iH��`]kҩ�X����������j��D�g���eЌ�QZ�w��� ���]�����~{�/ A���SϵIF��Jn����	e�s,C��������Fw�Fg��$���}���eɔ�����27H'�T,Ԩ���Ђ��g�˓&����b�HS$uKOj݆�)��s��z�r��8*�������C��m1�U@�x������7R9k�H��O�����S	@��-��
P;&�,l^s՚!'Ӡ��4�,��U�Ip�����~	�E�����3b(�!fG�w��2��R�Y�}�L:�3]��^U{Hߖ Ț�v%<�~|��wg��Ii�_q�o�~[X��V>Fm>�`�f�(�cp�*.�����Q��FI\d�I��p��Wňb*Y(%e� ��,�}���W�)��d}��3���߬�~4nd!N��H���t�_�x�9�o��h��Q��>v}3���M��/Nw��;ǯ���6�0�j��uNjE+��ؑ���ڼ�6��&3��C#�d���`q���c�=���\���`e�w&���䄒�D�v�%^2�م��]�E0����z�-M2��H:������R��-M%X�����F�����1�E���>O;���+A�%�j J�N�)�U|PcR|^4)�����E�hG����X�B�J�������Ĉ8��{ï�AɝQ������i6��?5�7�Ѭ�s>���%7 n�o��M�(Oտ�Ӏx���|���zMFQ���E�]����F��>�H�1�yL�<��͆�.��U����7�S�j�����M�&��R�uDN̳�-Hռ��g���\�%z���� ��뢜1�(�1D��z��%�����X����B.M�o=l���ەu\��) /-��X\�(4�Ag L�y2*��p>��Y�y�j�g��.R��^P�h+-���zU���	z �D�dA<�(�}ͬ�A4����=�?����?N,9+���P����ф�����z��,��n�E��{��EIk`jO�Ώ��Ɠ69$�r�.k
�/�^�?��zF���]��0T�w<�"�^��l���������ٱ��xl��)����29}|,�:K1FS,F"T�����N�:DtC�y��:�ъY/��ն��j�mP�7R|j=T����D7<���,�JBPJw���r
?�L�����Lv�g�6�=��Z ����>��`:�g��x������څ�K�|wqs6kD�8F�%!�j��'��yhK�I��eȻ-���<�S/�����a?1s��2=dp�e���/t"M ���6o6]Q=s)e�M�1%J���/�������M��Xؐd$^װ�ه���[&9"{�]�m������M׹���RWBn���L�D�͜�������Xz>��5��ЌX��$0��h  ��,�}���J�5�s>@k�"��wZ�}{8~��U�ƿy_�R�o� ����`����u�%��v��N�`��I^���K�g0	�}�}�,�	�p摳�X���Xv�KF�i%,���dT�؉�F!6�0l�(�o)V���C��O&�����J��1�=�7gG��ᾊvF��9�a���%��ƒ 	#�2��ٮ�Pϊ.�G�K	��0����z~����s�'~��BҠhjv����.mJ�9KV�gO��x���'wx,����gS�nK	�C-��lt�{6��v:XC� ���k��)8�@�W�Sm%.PsVU�g�����'�o�2bt|y!���S<�|�b��H�sV`�����̼�ӕ0��U��>K��C�D0��/�s��ۍEU�g��3r�ͨG/Ґ�lJ���h��,��c�f����8�>G{��.����^H�.�&%?"·ذ[pL˓U�C�g2@�ٯ$)���M���t�R=}��y���Uy�ƵߠqN����Ì�;��Lm��x�}��~{���"K[j%�ş�%�p�����vdh���7��"Vֵ����ӓ`��� ˁ+N��kN�X��t)�ӗGR�G�����f ��ܔCy��2���]����͆�j��U�Mh*���R�+�N-Rv?P�kG~�5�|�$�|Xm��Aa:\��=���s����$M�Y�C�I.�v�'������bv%��Ѫ��������7�n-��qCU�p�h��΁ӛ�
F��5�|+iJ!&6T�6q��E�@�p_��5vᩢJB�� F>��-Pm>1ވLO�Í�׃���2��'��9;�ߟ_��@�ҥ���tE(C�L�q�-�E�=0�[����zh6E\Ws/�T�eɧ���ʈ��Z�q0g�:7�x�
���@cb
��Y��������E�ѐ�Nkl��o ��چ�R�_R�^7@B���WB�<������5vGau%�L ,������`C�%QP� F���	�1��u]<5��N�c������S	f��ȘJ�J�e��+ߪ���;Pks��
��f��/�TO�:X�J|(3Psp��W�tà%IW�IC��DY�jRȫ�B��m��^�$?�W���u4p	Of��W���Y���0=�u�]4��fQ�"nd�6�A�5�a��%��U��.�:C�A����V�ɾ9���8��2�N��;�`���Ѭ�죇~��ūW�c'�:�\b�&@���2���O��)�5-Vj͙��[yտ���P�(4�Y-)�{���4���L�W7L� .��!0k�������k\�dߓS�lpo��N�zə��j�����-��7�BT�u�e;��!����(�o��ȅ������M���">��p�AB��  �`��%��^SSt�����ڶ� ���i���59]}�} �b
w�s{N�i0c����Ț���[!��Ej���+;n������G��7_t��	~/o%�i�J�7z�y�0�+����q�߯xBu�o��81�Y��l.o�1ڸVW�ݨ������M���C�|���c6�:�6� lsꦽ��댴mk�֒��k�o,�X4�o��kKEb�R�9� 3�E�d3u�fS#V�q�=
	X��R�Vy�ֹR�4��˃�+z,.S��s ��r/�K�6��x#B	�U�EK���8��	��BM2��(&f	&���Ǐ����(�EQ1ޤ�
w�m(V��A�`��ʁ_�em�5�&�uf.Ы��H��R�
&G����^�b8����Lt�h���[;�%�`��rM�I<���;(���'l�݋���3�Ľ:��_ �&j��Ȅ�73����g�#�|(��f2c�������mA�*_�9&蟔!ddI^��<$t��f���m�/O�R
�zG���~��D]�@�ضt�B�k�]�Jc���N�w��;p��{�@��w��sbVSB��~)���ߵ-�Ɩm��Jb�W�?��Y�oIB�)D���qG�B	�������P-0�cl���DE��)�#� �Rq��C+�-�Ha�0�D�c;�jʣB�h�0ɽ�Xi��=Ч5�i����;"ht�dM�"�T������ev-�c�@��LBF$��D���b�[ӽ����[�I�O�H�b#t�e�d�Y�����.�H�!���`�1F�q�O�˱i�@�w�}�da w��i3���A��|H�u�$}���j�G���f7Z����`���Ӻ�zD���t_�3ikξ�'��w��[�{�Bk���'���ͪHt��%�(�Ѥ{�s&ï�6[1'`�j�VO�A�vV�f�yd@�v��ޞ
2F����'g����*�o� �γ�r�Y�0SI����������4��h�z1�Ǎ���bSy�%RZ<��nQ�_Y����{�Ѽ6�h��%�/�Y�i#���#�{�c�/A�w��:,*2Z$��8	S��<�U�0�����y��N�����0��?�T`��s���������Wp4Qj^�}yxe���6��$�vR�8��3��1���x� ��=�}9a*M��6�O�+�M�
���z���=�%U�M.��C�w���֗"����"v�ʾ
�0e �[>�i�4�<<�[1�g���"!�x�z�K�V��%����ڴE�c��������_��9;�QS�!A�=�辻�BK�xu�~I��`{�i���:�"_j�ci.tݩ~Nakb�.T7�X�7�[|���C�B6M����U�x��i�(+RS-�-A��W�g�m�/�{/b�x��2{c����z�ԍ�ݹU�~(��̊K��38;��L��a)w(�j�g�3��h���ڞ2�AX�xHH�~�@�(��5���q�ګH����+���|	Vxw}��M{bu�i��0h��gY�̆ѱ<�H�!*?�CR�bn<��K���a��Ű��GN���升H�'۱�(E�М6�%S�K�3�`:�i�QB\�q��yxD[�r5��1��]�	~�"��l�aC��cxT�J_�CbK��V�U�Ԇƣ� 5m��3I��=��f��$޺i�~�)3�#?jԭ�� pB�mp�b��T\n��-�&]�2����a��`d&+���\�����	��#y'V��,�T�l|^�?�k����S9/L#Ü�)������AVc��n7��8`�0�6ƪ�rM�jQ�N�nQ�lġ1���b#dxh�Ŵm���'%�C-kE�W�T�o�v�BL��ɮC~�x��f�|�ϋs��L�ۢNE+|gRR(�����X{?#������m��|����O(������j6�Ah`R��Y|�q�EWh�����|�;�U�3��_��ě5���Y�U��z �I$V�Kݪ�$�#|�Yd3�aW��b��hwcB����N}: �z��:��� ����>Z���Ui)�M� yl�[/����_A���h�l�/����6z��W�4��6���A͗&}��sS���JKc�&���oz�pk���c�P�Z�� ����dKK�|M�=�
v6 s�׋>�_w�,�o-8��Y( ��&������{� �)5T2,|<l'=�����xT���������Э��j)��y\��/������Zϴ�N@��5	��h�h��Z�X�N?>v�![�߷g�R�r���G��L��J;Q�C����(�
�9w��nJ�U4��];��6M�������i&4W"���o�˞C��B&v?��;�j~���m�X M���c��H��2i
�|m�d�k��B�uf@:Kd6oe�{��"�4�u��+�A@;Kj�(�������^��	��[��u��O�J���,��x@ ÍO�P-�*���9K)ϣ���/�H�����P��I{���swg�Qbj,�6�bF�IX=nZ.���_Llz�K�l�+j/YZ�a�>4 L����L�N�>�"hE+u���%B(0�+��ҵ��*��'v�\F��rH(��5�D{b*�L�D�3��~R�X�V�sy��E�z�{L}�H��� =g�J�XC�)ɳ����f!�tz��? eFaD�ǅ>���}�<E	��9��W��!��굽�q����&QV�}ա��1�E8l]W&3�^�(N+���r���m
r�	�<�p�b%*�a��o���a�r;�gCjץ�ke����~�%7SsH��O=P�:I�;�~
k	\IR�̵q'˲B�}�T�5��N�H�\|5�i�ȿD���n/�e���~^�������������b�zF�I��H��[g��g�94�ռ� $��ݼ�6z5��c@����Y��Xԉf�N�������}D��N]�īԙ:L>19@aCx�;U�EU�I+a���aknz�'6�yکʘ�u����:�|��2�K�B��/0~�R�?��|N�M����g@��5��y�ȳ{��j>.�ï���dq+�kS������"ݍ%^uZ49j�vS� cΨ����~9Jm�̹����H\��\n��	m�س�{�=�:��NT���/TB�-9B�(�D.��v��= ��sF%��5������l�<?�l�FZYX�C3{�#���e������S8��gE�.���FE�8k? f��L�%��� �qq?x��A�K��'(ЇYX[�4�`����������]{���qX˷�ǌ|Ӓc)��d�m�������߰����Ƽ/~Aq��i�ܨ��|�p�e��(�z2���P}�Z��G���Lv�V���;z��Z$'=�R-���� J߻�S�E@���� ����g��~�Hw+����5A�j��E J8��ꌖl��sRrB�4j��_^e�� �m^����p�T[*x5����o<���,4�����_��}�Q��'8���G�a!���E]�����IR2�8t�]�Ӧe}������ZaE�{h
�	QJ^.��P���R��6,l<}LքzJG$ɇ��b :��c�<��S�83�h@�|[&pvT:@,�{�
�Cέލ��{E��iW�OZh���l�;�F�L�Wɏ$A}=9R�Џ<!F�-��ѱ�:ӄ�3v��r��T��#�17���>a�:\�?B�Z�`��Z�`%L�D ���^1D��bY�-��a��EK�>�~ָ�I���������ٴ�cDLQ����;�]4A��-v��vY�fB*�\0�S3�!e�%2'+3%	x�O���p���>���-Px��l��L4�%�J!\P����ǘ©D;���Z6P�] ;)��s�̐5���P�u��r�f6<e-M%/��~�K���-�p�Ⱥ>y����q�Od���`r-2�C/p���鮓�T�%η)B��|r5��M�gъ�g	}?0�ǟ=Ԁ/����S��a�3]'��\޼��9��>��R���As/�T��*E�Y[S��-�y?�G�C?�	�D%� =��*�Wi9��m�s�C�p	f\�%�M|B��ɡ��,Z�T�F5�]�\z>J�(���-Z�?$�
WZo�ܬP�4�t���sL�����&�jP l��
�7^[��x�q��j P�/_�oX�|�S9���[q,��{���gNH���6`�w�����2�!r������0Q�,�d�4�������LQkk=�¹�DY]w��tقD���hbg��r�ep����:%����F=B����:���k7TO�}�c�1 ��b�i3�#y��`j*��0N�{�m�����:��l�%!������<���f��W٘���W��F#7=Xs$�7b;F5��c&zO�/�0�ZU=LX�O��L8�����\�����CŜ!5�� I��C0W� ����Թ����jН��';��-/�^�Cɦ^�
�+�ܜd��!��vC �����+�,�ɴS��K2@���ζ���� t����k5T��"�{?���)]M���X���Ċ��cL%�pi�5NA�I���YIZ�Bf\%�k����t���q��kn7[�QѪ�x:#��h�yZX4a>��rJ���$�9�4D�ǲ��!H���E�
Q�D�'����O��*�@ƙm9��F��Ϩ��m3�� �M#D�ٴ�馯� �]n֥r���a7����K�ׯ��G^14Q��xÀv
`�j)��Nď[�n�K`1n�މK'���QOˠ�=����ಱ~�0eL[��y ���x�ܡ��)M�6<Q�8�Q$�o9�$�����C�m�d�m:�-H1�4����'�b��v�Qp��7o?o*5���A}羍��	����q~�m�v*����HĶc:N��?�D]~�����D��t��~�=�U�z8�u5>���
m�es�LI!cb�nv�9v��6a@K���`f_G�k�F�u���ܴ(q�XĀ�Ȏ�@1�%5�+N.0�Ri�N|)ܥ�S���59g;�5�1(GN;�(�e�|������]���c.��S�s9	PR����K��ہ;���jq�զ�� }t0�d���-�&�|��H��&i�*n�H��J�y>'=��(��X\�}�`]�Q H.b�2r�����s{�k�t�;�����W0m@�w� T^��$L��`�� ��n"��Ѭ-�߹T�_�����K*�`��/O�4툎qV1�^�X�]�V@z��{᪥�`���3w��,�:��IQl���$A�wǽ��v�N��&������vKp�8���6��HA����� ����r�g>��� ��I�П��4��T�O$m�?żRT��~�}�z��W$v�0�r���ői{�{��'A��&�Q -���ow*�x���]��2�
�߸�� ��`�>�#gŇW��u��VJ��݊�En��3!`��${�A���LI�n��� ����ݒ�B-���hņk0uL���q�����}���"Cl�8
��ǀO��O��3���wU�a 8�Db��N�����.���~�svံ(4�EН�8x�s��*�)�3��P��Dm�V��L�!K��?�m=&�6@[?������&��Cѭz
|*j�h$ۡa��oV����Մυ�m�Y�8���o���6#W���@����F'sƇ��W?�I�Ϋrާ�6��6�j�4J_A��*�v��Y��s*lm����T�(��`�l��)���'>n!�|;4::��J�����~g�0O��!��%Z�/���}l����K`�����P�}��"�[�5�n�,�q��-��ө,�Ȕ���	��q
EJ�^�B+'�a~���
�h�&��`���}���3���`�D6s$a�b�t��հ����dc�/�j�Bi&�]�
r�qL�d��P��c^X���F�����MDq+��P�bQ�nE"�(L67w�Z��jC=/]W�ui(d��JK�tǳ|�<�eNx���ڤ*�7���i��Xy������$��D�\�J/�/�&�moO����@eh�1�*���i�ʦr��`�:nT	����oŬ��G�U���&AE�\-Ĝ�p7(�C��|/��񖺁hC�TC��׺ ��G��0�g���[���B��݉J^�W������
�z_����Q�\:�_�����Ra�i��I�<;Ę��C�S��2nsG�d)�D�t��6�^y4+���vp��ұD�s���E�/?��I�����\�Bj��%Z�5�J�-.��Wl\���.���йl"ĥ�2S^BJ�O]H�J?	?�s�����tp��RZ'�g�[5Ƴ�F�铠�o=`��ɔ\^MC���D���h��&h�Q��Fؑ�������-��K�,�Vұ��� +���E�����N���:�^p�NB$�/��Ֆ+�@����������������[� A=��¬�A�J���W2(��ҏ$��kGu�zӚ;�5�����3b�ൢV0WfE�i6�f%�D�$�������S|{�X��v)��tG��@/�ݔJNc.�z��l#8�B����xiU�TdH��5PJ�Cnd-|LjL�>n����<��a*Nq���vu�Z���@gt�c���K!`O7��ܠ�����q����x��p�=��(yj�eǒ�^#1p�
RsG�f=OҚ�����juAD!�@��-�f(�8D�|���֟�j���������V�0^��L�+��&Q���:U1{vd���g����R��oFѵ%�����z�_�~�.v��hF`�Yg�h7@xV�4���8����5�������Ab�҄�ܯN���%�;b���XB�J�x =�SI��r$�J����̘8D�t���Z̢��a��(|G])b[Q{G�5?!wVΌ��
pkgT[��L�!g�٢M�f����Q�Űv�Ɔ��	|�p����;��0-�6}��jL�Xޡ���,�l�;nZ;��A"LQ���s�_�.ą�2) ��~{^L���gyU�i�Z�v���6ҙ���_%���O1��6ك�;�v"U����ٶ��^>��y̟2l%�5lڭb}H����"��C��<L���(�c���j<�YnhyVRC��D�g�����B��{�����l�2S3>`�{���o`���	3���@!�֏wj��8�� ,�p���� }��{�\j�)����ۍ	* �EN�|�[�,JeP��9�-�J}��Ɨ$�˥f����@`�(������B���7�h���/ެ$�u�FtS�]T�����;c~�u<�%� R�I���Rr������:��A k|��6EP�ej�((�P̺��ψ��%�Zx��Ǐe�ɸ\.� �4�5�3O�r�R�����	�~LA�n#�pe�q��F��#�HBN���N޳WJ�����kW��L�U���}�����%�q�Y"�(����c����-:��ap5�:��K� q���Bц�*T�Yw{��?�ټ�� %0*�k8E����Q*z����i�s�P�-�g�z��.HgiR=�������1��+0�֋�{�����\�yi�Q���4�lw٭À��D���!�$�َ�-7������]�
 ��SYH4P�	�]S���^��y���PXW@�B�TN��iinO��5|P���v3���iD��C޵É:�Uˉ����0�n��E!�
��'Z�{�����D4TJI�� \�_��Y�lw�{p`2{��v�~��ݿ��|#�ٳp�*�/�/'wߓ([��^eV�s^��a�cL׏�l(-W����;x�\�AC&�0���e 7�O%����x��X��0��.����\�b�_�*{
#�%=�_Q�e3sϻ����X����=��s	%o�G��o��1�-�n��~EqPх��~��{��F�S4ӌs�#=�#^��I68K�/:�Ԑ&��v��hMc�]��|�����E�Q�j�:�Fw�|�Q
J��s�b*r�m�Y��?`����^������2|��Y�S��rb�V�'��Aʼd덴c�dǶ:��pR��!h��Q\`uYGcϴbQ�!"2�<���D']�X��bɥ$'�e�7��GA�3C)w��N9�_���i�}D��%��i�2~K.0�2\���WJ��� ���x��p��tƮ���C�-����=�>(�2l1J��L��n���|G�	uL����.\�%m�� J�����>Xþ�w��[bS��k�X��A�u$Sq5��+���}U��\f��]z�!�踛S���6���A�V�`(��	B2L��9�w��z+�IXM�U�N���\�%i\1�..���IL92V(	��㡆3���2G������9����>P(s�6>5�΂BV"IN�%��z�|�"����%�@镎3��F�?�K��m���+��¯�̮>:�	&�q�v��ή9k�9�Ů��?�".E���_R�@ߩ�d��{K��>�hbK�{~e��S��Ge���&@��F����� t��J��c�{-�ʥ��c�Mb��<XU�|����_#����|�aߖws��LCօ7.�
�o��|;FQ�oV�����&���`'2xS���mB��E�J�]���*"�Յv/��	����H���W9�.;�N���l�Գ��a��H���ps9ʰ�M��"�B~��:�Q I<T�����S4<eP=,X���&������f>�F�&I��zf��'M81޻_�����-Q�9���0��Ӡ��^F�h',?�+��#��Q��Uy��av�<H����כ�C�x!Rv�[W/U��E�ٙ"�pyԩ��g�, �����&X탘�-��j�Lʿ��W��Ѫ�K���gM2|�����Id����<�K%İȻ,!�Fr���&����J��:�
� ��vh�J ���Ft2&���BZCY
�MM���҆/g�H��ǋo�wz+��gX:!��`/�p�6u?��^gB�,%V �Z <7^k�D���C��YdU"wc����v�3{����E��B's��V&��.P�0s�Q�t&�(�{K���\[�㌄F����Q�tRaㅙ�Vy��ᥘ��	t�$:�&7dU��%�;iэ�}�k��\����x�'<���y��:43q�NUb!7�1n�v���#u�\�H���Wß��:'Ȑch �c��C�Ț�u��iE$)~6��)�i���a�G�UF6��,
֦/�Ł�V�?mޜk�ڱ�Yp�(��H�I�XO��+]=4�b��8ͧ�azW�~5�e�$�s=�(U�;qy�m{%OK�[K��3��<c�6��)�+�(�/aϑ�/�3#��j3q����9��pp��7k�A|W��s9e��B͈����7PAcb_G�\]en�q� �>�Q�o�
���M���;0+�7=�۟v�j��	�ϛG�x����E�X@��ڸ���W�,��*���Ubߒ����TT(�p��<���t$v�� ����-�쉲[�d'Tչ�롓Lj�oiz����C����ʖK����xP��uN�.)��/�Xӱ�g�䴝R����&^+ N�VV�@G�����v�����䠳���,�+�?����69�n�r
�vCqþuQ���]	�4�`}���o }���]�k�5���h���Sj��XSY�ՅÀxJ�j̨%��{��޽����kKҒu��q��,h�iˮ�y>Bg�-��4#��d�]�ܮ.xG;G�������(vDB[�k]Z�)�&a�����J�&�P0E��ri/�{m���ۓ�d��0� +�FROa[UYT�����J[73��r�?zU�~�Rgry|����J��	�,XҁS^�zF=h?$hL�8w�y/�`�
П%��opk��@��Ia��\�_���.�%B���T)�SԎ����T��=I�'��s+�4/������A	����4��<@Kt�S�G�q�b��ٹ{"F�~R]�´t�%e�ڵtr�[3�����u
����jd�;���Q�m�����ee��LT������҄�1i��������=�0���xh�E XƵd��^��H���O7���Z��O9S�KB��ÁkE-j?���-2�;��g��-`�0��&=�rd=2�V�l+�1m���� 5$��>�K�u!,%���|4!k�0�uX瑦�����@./lkV\�\�.��,r	��b�uhgVwy󌬣d�$�Ts©iʞ�~�N"|��U�� B�P<K��ZԇJo��Z��� ����j����{pKV�qI>]���N!��)�,����9��i�L���M}� �����4��Gh�� �'���A[-@E0b$�(�k�v��1�d�#��ޛ�.
k�B����$�Q��#��?j:F�Nvz8� aT�@�L̲��8�~�T�Y`��!<a�}ɶ1A6�X��2�?������{c�*@E�U$?����`u����N�G�i8��Rjk),�*I��i�V�:q��*4#�H�G��Z��A�)>.}��}X5�|�O��Tg�c������5�]��l-xtc�y�"�?{�pƤ��y�����0� ���|�g*S�X����jM���ْ�,%����$�c�|2u���:�u2}b��Ϯ��u���	�B�.)$�=	=NH�?�b��G1�n��+�ّ���}ѷ#��S�y�2m��}��?�%J���e��"y�ח���xi��|��Wm�����P�,g*���q�>�rB �}=Y���;�T%��VtKpkɾx�~1�a��ۼ�4:�G>�_���(�bZ.aK %U��[�!���sMRV1���u�u����eU/�f��E��)��i9 ����#�u!��W�y��[�����A6�i�K�@ ��~��g���$~SP����/��'�<|��U��j��Y�ve{�:桢<�:���(ڌ{'c4�F
�ꗾ�dIZ��ᜬ�?p��r87�%wM�C���4l@��0C�`e������e��xB��	��uB0�YQXѸqDaJ�v�ͪ�Y)����{H��eT5t�Ï ���gh���3����Od�`+d$��8�[F:�C�M�-m�E���Ou)�2�V5iE�,ݭt*�%�����x��y�J�|$*���4Y!d<[ƶ�d�>�k���#3��Hu���+[�ص�<ݑ-W\ϗ �7��%A�r��ǅѪ�)T��=��. n���B�H��9��x�4�gR�[���]$�y�d?�(ow��Ǯ�oT��t���`%WZc�y��G�qr��<	�:p�;BoJV�(;�]��A��!�'"<� x�G&���L����)�As6�k�?;��M�
��Y�Z�l�����Fs����sfG�1.%�!Ua(w���P!D����[1);�gS�8���ɢ.Wd��BO9z��r����ʦ�lxn��5��q�;PP����A����R��T�,���Uݗ��Y�V��M:𸉳���KC�/<PO�XLs�J&����?��f �r(ZxwV/�^	����M\R����pC����/�'s�p�U*��z�D�
Wh�,cE��l|9��S����33ϧ�٤���bgĠܾ���0AW�ʠ�6
dA��%fL�������Є��Ky��b�sv�ޚ�ۀw��o��)6�ǐ��A��a܌T�J����4���"p۵����)Մ+4����7!ʭ����ϟ��љ}QY�t�4^���-��=��ݾ`=-z�p(�o�hѽVh4�^�@8:�{�C�vXh�d�����I��PEN]K{��۾��y��ހ��D�4�j젔�a�x&�^�3�Nl��h�q�j���p���@ܷ]0D1��J��`�o��������آO �$H�{J0���g����sz?�D��}��nev�)��!W��`%s� I���ךt�6oy���� �*���El�j��b��!�txx9�)w��*C~���ۃ��U0xn9J7	֔^B��$�g�)��s���,Z
��_�}!�h����֢9.?u�\��L�hq{��$��}�Y��N[,����3���V_�-�+���Xӵ.l?�F����=n��2g&����W8���Gr��|Ҷ�F.���R�����E���otF��5����ٟ�1:L�,)M�"�{���r��؟!�c�S����2^�J�Q�Q�#����v��^̈�)���gf@����rˤ-c�YL���h~D�:e�Ta6#�ޡ�<��!.܍1�;;�� ����!5��<�1y	������o�h��bMq} y[�>�Ȥ=��V�E�{!�J�(�0^́d-�	c����/7<i�j�G+>��<3x���cK5M�Kύk\7��@V���ZL��Bs+�����晓�]�j�h��N!��ѻp��h帊MI�KÑ�	�_��~��
��O���0o�̔j�&Kn�#su�~�[{��7��*���U�~ Z�R\�Y����:@n�q�"���~�I�E����k�m��v��G4�(� Y���7T9-�ɛv�LB��Gd>ev_r@h>R��cp��e�1������O�B�ۊz4��������z���H���nS�7 !����� u�� ��z)�|�Y���㌄��HQ�x���
߀%MD��g`0��p��3t�%"��9bn�p��1:�Z;wE�6�a�_ɷȦ��H���8)���f���U����*>IXC��L�t6�RDׅ���%u/�|�ƕ�k��b�����T'�]�E�B�dp]�C\�@��T��)��\{=����Hyz�N��;VJ����H ;`�Н����O�a����!��@NXr&a�?�\����Z�:�}��瀑�|��.e+��]a�4�7K_��I� ԗ�cci�/�Ϗ�u�l�����3�k9���F�b�>����T!^H�����>Vl��K�K0 �H�]��9;� a'���g.���F�:;�F��,��8f�K*��!�ў�ҏ�3,�!�*��sQ_Q2��o���R-%�[N���<�-�~��ji�Я*Pz��>�r�cT�,��dh�Զ�g����� ��W)��g���*�(Z��R�aA�u��Pg�����bm�������/ ��ʯ"��s��1l�!=lG�09A�¯�z���=G�W�H���^�b��z��uacS5���g��V*�h����U���^��s��*f��,���Y�}�x�I!���@hK/[ø�m�r}���0��'�e��z��k>G�i��Zsj� ��uȆ���ג�O��%�+|ӻ{�-.��'��~R"�&��ٌ�3"���j>J�PO ��>p���U���`R�s'��Ź��\R����a�_g	�k|~ۀ�l����"/��NoƢ���n�#�U$x�u�^��|��R�L,9�)�_ۦ|�i'1yj4�S��w�(�2��������b`Q����k�D����3�Pb����T]��'�(;�T�'oS)�a��!�ym/M��!Y����v�w�7�勔(�͹�L��7�H��@=�_���h��^�EW�:�Wڃ�W6`�vx��3���[��[��]6��7�!���w#�2s�ҟs8Y�E�!��x�<�V�6E�rl���5��a�@l�>���!A�����:�{fN�v����M���h/�^AP��|�e�.l��e�p�#(����a������c��ۍ�b�8���?�]�\�G�Q�q[veI�n6� #��+CŊ�nD�N6e�BOo��*%W:�H\I&{�.��������D%c������# ���6�T�^$��D�-I$vV�c;Qq�,Aߤ�U(���S����l?�iDm��hS�o��N��2�����]eЬ`b1�D�:�Ǵz�	�@�uC����,�31��[�S)
�wz���D��pl\	�&��@�K� ʩ�N{.P��m��B�Mʋ�W4�%��%��@�{� Q�aEu:K �&̍����8Yά~n�`\O�d����&c����3VXk�R�(d��L���w�`�A_��mNX�[���-�v�ñd�.�o�)<��V,%��J��O�O��!��
B���y�"�Dk���������'t��\Z�,�V�����m�Z�z��P[c'�q�	��~��;�gx(mƆ����1<��H�^K�/螘n�ĭ��Ü��DS���Jr>sX��m�x�E�H�����e�C�;KF^y%��N!PS,k��Ӱw���M����W��+ٚ�����U��_��g-m�_��,M}�	0��+�kI�U6�p���ɫ!����^29��io-��N�W����������.�
5١{m�vXMR�T�����6�8o��W�zq����\2)���l 2�<}���^o}J��w��(ert1F�i����tb��)�h����U��l�{Y�� ~=Oܒ������ � fW�t�Sl�2X��"�ˬ��_�(QP��=�AX���,�^A��2��K�H��*��r@�䝢�
}��sQI}W0��PA�g�dH��R.����o�=���ek4��s��X��R�C�����J�t�nj"�c0����>��c��b����
{�`庰��łܺ����^�I��I,Q�J ���n/�QK�4ٛ�m�2e?؉��>�n�d�rA7�Q]R����"���J۪2s����ie엞�>��w�3H�>�e`�?G�%
�al��; ��S���:��zi�D��qb�[�m�ؗ��ʘ>zܨ���b�zn!f�ʨM�X0�/��b���%�Ũ�g�g� ̈	��{��س$�~��[Z�~,��j�?��	�d�G��h����?�N��]p:tA1�AW�VGNfQ{���/�g�!�@��J�VN�P�v�\�kl����C3T��"�7��4��Q���� }�>�A%�W��>����o���D�G��tҎ��{�hL�2�nNv��h�!����p[���(v*���/24r�Iq�۸�ڵ9n�3�0�d�Ǻw�8�z���ֳ��>��f'%���* �����g��� �ï�rp��3k��ٔ��b�ŵ�*'P��:S�G�&k�R�9�-�4�Mu���9c88�?G/U;e,�_��DKR�5f���e�� 0�G޸�jy��eh�x�p1ztl�5�8~��A19t�����)-zJ�L�}}䥒s�@���o�u�zI4�����N��]O˯!/u���J~+ލ���L��q=Ή�v>9?��w�A����S�Ddߤȵ[�6����y�<V��uF�^
P&,"�.)��q`,�_�MĖ�+���Q��Մ���o�����[��l��G&�+�H���Ns��/`���m����ZҖ��83��r�3f���cq�.�>�L�O�O�G�S�N|n������=]2!P9�p+�`��ҁ5�<W!���K:�������ޢ&��տ�MO��;{Sopƴm��[{�=�*��Nxђ�O����!Y|�4w<DaT0�(��r��㇖So�M��T�]�>F��z�>��ԗ�����v�pgap���`t*��Y�xk���Xq���*�'H\z�A��$U)Y�j�5	�n�8�.FO C��{# ����;P�|m������9�Qީ
~is�=G*�� �K�FF�' X�9��l�7.��H��!�?<o��]�a2�rR���k��[�$��՚k����	��l���͕���5*1����t���?���2L�DP�2�u�oS��h���}7���@�����Zg�h�Wfo��d��5�׬�&Ž�4����P��r�@r���0�Q.�&�c��#6d��jⴓ/\*0��x}�S�NB{�I��j4�a�Ğ&�[�Ҫ!�m��q�Q�:C;�U�Q߰�z��;�
�)1u���SIrB.��^��+`�W�� ��L��Zů;D{�h��3���)ZWYS�:Н�wp��B-]�5y_�{d2��#��l��e��yM�mv���ܾl΅���[����G:5�� ����4�e�ِ��ctU�'B��w�r����h��(op¶�:}:���`[�Z�O}�_r�Ⱥ��ڑ�N���:�R��eg� �N��'�(6M�DXI@��p�H>q6�I��(R���b�Z' �j~�I9˹"�B���6�8�4��c9� J�-A���OO���^���?���8�k1/����E�)�ڊ߭Hx�u�%�R��
u��{; )&>D�V�z��S����a2	�cSA�󡏶vs�8�a�WtP�\6��0ڪ�_� [� ψ����$
�A��#)��e
0'E2�ws �Ү!a D�O	����{\�ʲ	�k�T�5�����y�/���� ��1g9N��ݤ��8m���ݤ�eC�f����efY-{�@{I����~X����������^��+�Z�u�n�k�X᣼D�����Ŝ'�(6����~M`
����KȡSQx@���V,�K��\RD�}�&�'j��Ϋ@�)�&�n"�ն�^x��N�ľm��KL�_d��٨eҹ�$�2U?3o���O���y��k~�>}����1�}!�����q!����OT���ј��0F�׍Oǆ�%傅�c�Ķ����y?Y��l�A���/���u�+�F1�c� o�X�\"���UF�S>����;����D�RϿxx� ����1*���[.���C|跁�쉚��V�*pv��=,0�0f�(Ô�$��QX�'ЯC�h��e"�{�b?�ya��e��@R\�iy�h�Et ���&�5�([og�;���#9`�90T�����z]6�WY��(�50���-6W�oG��szRm�\��y���}}��l );���z�M���L0)ÔQsFbls�ȭ�v���:�"j��͟��@�ɻ�FM M�*{��#@��+`��f�0�9��}7�E�f��@R� 7����M&��p�)�e�<�?4]";��~A��+-���Nݣ�Lt%+�wQ�I����E�0G������ך����^�p.1c�3�*M��86R��L(���C͐�w�1�+��I4��-3Yt�|]�З�ZT�lI���/�ț�b���Pf��V�=�Y��+�f�e���)��Y��-g�=��]�>q-X�Z�U�/��[�wi��yI��8�B�4��p(�{���$�B����o4�~��69�Q@���?��N�rBc�c� #k�)��<�&/I;S㘏$��΀��nX���<HG�d֦�Vw��5��`����HX�Nu�3`k����f�8�pZ9Z��]�젛��l��p�l<p$���Y�xL`��q~�7�K���\��,����w?��]H��?��8pҡ���dkz��M�`�4ϳ��T9��lbF[?K	��|}���٪�y��P��Q��$8��ۯ����.w[!�6�g���e�K��Ss ZY��#'1"�@D�~��s�:J{<�3��4S�NƵ��UǄM�v3�޻�b��v�Ҭڡw�t�e���1{V�ͤ�	�d̄1��\�ö��׶�F��|���$?��
�����P��<�Ah��ۀ)���St����]�q�F+ �}�)��6~?̈c�2Ӱ����}��Sŭ��/��%f��sL�J�wb4=��I��䙋���/{�c����m��jc��KQ���L�@-�zk�cT�ر���^28E���  q;";	[C��,��S]�/U�����d�QJ�&h9 M���Dq+���Ӫ��9�j�`4�w�O��xr$���/'���a�?j�z��d�C;se�A��u1��-	WG0Heɬ`��X��%�R��r4�N���KyS����Rtl5^.�D.��'��y�����l!��줥�d%��P�!����@�'� �bzA.��ƌP��Rm��nǑ����)�~u%�Щ[.��}�ds)혞GRWJ�
�(=������a����(!��p;v��=��1����o�K�,.����x�#G�O�Y�ƴ�A�Ղ��e�\f^*��{K�CC�\׃�G��و�C`S?�w��Eg��xͅ������1����^����2���I�>	%Y��ǚ��I֪�tyI$��<����|�	��B���@���Ӆb�Zq,�@J�DN�����y��C?h�2�J�1����nc�We���Xy��wn���$�`� ��`��"�3Ԭ6`��3��M�%��x����V㥜�7K����K�X\��4�픐V���ĴT���u�\�~���;�#:�S7b]#���:��D��6Ҩ���,����4U2�B�n~�J�n�vx���!4� �-A��Ѝ�'-i�.V�'6�	��a��:����䨾�9M�Ή�a�rnE/̈��
�!o���B��e��WLl�0@��L] 0�P_L��b:�B��?	y��ĶP=ݠ?F�,j�"��'���@��$��S��=�����m������Ң�@��h--8o��T�
�
9LZ�ؑ�Kz����?{q���d��)h	l*��5�N;_+Ƥ%��!����js@��h��a��-n
�Z����`����]����p]������\Y+8�=��]��&q�����^������N�h`~4��62-���?���\����kg/o�r?	�q�~i��w���l	&���bD�2n
>��mnD�f�'�?�!��DÅ'��X[����I�l/f��C�}s `��3�o��*'���ZD��@���mf�u�h�b��=o��fX<�5[ˈ�/�)��O���P"�W�UI�f���ֻ�G�4�<��R������X�ړ�׾ ��M���Lf������L������������U�r���H�"Q�v��g<L��f_ٞO3E*Cm�A]�
�:�ԘJ�����ug4L]����9D Ҟ���}]9�2-B	���
'?�C�<ݷ�%���V6�[�ev�$Uo�F} �(���&N/0�脖�������=�G�v��sn���p�����M�8�q*�z��N���(����[�J\�5��~:k1���ѣ�ul)>PE�y�ǅ��L#[5����OL�F�ߔ2W	:ō;t�W���nC�R'f�����7ι���G_ҕ��@��:r��v�����oX˚�^�R��
�o�!��ʶ���n,@�1��x��a�i�fň"��PY�FpI�I]	���| [w&�v-.����)>r��ᏏYd�� ���q1��b>'U����vOɌI��O����aȭ�Qk�b2���/@mkh��qi��W��Z&��db��?Ϋ��e�4���!P��O�Q�0jO���Z��qϢ���5IN�L��x���5P�C��#nX�Gÿ�5��"^cf��c������d>αג��L�����S�FXE5��0��S��T�q˯n�=�"��G1~����@tP�8�*�[/��5�Vl����5��+����<EuL����ؑ���UߩB�R"р>L��a����(/�1v�ir���t��3�gT��$ܳ����<
N\/'���f.n/�瀎8�����
����j�"y.��K���L��(�Z� q�҆�S��Aשּ�bЍ��'�i~B×�V�	j�F�+�	�T���"���񨶄�qҳ?Jd�P
�����7��J�;�D��%�PM�����g�Zv8l��3�y�љ��.��NQN�G{�:2q��e��1P�ذ�pW��˭ԇƢب�::#:�^��u.�������-k��&�P��@:����Ƽ�y�E_���zbU�} n\�H�窋�%&��aU"r�:�l:�&o�W��Ω%kR�]���~�ax�B0�v�"/��|���ـ7����=�	v̳s�0 �r�:�>���.�@��vSH��9����T\g{�8��.|�^����ǻ)|���yړ6��i�)XQ���*njv�Q��S��}/�\w�Vd��ųu+�Ҿ����+F�+��|2͑��-6�w���M;�d���;߷i���6C��p��k�mH*[K�E���8�P]υ|�uh7#�S�)ȗ��Hn|nؓ�	{����
��9؆g�(LCd#�G�|9&ʲ�o�ax��9qD6~��!�z�����|��h�쫢 H�q���88q��'�y�PC�ryΛo)��Ɇ���w��\z����}Rt����\���(�qr,~�BIu����R��+Jm��u�Qs�E(�Yw3떕g��&��|�����U|8@� ��sK�g�s�(���bfr�ejH>�ĪZ2a̿t��R�E1�1֠+u���+�2QOFA���!�g���_$ �:��nAP�aK(��JDُr\�6�P�1g?C)����`���Y�E��R'vK����q��Ne�H4Z�TTI� ƶ��T�L�����F�v�H_�(�~D��rH��ѡd��$�Wi2�ު��w����@0c�;7_��P4����j��R�;�ggO�_���2�B���������l4v;��)G8�|T
-~��DDH�:7�2z ��������z�Vd�I2�Il��P��D��ga��h�J�p]h���5@V.��o_����Nt_���~A$��s�15"�\q�{���G8��d1�^�"��7'M�f�͞*cT�;��hвɻ�¿rG,�y��)��|�5p��'<K���y��M?yޫ�4���c�u$U�s�	X��L�$��-�����,Sn4.���z���Or[J�4}iIK:;���@�BX�9cD��{0_^�e6���~PӜdl|�]�y4�?A�Jª���×�x����&�bL$B�p%��r�Q�1��h�2�	�S��I��<�d��d�4��S]����m>N��e_����%_��l���[ć���g�a8h���_ 6J�]�ę����6�C��=����X��6�C $ާ�]����9|�Ƣ��`o4�O�,:�F1$7o_A ��ƫ�AH���w
�k  ��M_��:��<��V���g�]ػ]Fot�������\57�ƅ���]���>9�WLCoF|y$;,��Ç���> ��̶�N�%R�j�$����U�˞m��fH~J�����eD��J@F�7?mH+;����)�*7U#>c�OEc^���������<�$#�n����'������N�}O��U:]E$!ߧ�<�o1r`~D.��>t�u����l��<�ݮ�<t����8���A��n�{\���)$�;MA��JV�PH�vy?��iq�M��*F B�,�!\�����r�r��)��v�h�5&X��w�L�1�]�%����(�D��ͫ4q%Q(4��!�-7�-m����$^AÑ-e��YC)���,�0{W">v��P��aqޡ�*l�i���=u�~�Luڛ�D�f��W>-RT�_�UW@��W����f��+����l�����/ �T�u�a@�i�ZF�g��:KB՗����!a����d׊3.�7iB]vhY}&2�,G�������D�������i��q@V��M�v/��5���twkmXD;S�s��,/�^�\�E�N��T��P�dp���Х�c��"��h���=�u����Ӈ�]B�b�^h[�hc*|�a��
*p*���R�h��|�(��bβ��!�|��ɘ����>��A�Hp�M�SV�!�3I1���ԗ	��5���K�ۮ=q�þa� ��Q��d��îH��<Ƈ�J�����_mÒ�&���ъ0�.Ivp�o�ד;8I�(��oϟ��I\iu�U5�͸��E̮b������f>�:@:�L+�U�Ú����y�D�Ŭ��-��y���g Sz"&nt���)$@�yY7��y��|`�*��"��k��7~SϪ���\��;g�)3}���
��#}�Χ �l丬��K����zSN��*��7�`o�u t�;��E3�ܑV����	f�.�K��<�?N3��(��J�
9	|s��B �6�XmMH%����?��d g���O��h�J���/��x���g��z�K	�z	UA�&5jϬ�z�=L�0���&g�5Et��E���w������to3E]&���̚�0��<���_0���j��f�� QN#���@�Y�P�C�k��
�" <��}�n�Q|�dg��������WKJ�9��]̒ߞ]�T�/���;z�I)��������������5[��=]�_6��Jg���}}z�64-�ۺ[0�"���C��'9Q�W�����2`�� W�L|������_��öA/.�x�O� �b���94��]׮�l�op�\6<,�lH΂����׵���������51�B~w�be��~{g�d����N����Z�;T4@[��!��F{y�����֐��v�s�F>=M[p���5���oMˤ^O�AƐ*��`?��0�xｺ��MSĩ���$0�u�i_�ŀz��X��r�:U�{"jP��ĺ̫�z��ڿ=8���At,XJ�J���� 4�Qyf�5�ﹿ�h�%׈�N�|��f�}q�n'uFX'���$$�J{h�X?�b6�x���~�|a!3b��x���O�u>l��Th���Sţ���,	�߼�2f=��5'2�5A^/��٣؈���IY~;NbW!c�������lC�V�*������Ua�aЊ�
�R����5�:�X⩰N���q'���A��Q�1}�]�7#8��VW%��H��}�VDp�T����7!�*4�B�_&!+�I9���,B��U*�AY��I�ȕW;�*W,�[��A�IT���һ+�X�� 0�e��ž��=p�B����7�p���q'�å�t�,(|]�.S�nz�1*)|��Ԏ�?,��aa0!P��8�ʉZ�E���\ ���6䏺�e�)钦�}7}���_x�a�3Rb����L�����W��w�h�ح�VH��\z��%
lMp�k�3Oi��Y�%�=v��������"W�H2 ��fӠ�@���e8�B6[���>�!�����]w���{�k�g�8${ȌhV��B�|��K7dI���T}�^�pJPn�U�*��j�d /EӳI坦�����)���"z�Z\�]�M�A"%��l��2��f©\cS�rM�+�͠�1eGN`ȋ*�#���Uh�Pl���E�Q�ݦA���|1�HQ���-BE�į��()��N΋���@q��հ�3�礄Vd���c�$�NԐ(t�S�دc{R�ځc��>�\$8�ʲ�k�i�8dd{7";Fv�C��e[���FXnj���0U�5V��Z�S%z��xrм�^4�F%Ri���|/���a��Sb�':ޘ���q
�2r���ټ.�������9����_"���>g�Ǡ�%Mi��o]?P1o��\���"��K&�zT�>,:�&�ð���)<ugʲ7KkF�e�+gPI��	o�|䂯�S��2@�&�}C�)3�;{2����RO�G�(�z��t�Z�|O�]�`~#۶"gr�J����f���@e'��ٿ��q�����)�bGV����^7����}�UC ?S���\���8@�S�:\�e~�䫤�o� Tݖ�1,���a���K��}�Bu��c4H��$�����eC��k���$'���S0&},W���(��ZjQIP� ˣ� ��B���%/�E��{��a��������?�a/���mُi4�� 1����\B�Mp`\K����NU�Ðh��qԷ���#��n�e�E2R9�V����L^����f�U�s&�����P��Za'�pjh+�����|��w_������������LH�<�7��l:�hǢbN�I���r��{"H;�J5�ƿ>%�>*�{�g]sN�\�M��r�}���9�U7]��+�֬@Y{��[j���?,�y�7�(�x
G�ޯ�}`\^p{��;�q$�c����5���f���~/��D:��C��_,;!����vг�_��y�O�#�@� 7:���9D�"�-
y	�Dˠ�hOL&��'ì�ܣ/���Y��<˨��>�k��j��誄����"4����߂��W%��޶y93|j�G*Wb�n7��[T�*/�:���qS��n(����E�X�?��R'�;�4�UU1�<J��v��换K�&��wg[b�� �?.�C):�W�>P�_�q�'�<��j0����8Jl����"	�w^Ɯ��ݰq>�-�99�R�*��+�VYO���`bF��%���O ~a9���/�)��Gӎ�.��N\ځQ�cZ���g�}9Ay�{�<����;����Dy�bd�m�@ˌ��9���`��4.)�#א��]>(-z(�Y2;k����&,m�
3�3,g;��o9c��E�w� uG8�j�\E��#;�{Wc��8�$����;�cx�D�׷m�/CҰo�w��0���|c���{��<]D�U���jt�&[��C3�hc~Cp�����[%!���z������ԛo�x���'�Aj�E�u'���ut��3�~�1u�7A���ܱ��E�(s�&��Xu_2l����{�x<����."�[㌤�˞4��� &�v��miɰ.���D�J�,!m
�u����8t�	�C�8̹8��[J�U�YE���#�dP�e�$0hj�Z�'���7	w@D�Nw<��D6�6,�J}}#��>��J9��&�O�e�OEA�TA�����.�-Nt��ܿ�w�O^�te���{=������x��V��5C����MK���1"Bc��)X�h4
���9]t�yR*��fmq�0��'Y�KW,�
;�8���_;wW�,����h�wa����0���6�*��xE0��/�U�Y�"�W3����y/Ǫ��T}|?�pJ�gAm��Cbm]�ȿ����EI/ŋ|D�-��NgǊ�	�8��M�彨�i��Rئ)B"Z\�f �uo]��婧�ۇ����>k�����$�u���yu�g���a(�3�0<���*6���T��aU\<f.U;��/����]�m]ۣ���"U�G;�]擫4��HCZ�`��y'K��%m��c�R�iN!�c8��3f���W��?����*x�����#���Ec��Kinto�I��#�$�A<�w�9��N�2��+ɗEˁL��}
�-8]:���H�S<J��jN% ��V	�d;dU�o��S���<Q��,�^Xu�3�64q!������3��j��3IމZ�D((�j��]���q;.N��J�M���MJ��y��Yω�ܖ��~L�_A�
�m=�?�������y�����/*��~vm3y�%�&t$�a�X�L�a�P�D�6��-Ⴂ�t�V�b=֪8���퍒�.�׫Xo�-����8ls'�f�Q��8sO{��ic���]���i%������fC�&Hٯ�ޝ�AS�?��`��y�?�r��82�@�	�J���z�~K��8�Y�*JJ<vǍY�>�^����d萪��Qƪ<��e⌌SQ�V���o�7kMtE�� �Ѩs�"zd��d-G=���t ��0��Ec����;D?����������V̥g���6t��a��]JTkR���쇩FZ���&�$M�Ǎ�f��G�L��~T�凾��8�t`�����qG�	iy�N%�#�׫@&��"���ZΦr��rt�V������п!w]����˲���*�#M2^.Wh�l{�>��'w1:N��c���{#�}	,���pM���/�S>��A
���SO�*CT������t[������Z���a�:��x#�HiT�WW-2e��L#uA�=����&̈�IYkUN�%�Я�ʒ���'��e�q"�a���g���6[}��h��ĉ�H�\]��'�,��p
�7�	gӞ�z�0���֪���gq����K�9b���+D.PY6Wx�@�5@4
�TŔ(x�Lu�Zt`�� �_�#g=?5�\�乪#.��j�K{�K䨖��n�D�
�F����ރr.�a�'G��l��ga�*O� �g+�b��NMS�J!��C�$b�ݔ�]�~��l���C�c�Mi�G}|g(�r��ۃ���qU��;!z�+?T2hA
�S\�x#5������c��A�S����4g_��#�h�N����X���7An�ӎ����&�6��~��m�K��?Qܪg ���2�m�s�v��rB�l,�"��N�#���{�x�yA *�x��X�w�N/Ah4�z,4ԥ���Fm�W���%����*
J0��dd-�}V�z�����5�쾇R"��o�l�N�}����|���!!O��+P!��s]���F5K����l�A(ڠ�=n�]�Q�������0o���u���EM�k�������pJ���'�LkDlQ�z�4�w�1g��Ve��ٶ�e�k��*�u��w�HZ!3K�����t����q����"$%P���!�Y�i�͊fT�Q�I���������~��(��l"U����/�0d�y�X�j�e�����З�K��=yƁ��A�$�W+���wv��8ы=)��i߾;�/&BU�+�p�����}��#����d��I�n��{$Ԟ*-,`�CO��=�{�n-�;}����|��;wD��89$}���<[HHx���PgP�e����v�.�8��a�z{�<m��#���8����VC�=�<a`[w���Ǧ��@���n�>
"(Ұ5����@���>yHϑ��T�Z�P�r��19���m>yB��j&�('vgx~8�b��/�V�pb���o�v�
���r����� �@��S�.�� ���/m��`T�}���	^��Vj:�Կ��0�-��v���[zZv9Qi��8�Y������*C�!9<�Xhs93d)�v��$��}�)�g�|���}�aE)�º&�W�KȮ9����q�`��[�N6h��+�b ����1:& i!ڶN���ф	�:ַm6 � �3]5ܚn���H�~��nz3�\@,���D��N]��_����R�AV��tfn��׋�#�;���D�.!L�,��0��ːw��.����ԡ��1#�Wpj���GV�r�I�T�ܒM��-�ѐu�L��X��L��s��.�g[���y�����xI�H�gz.\��U8��xY|/\d�+�_b����-tv�Y��v��$:t�X@����D��q�1es��+��ki]���s����(���>��&���C���\K���ŦQ���ѩ�(��,ѫn��D�y��O�^l�b{@��!�X��W�#-�a����Q������s���c���ح��V�͹�[�*���������7;)��l�Q�|�@D�i�T�j	
���x瀿yOϊ㕔�A�TU������;㢭t;sFK5���vŴWC��v^7��-�I'���_��X����]�b�h���� ��te�E��U���$� �](�mqw�dp8JΕ�(W���I�ϓ���Yr�j�>�I'e͝xy���$ڕ��G�=�}�@H�>":�\B��D�9B!/l�!�n��x�۳�������xO�ߠ�%i�C����.j�~�+i���g�1�V�OO^x�����z��H=u��$�c�����\+�>����O��	d��<�l4rJ�5�@��P��R��H�-�Xo���'J�&���Kۏ������`��M[>��Sr��E<P����A�$r���*o�	^���Pީ��l����:E�e6n���d��&Â�A��4S��;S����R����J�5��fg�u���A /���eL�M�
�L����1{�9�7q�^��f��J��X
mt��<A��{�ni�.~Q7�<<#���G���#q�c�`=ݤ�_c;�m�����8᧊G��B�(� W����.G�n^N�&>Xy�pw�G����eyy����l_�a�}ξ���A�;�������$�j%��8��;Qq4�}d3�n������Rz7Rn�A1\Q�BE�|q/F�8On	�j,�3�m��&�c��zeJ��4*?���j�3��>d�뇪]�{����LQ�t0LB��E`dd���eěH
�d0��j��+���ӡS��1M��f��d�%1@;�����,BG��[����(:�A�g��JK��g��	���W��
yǹ|8SG:�1�w�p] �^C��k�WƑiWe:r���E$Asu�M<Xj������ C-֠0j~��g�jq2P�9�4�������TҜ��$ȶN�;'G���dޫ�w�f���Gz0�M��n���!>�K��M�E&%N����Bi���)/��w]Ek�v��7ܮ�$ɾ�+ڈ�Ԗ#ǌs`j���X��pctt���$��9b����i��a�74J��=V�����@�>��r�G]�/4�Ml<���AA�U�^q�8mhX��	���|M(?V��T��:�@�=c|�r�f���a�a*єߺ&�0���2ma�A|����80 �����	��2y�߁BLP�W������a0�g������4���A"��L����34�X���̵�z�顚 �������9�󆳛PCJ?�A�5L�~4��wq���[�S5�,X�v���m
d~F�R��NM�8V}aq������2t������۶ͭ��;k�	&� �7>���%�0lK��Sp�Jp�b� ��L:��G|3�j]M����Y��)P�S���;��H4����;�'
�{�WNW���m�
�AK^����I����2֑m �C��!K�4��i^5\t��S��c2��G�jwdWSR�3���B[=@7n:{���ӄ��5KҺ_&����;���d�_�X���>�~	R��4^Q���_��ӯf�$C�g�VhܫX��xn����ڒO��X<���E�3.�ĢA�پ��Z^�مE��.�w%N���n�ϖ%A'�0h�xG8%��R$�ia�pd���{��2�������2n�$�h�P��m�%q�Ǒ\ �GS�P���<�:p-�;t�AM?C���� Q��w�*uw�]Q��}�%�K�H��n��VM�%��$ɾ{�tRM�^NI��Uҿ:}X.�ߵơ>��vB��y��s"�հ�7���HfZ�*�|���k4�2b��3"����Ç�+G�20�NV��ĭ��O���e��U����Ŧ#���>9������G)�@�����D~4��?�ĸ/��OX�.c�_�
�w��|����>�Q9�a����(�=p(n��!��t��ϵ%���33����*D6W�����8�=��f�LX��ϊĖ��n���cf:q"�O���f-�����V���WSz�ҌHcP���!������q��/�G��	��{:x[�Q�[��edԿ�ZI�ŷ3彖m&�gj,G	Ԁ�)��Х��D<svA����x���>���#'t� "Eu��XKس�xp���&�%��-A&��;?�^Qm�ov����Ȇ��S(��(��n،�j���s�H��PQmвN�fh�u�2�CTk�����e%��܉Z %��a|�x�QIx�����8����?��;�c�I΍V�d�Voc�4ِ�p,�о^��5�;�n��!�5!Ϋ����uso�b���ff���^uO@��%��R��!�nk��I�)Ս���X#�?���yv�Xp�<r�ɹ9����� ��@ɸE�Qj�+�O80�%z�D/����h�-�CmE�'�=7���:
���L�)�%"��n�A���CFS+�(^�	T�/?��$��ϢAo.���}{a��vXʼ,�ڒE�8y�
G[ֆ70Qs�Be���@��BV������S�n]����!Xx����f��JQˆ�S��������/C�sw���,,H������E%��G�*(��}d	�� �馨e���t��Z�<RE�YT����.�h�_Js���t�,b��,�3�I���`�RB]�﵁�@�����M�:�q��_����7
���������5̄��-h��L2��:�KP�-j��s݃���8�П����Rp`:8$mX�Zcc��D�`Y�=P>��d�H�ė�}by����f�e�K��v�#5���0���b���^�&�c�O]���ʃ�� ϝ)�i��}O��qX`j��x:yB�����婭��GXO��KS&~��v��g:�l`ǹהrjSj뮔�mǣ�w���*
NP���?Z��3��
J>��VR
c���
[T	e��5h^��n|����`���{;C�<����X�d������J�>��	gxr��K��⤌���t��$yz(�.�pF�������R�s$�ݝl\6������<�awt��d@�Lb^f��z)�RC*g�:j4��"�XJ�U`3򇩦3�I���"�`�s/^YMn]K�.D��&?Q�r3yeN��6C��uw!쵨�Z�υO,S��P�ZT@@�(�2?�,N8LL�À�v1�U�y�Z{� ���0v�(l�t:�n7`��=����Uص���͹�F�P��Md<�2�����}���<@Q0�L��Y��ꑤ1J�ar�~�M��H\�#M0I�Y��r��˜���1h��&IE���P';!���2	߬�Ȼ����h�ܯ���qX��#��
��7��ћ�HAo�p�Q��]C_�3?�ԥ�������	|e��ee�!$�Y�B�&�A�I�K���7��xl��V*��2�U�GHٶ�(P�4���2���c��~�V��[��:��ʥ�T-��?+.]������c��:�7��>�p���҇��9�CԠk'\�p������mp�{ [ۡA��`MBn(H�(l.D	d60�$����^���1Q�u�u*�7��vv�>.���4,;l ιk�C��?-��(SR#��g��)�Q�wu�W*��_+�Znc虫���;��a��Y���2rj'�gX�%l!W���
i�I/���L��.6_�*0Vl<,�ћ��������^��F[������&�vT��,�n�mܫ���Nu���� ����_�ܜ�$3����
����_���$d=y��ig������ڮm�r���X[Q�k�����B�����b=��ȉ}`����r���!E�m��+��	$�����|�@b/��ٖ=��j�������²Tr+OPZ��z�SO�[���Y}d��06I��$B�y�!�XJ>�݄�L����*V��#gfJh��-p�dAFi�΍���~�֡(�G�ڕM:Hl~V�>L _�Gd;���x���]����ș���u:��v�h�^SC��`i�U��v:)�[�BDD+���"z2����@ Ư��$lSzY�tDu��gФ��m�u���N�1�c�3_�3,�� �v��{�[1�.0����S��H"��LKg�cd��<;yȁ�7F��\R�i�C���Io��W�ץc��l~T��;[�s��zo=R_�Bԛ2kc�~�_���j�o� �����n����L���Z�Xat4�|��G�$4jU����>ηf����E<Vb^�7��EfG�\�1 �SP��"'���TfK���KG2�� ���ڤw�����u�@$֕q9�Y�<�*��y�=�W"�	Xte �9�2�Xa:))���1c]b��&�s�sR��ݴ�ï�/� ���pF�qOi&�J�Dv�/;9���'qK�j�MA!�_�1õ�������P	CTٚ�<�iV8�0:@�q��,����ے`�2� ���D'���*�!�!�� @1Hc!����p���R�m���O�I1��6��;a���[��,:Vb��	�/aSJsl���nK@d�mЁ���u��3���س.���!o�q5t!ONi���;:g�.��Nt��B��R���6;[ʤjd�f웵�Ɗ�h �X9l��C�犭����1<�!��C���(H��(v�*� U���w�Eb]45BM�F U̬�lx�@�+�0�GWd�n2|�X�\���6W;Iu�wp�dd)?m	����t2�rp�:%�&Y��[��1(틑y�q���/0g7��^)�[�س��PV����&g��d�<�[��S'��TY;�.���EA*�_B��W�4u��ś���tE�_g�⏋�E5�`{*A�R�dT�߯*�N��q���� ���gK��A�S11VW�,=�@��	:���0���4B8
-�B�fv�.���p���`jק��Wහf���i��V�#��G��'�*[�,��g�X?���{b��
g�����F"���r �ϩ������������F��(�O�~z*brhZ�Ҡa�s<>�]н�6��ӡ�Z��@:�9|7mg���5����[�o��[�]�jw;�t���uc�h�apХ�k4��|��/kjaD�XX	:x�Q �P���-��X�W;Bĸ��u�� �a����WQuE�c��e� ��g�;���:j�[x؀ggb\,`���ժG@\*A*�ۀܙ��[l �"��P��Gז�?�j���8|��*R$� �^���|�A�M���o�S����^H�][�n���]��:"!��;R��2��$z=@:d�4X����aB*������Qº|:�J�#?����Có��Er�V�'�T{�t�?�>�)1�!�Of�W�|_�i���M�5���s��ǉ�����bcbeb��A�����4�} �j&�`�mO�uQ�Ae�L�߷�O�N����8J��y�P�~G�z��w�F*�٬�����c�h/��{"n�8D,vsv}����R%�1�+n{�o�@�'f6m�����(IۯѮ�,��{�}�g�;)���r�h$h������Y�RR��o2�Ѽ&��Q��b�����S޽��@�h�O�#s��q��1]��Vt����0� �gk��:'�EJr�;�dᏞQ�����z���@n�}]�Y/"�{���-�8QL���'�F4�8W�zc֔'c�j@�I��j=���]1'D���k�
����w��]��%l��u�jp �sH���S4_^v��b3u�+�B[aZ��,r��W�%l9]�X\t൝�T���N �Lա_�8F���=��+�ɷ��sA�-��-����@qA��x`���b��7 sD}�t&q��;�r�<Ұ8m�Xx,��kV'�"\# V�f�`h�}-�A��v)��<�rl$ԥw
F��}ã�xqNB������Y��t#R�H�J�}tL�->����.��H��aTkW�8 �IĴ��;�t��'׵��l��R�9���	�W�^T�+���7�Q��̳�(��
/5җ��
��@����1�}|l)�e
�[�7ڪI�Ǟb-O�/Ãl�?�6�}�b��d:Dף���QA�����q��z}b9ꦡ<�m=uδ�w$*:�h�gg�V��7d�2���m8�vR8��s򕠵�I�f�PE{h*pd����c�,�kz�y0\�8#�I�0��{M^d�xՎ�V_��V'�;CV�1?�sN�-�����ucF�y$6�"@gg2�Z�]�E�c5J5�|>�i�Y;@�J��K��-�wER�W��l�Ty�����A.���LP9D0IƮ�t�� ʋ ���@@�ْ��쪠�`)������(8s����H���gϘQs��ߤI ��&b-z���{�N#�{ci���)���Jדұ���I׵V��\��ד���[[y��/=��A?�76� Z@TE;k�1�RϴB �Rr��lr�p�|F��(���4�2�w~�4���L#�4y��̅�Q�:x9ff�`14�;R��艃������`����������� | �N$Ň�5y���Mgs��>C����JSSlC��cH xY��<� sA�E�k���;����)���Kڔ:}�R|H>c�?B��9��W��f��+d�0��䂞�N����E;�I-��%t*ȿ��	���y���)!pOW��<;�FV_r�Ƀm>���1p'�_��0��%Wu������A'���\�'Q�߄Ms)k���s�<�������6�В>^J �uR��F4�����W��	��L�l{j�1L�Eg(���*�f!�ڒ�%�������`)Yg�2�m_�~��c����
2�!n^�ÖRD�p;��}*ٿnI��ǆ�e"V�^6[�H/]����Mv��I�`�w��*z���=۱�&���Q���͑z���_vb���4�� 1�B�P��%�4N�<�ȴ�����SA���x���gxzȥ�s i��Kf!�G~$�e��ʣxzɃ�=�{+�dtsӺp��¥��h劉����!b�YuHYC�Zc2C�F�ѿ�?"�R+����t��x|��J
��,�#���<�R:[e�������?H�k:7$��
e0�C�\��l��/><l���l7l�`! �	��p�L�&��q����N�!#��
^W�[.@$�hK,�4�^],���d�_7���%. b�누^H1�Bz�TكE�d{f��]��L�}���>A|�N�7H�� ��rqS�;7�b9�i���@^���&"�I��8���{bV3TX�f㡒C_c�e�v,p<���6d�
,${&Eқt�`JDx`���v\v�*aR��yz���B��Ǌo^�����Y.�X��G﮳���5��VU%�në^�M�R�%VW@�V��W)��:����!�'��Y�68�ɷ�
�F�W��Ե�*�D�5�<�?��E$Sk��&��H���#�i�n�?gP-�;:����ِF�~�Z�M}�e��>�%/ze���j4�mP���駲�%F�S��D����������\`h�i�f\3.3��+�^���AL�b
�X�8�wcѥ�UA��; ̗��*���]�C� ��ۨ�bS�
P`�V����D'+�H�@�D�z��d�c�d�+��	��c�o-�7����ì�L�/.		�3�ml�!������҄��6����Ę�VT��h-ǌKU�7jң��q�M�+�F��oO�����mR��`��]ӿ!�z��%{�v��9A��:��Vv�3����M%È��C����}�m�)�ET�`�Y`K�Q�f�C��CQ�r/�&�$�^���IZ��`�G͠Qe�w&%a��͖-v؇�w�b����F�ٕ�E���ܹ��wv�ܗ�0�
c�Y
1�r��G�epW�8�
-�G�Ԣ���c@ؔ��sRb��'�v]+�"V�p�15����i��F���ǅ�+�e��u���Y�R��d�Ir�۟of���?��ʚ�ъƶiE>�:l���u4�v9��"������Pu�N> 7:��]ei-��Ә��.����`�E9����^�;"��������v�8�J��lr�X*n�P��O,y��L�{�����F�8~���y+_H�%j	\>Q�.�2�^"��.��7�� w߈�ذ���LL!���a&�����&^6$\�=���<��d�H����D�	�q��A]2�O�4����t��Q=�THw����o�/ľJ郥Zo:��Oc@����1rF�����I,���l�,�I�*N��- _�-��m./���C���;4{r1���36��i�9��p�u}�����q*r�L�$�i2���ÑD"@���)$Ʈ��xhdŋ�I�c,]mo��ClF��N�T54KM>*�K�p.��k8��?+�*���N�p�V������B�a*:VVD ��<LQ0��9CSt��M�<?(��gb�#�N�f�s�vt7�ї�L5I�G�x�/��\`H2R�'�GQ����!*���̝	Ub�k�R�i)ę2/�����_�Zʫ 2�x�f/���>��nPps���fv
���D�z*nA�8����nl�M�^�����������Ɣtr]k�%�O*��kX�����*-՘:jT�qޯ%yq��/ΉiHNJI���;>o��d��o:]'����E�EZ ��������;����Wф]�tHIYf+�GFP
�EN�s��8�P�)濏��NY0�{��U�q�~>�� "�E����q� g�9�	B%��D��C{g!��\C�ݸ�<1����]�{�x�h�lP��U��hj������ۿ�q�>(�<�o����.S,V��FUp���P'o�
�)���k��^�WXv ���4	���y�J��0U�Y�(����d���U��k��\J�=��>
��:�wݿ-j�3ӭM��nTF8�,9�X�;��˵_�z)��%�Z�N�g�	F�L����Q!�߫�]ɽ��׷���G��y�@�+R
j��(����j�x��ɞT�ȼN:"�dz;�\�E�*A��+C����B���@s�.>۽���������/��,n�z<v�ؤ�\��4�T��A˞Lu�4Sf�>�hL�=b�%f�:��:/7�������N��!8��	ǲ��;Ҫ�6\?)��m�6���^�%�2f�)�>�,!�AG���"��}�P��;t�avLZ�^�A3("B�}5����D�6N����b����'�����T��g�,6ad"�h�5_��u�!���:���͸W�.�f�V5;��%P������h���@NC�+W\�C�\6���s
�	e�=}']l�n�=�C3p��:��	�DzVg��t��������Ik��X� }��>r����C�]&Ji���z��]6�D��W����ĝ��~S��nvcT�W8��-H�C��:?�C���XS�}hZZ.`�*�9N�f�d�x��NA����Y��T�ҭW1��w����t\��MFW��ދK �A�$���~�gv�h&?�>w���� �}�Mg�梉� ��k��|�G���"ze�H�A@Oå���>;�ǳ��u�W�7��!�d�^:�9<Ӆ�*kb���pd=�3���	���В�D�	��b,#�+�Xf�MT{g��Z�u*���N�l�z3����KQ������3A��!�;��j���D�:�b3,y	��*L���.?|Q�J�cq$��t.�0�k{IS�
EǴ��Or���s��р](j���v���rGٸo`��?�P79W��%?�Ni�
�������!���>���-^�v�f����E�Ų/R����/m��S��~"4�s��	�U'��]�#��F���PϚ�'���_�����}޶���,�1Y�0�<e\�����a�=x+mpc�tϤL��w�0mA�
)�ʃ�U�t��!���Ͼ��I����O��|�]�(OL_�Xc��k*�ӨY��Y�zʺ�q��ce���ˑ��3�\i���]�KɊ�.1^���%~X���Ăv|
����?z���@��[�uhI��4>9�c����m�<�IZ�߇��l���cy,�p|�`x˯�s��fX���k�����n�{�Vg�88���6��ႛ@������x�&
�����-�A� Ai��e�� ��؞�t�JE5G?�^�7�����L����1���H��߯��Nֳ�kRA����V���򆔄��U��D0v��7��~J��b���q�B!=���v,���m��]�
FW9S%%!�f����UEu�E5�P7�+����xט������f��EQ��x���ؒ�/j�lspE���*:%�1x��-��Y1��y����Hу��B<�g����n���A|�����V�3��!`�q4y�3�R�;��K�X��m�ϧ��
X������ډ3#됣��S��z���E��ԣ��QN��H��@���-�N�;�ҭ��Ջ�f����-,a`c��3��U�w�����r���?]�H-���~���B�GsW5RV�#��2J?b�z6�G#Ų��4Q�4�]�����Y�a�ɪ1R�;�*[@m2u�x�g��9̡���>��H����Ԥ�~�r���N�I�Z<�W^ ���5��D��k\���64�e3L�Ч9�Q�����V�Y26��gS�(�=�J֪B��2��Bl+~�d���_�ֿ����F6�=`�N�"S��X�<�@X�B�R�W�j�0�*����)kj�D���AH\I>Mc�G����w�ǺA��y0��l.?}}��R���p����=�����T�NBr��(4e����F�� �zI�8*%񍿓r'�k��tY7X[@�J�t��5Ϋ|B��Eg+��C,��E� ��i.�NJ��-yE��`7��O�ª=Ī��ҭNy�f,%��#��7n��'�n��]���L&9ڦ�w���r�3������I�E|},	���[G��/-R���Q>4SvkI��~b��(���FL=����ŷHx]�-m���	i�2�L��l�� �O��i�)@����Р��n�����v�15��[�ݹS\I��p�����O:u������v�¥����3TB�;hϬ�t�gJyH�wD;��/��5�+��[N�?�&0��X��6h㵬�y��ȫ����P"uϞI!��?�F����%$q|tH=���]k4��]+�[X�'��vK��r��2��0s�8�*K-)#J@M�����)�E�X���k�F���'~K 2�vv�7zMS�1E�,1�n#�����拈��N<}��lJ����R��ޓB@>�>� ����x��T	9�g�a,&�'\u�A�6V2w��P��x&&�}2M%�ֱ̔w����T%���䅏*�[����g2�Y���(s��/������r>q���b������7�
�c�ǳ���>J�	��;��\m�:�"��Q�kQJ���9��T*�հJ��(L� �=������E;ef�d~��~n��$��"C��d�},����J!f���K�����r��2��֘t1�A�����Ƿ�L�` ��.�>��ͅkY��bH�w��x�ahꡭ�C�X0:$Z�A'Y��<v����*�a� .1\��8Cw��æQō�_�b~V)>%��z�ƴ?\��f�wx��Q���E����;�a�L�dz6Έ`|9U����/Ɇ�����T���Jb�0j�Y�_˃e�#��6�\ZR�8�h� ��8/J^*��� �d�P��!AFV�NU��Q�
>���D:�Ep�9�ؼ	E�q�)���ү^���d�o1�-��!_����{�y�R��^_cJ��$�����E�n�¶���7��bo��%��������C��n������9e���c����c5,����o�t�H����41����M��d��`��#'[���H�WF�z	�;�t��J$*[����%I�?�%/���C�Z�,_P�p��$��D����X�)��d ]�N�E$��(K0&#Q�&p-�eťd���\M��q�P��=�z\6,��U�EE���P��F�(ˬ�{�S�UXqP�o6d��u`��g�E�,Ɋ��Pz��g�/�Q����vײ#��d�p+豦�!m���	��h�:����������-_a�ƩJ<-Q����.\��LVF�P�jw�Xy,�����a�MPw�L9��X��l6n�2�u"?��tu~ �PD�(�T���#�':��Y񥀓��C�p��ۺ�/L�S�� �w�>cyТcC�	�g��������/��=ś阰_� K�;��/��%�W��_B�g����̒�t_�\�cӅ�r� FKJ:����.뒧��)�듶�$3E ꗿq�8K�~���Ap�@��[o�f9Y���w��7��oU �b8�U�mŲr@��n�g��S6�n��(�M���"tf�]�%��|��\�V�h���TLv�<X 5�E�<�j�a��ꃋB�
M��G��9�E��m[������B��"Z�М/�����3�Ɣ�o�)���#��[$�m�r���ݭ<wz�����?�����wH�
����о֎`_5n[K�8|��S�J����2���X�?�j~�y�k������b�`7��4��v��#�U���-��q���W�B1/��z�5��Ҏ���R*��42k�$�����Y��U�]27��]�~VJ+�����������P�#���fb����s���U?ƗH�1��HL�3�����#�]w9��ޞ�@HN�Ol��`g9�?�A��D��Ô �d�qe�;���t�Pp)�N���|X������a��������b[�J�Z��KB�e��Ξ����j6Pk3_CQ�̹��́���z�d#bɺ���Y��3����i�X]|�X�z ^L���Da��bm��b����4V�>͗S����si#+N���X�w��9V:��ď���Ks��e]x��KO�RM9��\~��Gԋ'�؜xƺ�Z3hlW��f�ͱ_�Qm)�eP��{�,��-x�-V��[�]y��>�#K)�dC�4��Wx���+}
u��e6�����2���᧢Q�qڐ(UF��J+,m�$ݧ3<�������!n��o����\���ㄪCrJYm�9���0�:�me�<�61�dҼߴj��l衑D�(�u�X�u]=�q�{a٧̯yّ@��qã*|T҄�q���{�j;�68B�G���F�ș��
?{����l�����n ퟸ���¢��m�߷$��h'���-�>�+E��'}~�Ɩ��*h�\z��#�G������8�-�2�=y��{^��Śuq,�+!�y�Qod�rъD�C�o�>���j��ZB�?a��ք�*b������\؉�hS�B���b�2ެ����rk�#��(1l��B�k)����3���:�WS7�EO#�c%OPun	#�+B�w�F�'�\�܉!����k�"P�^Yvv�!o'�JT�@�*dj
��pӹک�������ʤf�-�X��͟*�����ܴoEo���ֈ)hBl���c�g�Z8ѽ;��N�:hn*�6���9Z�L�K���m��F��
���E�p�1��6�W�o �`�ؚ�n���������{�o�M�k�����
i*�]�5���t�l`k?c(�g�w�W:w���'��0��&ku�e�
h��J𖞍�]�[�?^�%�����	����s�g�ԙ1�ha�	<�=�	���6�}9ґ� d�>#�sm�5��:;<��qCā��z&g*�I�aEi�q��r��'�i)@�<=p.���P��*_Z��t���H�/�lo�`M��T���П������6C.��*@�hq��Ӽx`���e�ANCy`@Xp` h
����H�KlOfx�B�1��+p��~�J�
���v�Xw?������\��L���P��MDB����C��-�@a�ZM�(0+�I�^De.Qm���fs�/q"�|(]��i���s`x�x>jkqR��ӳ�d!�tɼ�$����"����:\��[���%!.��7W΋���,)��!!9��F�_"�7�ɉU�%>��VDD]>�&���E�� �6D�lO&�������5����P����8z�Sߠ\�����z��a׸��c�.�1"@���d����P��}�[���<#Le�}��4]���k�>�G�־��֍�υ�'f,�����Θ�j|A�wwD(��P��z��Y�L�Z����`�C�+K�ݛ,U@sMs�Z�]k��96i���p�q��#q��L��d:��}�K�y�p�$�	g�}�YK�_�{!n5�Q�������2m���[��m�k7{|*'R�'�ί�� �xMv��6�y��k���.nP�<e��yeK_���I��nv�bL�@)�h� dJ������2�ݑ<���s��4*���]����{K��3_��n�N+���Ȓ~O������I[C2�2���7�&��9&�B�Ah}��*��!�B�P6����Oq��'��S���>�^����f\}e������I.�^O�z��ΗӺ����t�#����|R�(�����v���3��r��is�O��u$�^Yt��n%9](z���	��4�{��Rgʔ;Gc�&E0˗��!"�(qvΥZG�)�J� �LA��Yf2�<P�NO��sڂ�~����#��*�[9��4I�T�ᡌHyYoHX:0����'�z��f~{�!T��0���7��Ԉ�� c�E��73��#9l|��*���f��@Rt���.���)Y��G��bũ�cH}))���-S�+�ζ](��خ�To"�ٓ��$a9j�����&�j8����#7cX����r���l�h����t�jղ��0�f���=���KQ�9<�{b�N�񃲑a��,g-�+�//S��S�}�����9��m��FR��6��~�����]�I^����2���A05!��+�ūѥ��}��[�	yY�h)�\�im�$Ĕ$�N�y�q)���
�/l__���)-1|=	�!�?�f��6`�ǏSh	NѓdD�	��v�p~�h�x�Q�#��6��!+��E��/:S;&�v�ngs�䯛�!�iF�|�G�,�²�H�D��L�N�ɜp��yމ�ɺS��(X� �;#3Q�l��c��,B���4#z�-6D��C��t��0J	�J҈�����e�b;�3��K
)�V��#mɮ���u��&�
�;���w���矷w��-�����@�$OX>x��>�0	_秭�
�j5�ZP���J=WXd��}ES��E�!V�9��YcI8�7}��(5.'�.�0ۖ�2@������0܏HL�`��>�kx;/9ݐ3��5A�}��Js���þ(���u�7�b�������::G�q�9	52%����2r�oj.h,���*���Igc���I���8��n?lZ�tU����v{�Y~䡣���F8G!8:	G�q�����ۈ��A����[��z<�������']�6"p���ik���p'&�8��Dj��	7��+(��+�c%�Y.R�@�)ws��3����7FO�r;������]�8�x�N7�^2�S���I�5�a�p�.-�x�ۜ�zGMS'�I:��!������/�B�9Z�=cFŲ�U��=��vk:�g��a�����]�����۟�B���!��'������������uF-WnWu!�ﮊv�}�
�V�<�E�������y�8��s�����c��EHدԝ�8'�X���5ԙˍL�Z�_Y�N�b�'g8nD6�T\g�Q	Fvse��d� IX��C�p�ı-l���T��Z��Rcv�&������o�_'��q�Z7nF��u~/�Y�.��p�z9Γ�Y$!X�B eDf�Ǳ��i=+��H ���[�hr�v:6��50��!�ݴ��J�o'Ӥ�}�Ȭ�~8*����!؆<�C�toM����A��2O���,�q=&��fv��>U�l�̭���X4�ɣ���-��OY���$�kG��X���Eq�3�~A�ڋ��:0��L\��[g���ā)�R2���Y|N��`T���w7=�p�Z���X)��,pP��&_G0O��bR�z��Ɗ>� S�i��p9��=+�΢�.%�G���Q�@��27{���=��Y�h�J��^vs��}z���F����yO�@�թ�`����|o�8�tW���~�G���_�X�	�vy��{Pݦ��]���\�}Yi�]�o��t���N��'�����r�c���C ژ�*W͂�^��aN����!(��-��Tb�'��*��˸@�(t��#Tg��� �I��uB�(�� ������֛�B"�|���S����NJL�
QXH���{�����Rɾg�9��a�[���%����l��e���^m_� ��W߲��m_��H��E8�5��p6�	$�=h�.�U�D(M�t
��j�&}H>^|$���v�@���Y��p��LY�٢�7����'3{9�S��U��
V�;$���J� zE;�)�o�u�hr�*�+��fH��w`ƈ���ڡͅne�=��R�"�`?ԷP=�=+<�ORT���j�)�y`����3�zH=|s��A$�U���?I2����sD�u�����n�	������<��$�'I������ߙI�䵹���eBf,�򆉹���-n[J��v�0�p6�~;w��v^<�RO��R�9���6c����4@�W�Ұ�P�y����R���mV6�!��no�������oe�BD)"*�&,�I j6�:�,,�����?s5� �3݌�	�F�)D���ɜ�.6ARq�C���`y_Xe�f��f���{>��7�>~ʗS�ra�g�����+������R�a��3[[r��DRi����ӥ��ȴ�9����_C�s2����܈W˴4��F���\�Û�����ӑL:�H���=�?mRI�a���Q�?Z�y}��^R�����K�4�_��̚G�L����s�9�������a�}$�.��4�Oѡ�
�ް�өNi=��d o��AUr�|�Fz꓀����V��t�H�>}I�Wy���?f��G�K+жy��-$t�$�^
i�l�����]vy�;�0���N�])�D C���c��2Bpjf
[���e,c�����Wʧ?�o�7v�/��\n#�(=Hȷ:O��D!?;���*�U<�e�@�C��+��i:|TN��sFl�hh����X����a�w�Ԉ�V�
����c�߆I���k����ӓi �{�z8�&̀��Ʀ�Jh/���j,�&�t8����%;M�D�f3�$T��|@c�qp_�]H���U"�C��`\���`7�̧.�t��F�<\V��K��i�[ë:L�kLeca�%5���1�ZA�2�Pp	o�`�*����a<,��I�M<L���!]�2��pC�3/?�{_��.gV�J��03�a��n-��j����p���G��<�{�>�m�	���͂9]�G���yD|0�`�^Tf�n"AJ��ȓ&�s�v��;���:�_�B'�y�6��V��u�3p�m=�^#L}�D���IZ�(��|�����d�c��"(*"�X��k~���doz��g���~M���%�D�a��fW���]���}�@���ڃ�@�������y��dQ)Q���$o����WZȩ�(��hM��m�^i�d9���J�	�!�"uT^�`��ȳ(�,z܈/e�:q�e�=>e<���~;�����T�\�;(cĄT��CVp���v��@�r�Z����.�LhQ� �7}ȷ��Ɣp+y����9o��)&�+;�7�
�j�੯�q"�?��'�T�p���(��:��]Y�����B�J���t��&F�&D��x���13v��->�����t"g�]݇µ�v,���l�/��ؓ��DM�v�u������1��^�?^���r�Mo�>�}�_�-me�=�Z������C����u3#Ŭ:ǲ�n�3�Fk�\�&T�7��8X�#��D��A�8<v�z�(�>Q���Hg��IwRv�����M�6��$$o���2�n>t��G�g0E^y�i{�1�,܏$NYu�����8H}G8���L��f��2}�t�X8z/|��IϽ�c~��4����?-��O���;.<@b�f�V�B@���p��|^]~��}A���;���R�e�5�Qp��<p�:u��DI⣚}��W[�~��+�Ju������4Y���]`��B�e/��l��'CC�pf&?���6�b%=�+��f��k,^.'t����������7�|N{d�.��M-���<�4��Ut��� �Y8J(�������}|����E�$�&72E����ESg~X��/�9�p�ll7L���S�����\r���#BJ��k ��L��x7����:$�&W�9�Q���iw�f�/�5YT���	C�����-�Z�У챁b,o�������q�*�GZ��s��噍[	^�ʡ�O%�nn�؀�˝F� Ϥu��~ͥ��0(|���J8�ve����s�g���EVú� L8��j!�}�L�f�7��
�:�˘��q�N�:��1�;���Z*M�He#9|�'P�b�i��i����*g8��5 ���y8y�uD��g�;E-�7!��|�d�P���|� A�T[�J����d@���Q��T�e�V�*��g�P�_i�Y&���p��R�k �v����<���%��V���RDf*I�iF�]�Wۧ����m���hG�q#	�s��Ɂ�Cq��$���;�����շݜ.����V�խ�ٹL_�����9�|<G4\�C���;"j��;�p� ##�J`of ����c���3n�z,D�K�֥S������(�����"�B_�BԪ����i>W��ǖ�U�$5|Y#&�a���ݣ9u�\�ɘ��@8�[�~S�}�&b9r=��X�'���`��rt��Ӕ´D���W�s��-���Y�'TP�W�g\탠Fĉ�<ze�s5-�_	�PP {��W������´"�ب���(Լ@R*c@���� �9�Hxp�~�������K�R�����3�<ae��8� my,��7w��tb�>����)���h��R��fC����M�g��>�d/�T1}���C��#α��ZxuG/I;���D��'�Ln,?ވ�RGM�Ҷ�Ν���7W��+������O8�CO���c��7��WE&�Z���h��کBeV�o�����I��\�X��.�w���{���3*2q� KQ���}��'�6�9��bFƥ��k��e5\te��Y*������G;]N�/%5�`��R|���(���"=9�}��kŅ��C@N��A��q�`	��$sRo��m��Dh�1�̙!�:�����k?�K�����1e�`"���)W��o[���]a����Mk!�ִ�cU��f���G�ۙR?o�<R��$yAl�G!���R�9L'��.OD,e�����{�3?Pݻ�
�a���`t:|�s!sF��;����ƔD>�_�$����cQ%T��-e'=���Cj(�(i��6Q�|P18�ʈ��j�b�OCJo�]{��	}�X�T)	�Ov�����YH��f���L����}^��ܧ���\C1I<�5W[ݧ7���@)β3m#l$Q�JZհj��Rn|.�";rj�s��Ac:,�?�（��[�X,�7��������zK<��[U�G�kBN*�bA9g�.OPJ���6V�ש�^�uC8�p���>����u�BJX������A��A�(��f�E�Z9���05w}��̵��N�^�	,HXJ4�v_��%=#��L@��*�'Q�z���D�a=2���>qx�h'Z�R����N�SA� 3�n��-G�@P�����2��ɨw��wP=M����&�� �2�8:���u��D]��G:A\�s�4m&�A�(Go����>����٥I������ԙ{6Ki����^�����\��_҈Dƹ�0s���8��&���(�ic�-�sY�t���覐�+h�C��v�]�F�|���#�,\]|^`kqD�=N�ӆ���f��0<A?:nA�!0���wX����q��LS"�%Ϛ0G>/�Djf��r?W0q�e!EN�{�j��˨]�7{LF�j�!耤���8��[��^����%��4�K���e
0�*#X�]a�*��$�]�놏tNy�ץYD`�?))���}F�M%-z��xp�cbȓ�bA�EI��x4��,�����ǌ4g߉����x��/n�2���-��{&�DYq9gu.��:%�o���,���P�,����X��.'*��Ю$����^B��Xey���fy*�������)�y��l����:����s��I�q����j�Z��!+�*S��{p��@����^�pR�dA�h�'�������1 j/��f_i���ؓơ@� ��P�7��^��(��{c�e�����Gm��LuCт�(�9 \�aV���
>I��}0��Ǉ�5��,Q�tꅸć��2h��ͦ�8i�GT �5!�)��\��I� '�x�ۖ���Eq���&.2����)և�����]k�N���ҕ���㺊���" Y~���//�w���4=4N��柮޵Wx�y�On{Ku!�<Nv��\��w	��յ5�� 6�����}/Θ�d׸���Ŧf�#�0�z��C��T��w�����ߴ�<ڶ��	�7ґ7K�(��Z�\k�qĎ+�+r�.yU�c'4/������׋��
OM�k&%FA����A�����v紊n�Ǜ��aR���wQ'~<�4�Y��U
3z!�.+��\.�%�N�B�l�ƒg����v��1�$6�{\9�fC�+��>�z�ChюRb�֋p��Gt.�Y�b�؊y�B|�:h��a������ԓ�E��5V�3�/��u��'��g2��S<�i�0��NUk	63[<�(��8f���a�����t�ТP���K�\n�6����p��iQ�o��u�h�{<w�5܅ՔW\����Sڭ6���s���ω���S�[럀�X}�mӹ��l���=Qػ���]����|ơK�0P;�L	.�!Q�γ�4�����&l7HMƒF W�:e`\����,�S���I���.���
T�[ ٶ:s��	�ۘo8���
b#3�lxrhl����|rE�jy��r���k �HqXQ�6�` a�%��E�a�������HVB�D8f�v��H�Dץ��Ζ �$�~:U��p(�L{_�䴍�;�(���%q��kE{��_Ah�J :z���r˟=�����(��ni�+��o�r����B�p8L*� �!"2�	�����N2����	H���Z���7�-z �0D-�bx�).&m��[P�{� Hpx����C�t����ю���.7*m�����ݬ�\u6Vl��S܃M���E���\�gǘ�wJ[ag(d��pI_����'9ܐ�I�4��G�ǦD}t�'�.�Fx������z��Qa��1��Av	}	��ĳASz^��Ĺ��������}U*�+�f�}��|�f��؇[�X,bR�]02IL$��v�x����A�]ˣx�ۺ� %����h{DQ�0l,o����K�F�Dc���n��>�uM�g�hL�kL����r��Q�w,?�>/�ć�Z*�_h�=g~�P���)���U�'�E��)��:�� )p �['�Ul'}�|-�&jÍyı��B%hi�u��ˠ�ߠR�6<���*���FY�� #ZD��,�^rU���Ձ}h��F�{��`S�9���ڛ���>D�t���L���__��J�m�π:����j�!�t2?+�Sn�2��ك�!���.�i�:_ŪAq��:=�ؐ�'xl�ӭ��).��C��yx�T��4�U\\G�¢^�z2��U��&sx
7�_9�
h�e��e��C]�li�A�oAK�I�#?ȭ&D�w4;gfIA7��*,?3H��An�H�Ȍ�h���i��0b�6���y�,/�L�3Y݈��[~���t�^�]d�	�j�հ������PM��0.#
�D	/:��Zֈ���)K��aV��-g�,��FP���� �R8�g*,�Ȃ��Hn!����ȣ�
��5��� u��|Y�(�3tS�����2�>��eȔ�y��0�q����6?x��!py��������E2g6�v-z�!`m��j�8��~&�y��n$�F{���qHi��e%Q�W�1�r�����D���ggw�U��n�� �Л�x�aa�e�'d	`/�l
wp[�ѕ9�z��bѶ�ՁI�u��A�ZڄH�_�(�9�s~ 5:_��[F��uj|�uyv#{��R%�j� :~Ý
��~�s�����pư�
��h���݉�-�)Ug���n%�5p���z4�=��pi�YI<؜�^�$
�*����u�Q﹏��.�J��g��{�p���M��fUf���T>�U.lR��e�\R���;���-�`���t@��\{�F�B[2�!	 c�0饭F��dX��6�·U?���o�������7�,>�L#��)ȹ��i��^�qB��������k���{��^­�Fx��X�j������&��o��� �B�k;�����<`&��HC8��h?�h�!1SF��;u|E�L��/�������9��6%ko�W̨ ��\P'���/�w��j%z���?���2G[��������F=�*���D=w-�j-����HӾ ��Y���t@�l����������y�-�T�Je^Y�B+̤Lx��,�����oP��� �&޻�������P`Y�?7���G�r��"	B�0tB ϠUA���Aa��i��7��p�s���>�aC)�̬kb\@/��.R�=��G-CS����m*���Kq���#<���Rէ�a��;��pvù�<a��HS�s�����_��b)��Q��6�8�I�g%�zY�Vr��1�:�������� km,�.��{ԁsmG9��E�Z�3r�	j+���M�+�����1f˨!�ݦ@s�#�\���޶9�D�gh5f�@">�m��$Ss�b9)��!������^����a|&`2��φ[G!�<ʭΎɃ�!)��?W�I�"����ީ��`~,X1?Y9A+v'�D�!��y%��r�D~��ǰ.�1.?<���smz���"?�V��)}k�(;�.��'X��=:$]
bGU�u����뢪Z�ƒE�ID���U��Z���t23��+ ,��r'H�pS���Gk����Ю� ���0��YE��`.3�lC5s���*X+�9��������R�O�"��N�: �qh9�����Һ	�����jX�"�I��L�6=���_����dW����0����3V"9<K���ӟ�E4��嗥B����1�R(��s�9 0�x�K/B�p������yZ�>Q�j��%|�[1��Y�>��0��	o,�H�;{dߤ%y�%�aX�.�V|�&-G��X�������������X�!\��NC�p�,mm[<�5���珜q`yq�+!3��~�9w]�k����@�	��"��wG��ʔŠ��v?���)t|L�j���$���l��ّ��KJ9���W���w/��?�ȡ����N|��F���������%��i�/�
���Ӷ�@a֞j�$j/͎;�:'N���,�/�ִ��χ]����)J-w
������v�9����#��X��r���I�8QuiԆ�X�h~JQ%ē͛.qU#�#2��9>�$�/T؈zM".U^zX�ez�xk����6�R,�!Oiv�il>�������ϫ�/����	^OϼSӓu��Jz��̜�,���d�~��ȋ���;���{^9ɳ�PBM4?;ິt�/����",���C�>/@�춝<8$���)�}[0��"�Dt�P���l� ���RSL��9�"gy�7�<J�(O��GLZ<��s=fA$0o��q�̐����5��^ zљx��߄�5"��U����q)r����F��:���jh&�B,��Z-CI�_ϑ�
�2�5%����v*>_��+�<8 �N�����U�f[s�����ٻ�p��+t8����Qkf]��}��NDc�^�x� F�aI0�Q�1�@��l�|9b�^ݨm~�+�.�L~�5�`�R�.�ҭ�NǃbE���9��&d�2
����as���pФ*��U���(5(VJ�*�XM��{|��\�W���#<G�2�N��?a��x,���i����7�̂�P}`��̠[j]�DQS�M�D4��u�jh%��^֭��7�nM���:Nĩ�姠�i��ε�������b������������B��Z ��w�~��ٵ�mb֬B�gK¼!qk,�E�X�ރ�tF^��΃����Nc���R|�'��1�҆I�ɚ�◍�Q]�縏���$w��m?B�ܠ�	�c��*6ƻм7�_��s���M!�H���U�ϸ6�gƼ욉��t,432i*���B��ݴ�jpQ�]�\yg��o�k��j�,��Pݶ����	�f�_AT���~�oVP��I������:���_ϐ%sqN[t�O���N >Ȝ�8.��o��+w6��]��&���;G\9�N-�.��+U��II��2sB</��1Zn�L��˵I �,5���)���*ھ�`w�"��`[wH9l��Q��\��wex�w8;��G�v�B	�L�Tit�@����I&n/��+��ɟq�KD+AEF�sV�+ײٽ/="�d����/����N�<t�3?.�|�b�3�'�sC��eُf]w���-q�6�U<�i�� wo�ATcݗ�y��$|0RU�$W��553�MRm� ?�"�gG˜<m���Mg���&�y}V�=���+!
��dÜ��V	 ��_"��V�,A���������qR'��S�� h��r�����c�V=�Rmr��S˾AF,L)z��e����TH{��Q��t��g��(�X���`�5����?�H^����L�S7�5:�WNGj8P�r��T7��ϡ�l�r��_m) C�}�b�DTf��#4�m{T����&K$�,��I�����&ÔbL|��'��ɳQL���ŏ��^'�i]�%_��O�'R5Jm�˨��_�.�����_n�1�
�rD0SdMҙ!U0�t���Ň�b.��������;O������%�FCdD��ìm��
�[lf�[�����!������dh���&9<#���S������p�AxP��A��a<�y���e���"Oƥ�mFq�zK�����z�zN��i�dM�{��R��C�>� ��CH�\
Q�X��g�%x/�Wf̹S aL�X�v�Z[�X|��N@Up��!�p��w� h\9�(��p���c���� i�������Z����n��$�HF��1��t�'���փ>_�0���ɏЊFqw!g���*^X}��W�:�ӓ.Ju�V���E}���m����OԴe�zwo{�Bʟ�&���G��Nt����jɝƶb���wF��̗���� ���z�eS/H�6K��Z^���2�S"eZ�+�;uC��r<�:9�o��ʏ2�+��B0f��h��F]�,��H���H\� ��;��ɔ�q1��2x7�ݱ�k� ��[b4{���)�i\��1�Z�Im��k1yNv6�e*Q�A+��(�B��vo ��Qo�۱�����!�[�׏��\�g�wd�?��z�j�׷)ly�$�Hx�^�#|���G�AyT����-;� �'vW�N�J�n2���R�C��J�ZC�����,BrI�D�3�Q�{ �� ��+�L�6Xx?ë�p,��o�c�fy�:#�Guo,&�*�0��v�C��#cK���&mf?g���[>�K9v�Nt5��o����,,^�_�yү�� �4��0V	�����8(T����*���)�Z�\����	��+�.HxE�A���n��36vr�AdcT|�V>F�X^���p�����D�W@1����]t
���!˕FT��_`\n��z���G����\_s�6ʡN��y�[Bh�`^f(�q��6/�dLx�"k����Gw�Aym�c�m�`�����%���hp���X.`R��4]�n VY���ĕ��P���2W���W�j��� ��v��N-�
[ζ/yy���>v����1�n�y��h�_P�D(�5'v��ԖI\����r����x�]�Y�����'v�����W���nt�c��%x��-8���qA���?d3����SQ���	��a�:(m�0ؖ��b7"��30ۡw��=i͞J�ye��|��Z���$GK�2�<�i�����/y�+��-f�4dg��X����9��s�
FA����d���"{��:h��F�� 2���Np��Y~�B?
�kՅې�!/)�[�S8�����z����a�U@p�7Ƭ�`K�M��*��LY�L���f�,�6��v���V�l�;�"�d3�y.����ta�G��67�𖆗�&�h�ʤu�~ɲ�k��V'���軈Hș�q�]��ӐG�0��;ya-Cs�x�'������$���\A�$<�u�|�|��{�d�T�[U�Z��ȹ�x���G֯�G?��R�����Q7��`�ߊ1*t��6���̊�1��6�	*1���\%0��j6�s)X/5���`�qH	�M	, �\�N�ޅM�ڲ���!�',�;n��q�Aw\�����d:�Go�o��2�40��G��	}�m��Dj�
�n`3't'���� �p��� �m��>�\-��d��A
{#�̼
�QY�?A���~��t���!��h��ܥ�?-�!*$_3N�u������p�/�ħ���5�������HC*�j��	��mc���5�pk�q���Hw��:�n@ʬ�D��O���]F���tI�t���)0��M�66���%���׬�:Z$�1�YO�%jK\�mof���Z�
���	K��A��=z��&C�N)쮥����VC|Xj���=��n�t��]�dC�ӫ�&�;�����P}K��;���Gta첤&��Z�֭!��n)l)�I�e�nH
�XV�"����Bܡi�OH�w�ؒP�I�l����a#>v)��(���ߨH����K�l�	)8f�_n�˶Yol�*�#���d�̯9P�s��&,t�BY���\��8jp�_��O���K%G
���Wf���!(C��₰W�х�)���ެ�ֲ��J�8��$3������6��̬P��ЇcU\�b  ��TZ
o�7h��ݎ��J��z����Dgn���dIf�D�<�)\��|�}���L�Ğ�{�	yM�	�g�����C���R,r��S�ۭ��;�t2��1�a���ɧ>�[F�	�(�t�)C��'?�܄����z��0M,���bXU���m�Q�J/o�#E�u\�p��ev1?e�&��-KQG���k��7U�M�[y��ъڔ�N�4�/��SO	+����8���$�U�)K����E�w9x����	�x�Ѥ�+k�ݯ�䥨͙�[d�.%|�7JМB7��l��T����.���ٺM#g�7W���HBFݙ�]Y��J���p�x��7m$��������uZ(am#��a�$~Qn`_\�u�k?�?9���+���;�m~	�x9���Qヌ7��$?^��/E8������3nӬ���{I��TjKxP0�q�a�~�U�@yp��p1��e��Ng,�G߲�Έ���8���q�c��:e�g�}8�j�4	�/�gI��a����9��Pr����[�4m�� ;;�D/�͞�JHm٣�D�"��|X��	�n�L�Q���P��%��(�d�������Z=���
k�.�=�Ο��2�](g�M���Vu�G:7�4�!w���
�u�U믰���a��eE�`+�_X��pv�e�,M�J�����$9���!?�-co�-�}�a����f�}>�l~�r��i���v�~��Ꞓ-�>�0i���\��3�w�쏏P�$8����I�ϐ����vf����&��4]����.9`�ܚ2���U*�-���ue����DA����\��$z�]d+�en˱���crB�z����2��#4��Y<��JB�n���}��h1.`�j_�,i�X�H �̟~g���z��گ�qpJ�^M�{&]�����&�_�Iş�շ�X�f������P=�z�	�p��$�IbC�(?��iG���[g:G.��+\M�"�����P��
zt����tY!��ߒ��q�Bx�T#:z��|�a{�|�H5��$����c�T �$��W'W}�WsA����F�g(n
�A-A�^�t��7��[����I��Y[�i���WU? 8��<zq4��Lp���߬���r�Y���*�8�f���do��C�i&PIJ�H7���oۧ��+�1+���v!��m�")�S����\�^k ���l�^�d��}��{��z���>``����`8�E�xyˈI�h��������b�Xv^�Q#y1z���puG���MR����Z!+~_�'�c�0�����1$.o���A��1��8胸���`��s��,�.�E?A�zdY	���`I���E��W_|t�w�TD���%	y}�=����k���Scj$�2`�����?���Z}�m�u�Ǭ[��՚;�2ї��Jk�����O:ڝ�,�)Dp�";!E�ŭ7��SR���Ҹ>j�˃���~�*���]�?w������i	��i�C�pݾr��񱸝�7�4='g�G��A.��l�n����j�ţ}N���i����e��6�Mԃ���� �����V=Tkޱk���\R)~^��ocH���,�k.hM�`I%����"��>&*�;W��%�=�������L�x8���O�!��Ή�鈡����vW��c��n�	����ѶlW�N�*.9 �}�2K�r�y@�6�8�8ƻ�X�R�h�O1�.%���%���s�s��y��.F�	BMz>=�w��B���Y�'�����Z�z�����z�PynH�<7�P7Ca�y7�F	�^���Kɥ����Q�"�� je1��Q���FZ�!��9�r��i*��g�HU�O���k�O���}�3�3����!0�z{�1��E]�ʉIoUMA4�:���YVW�(�����d�["����{f�B�:L ���u7r��7�e(]ᐽZ���-��ۭ5#��cJC�h?�����	û�>��w��LI��o?�'�LO�:��ct�Տ�{�/��u�=� EL�i�JB���.Bv��j��Xm��i����� ��!*y��JJ1]�b+d b��5y!}�*�M)�P9Id�8:�X�]�Uo��Xcia�V�N]`,B�Hmb���h�e��^T�)rB��O�S�jwCVKq�v���ֻ�������M��'�BTK�_���{������S��M�˺�C����E�_hV�CeY-�"�\�zT4\y�:�����M�f�LUJ����B�����#���ᐍ��h�� �n����"����7�`�7�N�����u�7]~�%P��FT��U9S�Y�?a�j-Ҕ�H�A�4TC�e��	2�>E�.��e�e�L���qUגr�\h�FA�2���k
5��}2��z�I�_�]�X*����0].��z��t��vn�i��3��^x�i�4ka�c�MNv��ġ_jD	|c��ϵ�t8;L�!�8r�;sT�D�1(���^[e} ZA�.�:t��\{���� �����2Q*ER#H��!-b7����B�nU4��v{�	��Z& ݧ���L�V��Y��S�;�.�m�a�;K8�f�Y���Z���+
/�H�v���z�+�d�9�������B[F��䡆QnU^�0��^�oU��8H����r�����ª�~o��9�AN�p�>7�o�[�E�z�I�_߲nU�`���ۃIz?jK�XZ	�<��OP�<���Gw5�UgH��i���y�jH=ҡ��~w�ݚ���Ƚ�Q����*g(��x5L�?ֱ��{\��_X(��j75��d<ׅ��4��:�L1�;ӟdhI5�*��Ȇ�u��תj��"�p����^���!�n�iga"e�W�,Ggw5m՘�7����SeO���S�l�f��~�r��o��Q�9AN�MB���?Pm/�b�+W#	�p�wr��9rU����� ��МT���S�����I�郈�����o�^��s��l%.̠]�X� H��o#�"qA�E	�V��u�1�݂Ҍ��4��}^����|���h�O&�R�^i%?��Q��B2d'�-���o�4lu���`uu�m�^B��;>��2�G�F���]v< "]�F��2X��f��D���ic�WU�����u��uI��PR�4��7��_���t�7��E�*��%��e�h4~�m��y���X%�	�����J�5����i ��?e���ZV�"��OAqΊu|��'��۝��v]��P����>������F-�;�X�#�]�~HǓ$b���_�����u4I�cO65���O�h�W|Y�j�'����fa�����7��e�pc�ӡ��̤�
�.����	�b���Qv�,�9�''��F"��,��*�����<F����b)4p�ѯ����k����`�E_IK0!T��ad>c	�iS���A��|<U�°��!���%N�Dj�V�k�G�C|�ߖ�N�TNrӈܵӀAa��j��4�h��G����̿�%9��<�h���I���~	�PyyI�L$�6{]:R���-�H"N��o~������h �P�ֹ�1��y���~�5��'�\i�7A�h45�TI��#^��O˞Z������\��l��ƅR�B~!՜�71��&�u#$����1	�e22�H]�'��z���W�%;�\H�^�A+�?Z�#,Ts���ܬƳ�K��ܮΰ��5�-,��&(
�<�,�8Y�z��}_�r.� ���v$��&]?��|�1K���I��Ŧ��LΧ]^�(C�#*~���G�ZW5����S��ݸd]�U�R��rǄ���Zp����M�y<�MQ��%�ǽ��Nވ���|���T����D),��/����N�P-��ٹ�;�*�+�$�%�*�߽���w,6R�CC������~������u�u<���.�GČ��v[��6�+=D�ہ4�m6����fY�M7eK��5�Z��o4��w����`m`<8��|�s���_�$��^@�=`&En(��P��&���N�Ir.��rMAS�>��#���u�u���ǧ^=)�?":4��UÂk��zpD�g���:��_��+��{��@�B�f�U��{�#Zb�������n�j���:鏰ER��Vԟ�ݼ�W��Y����
p��4���)Ǿ�(�:p��V���A]��(.�wx#���r_�O��ı�<$U�-�:���a�q���Qx�C��ny5�;�M��j�������})<`�d&���T���͏[�L�ݾm����g&���g��O�������z�JL�[O��K��,�l�嚤��
P���A�(VS�(��ͪ�^�������:� ���j�����T��S����PI w���TG�����i�m˴���� �M4�<&E�~X���Vdt�������ǥ"�NS��wbw�ouQ 
#�?����V�t4]�3���?z>n������+	�O_]HȰ/�\�(2!0�^���bUu<�!�&Kl0~��W+�Po�43GP>��h��v�3ٿF+n3"�ӧ��߅��#m�S/O�4�����g0�nl:����Y��_��M��2g��_�͠�P������-�B�v��/p�}����x�5�2�6�@�Ǔw�s�����������Y�N��·��,'�$�7̖�����5w�GVb����i����_*����m�h�)�J��"�mg$�,��(rپ��dM55<܆��Wy��A�VȬ4E]�K�M�.��aߜ����3�G[�'-{l@���MV��#�t�?���Ҿ�G���>n�+��0)z׌�ܾ_W��Xt� _|h�H��p�	�5�����$N�Y��J��ӿmD˾�{�#�*9��L�U|�w�W|n�[�V>�YJJ���n�%��V�4�
�)h �N�$=1q�MTtp��j*���K��O�X��d�8�ƣ�4r���/��~��Y�Q(�-��*�&M�<ed���	�WB��.��RLn�-:J3��<˂�Wp����sm��%{e0&�@n�!U��fQxp��c�t�]����?P��l��X����~�sݍ�{J�V,�*�M�<������.Z��x�ɉ���*�*� �,�WLd��/�)L��s��_�.�+´;���y&���]:���%~�n��U��|1�[�;��H��X&1"����� njַ�[�_�cd^�
�;��^SM�2 P���Z���}�T�0:j�M հ���E.�'F�.�f[h�����н-!��鑄$��B�i�R��[�V��Gg�_��L����<x���b&):ik-gQV��":4XN����N�j*t��w��8���i���ˑ��^b���43��y��|o;`�#�.�=QL��Oދ�@`\^��ȭ2ү����<,>�Ȣ)
O����RɮǪϦ�M"�K�w���'��C�
 �"ú)�L��ʪ)�=-g�������	�)�T>����rHĚJ��9K�͌��i�4�j:��q�#���=DW�� �N�^-rL�p�@�U����x ��5��$�z+$^Qov�D�6n�`��=��[�/FdS��r8c����"vz����v�,�́PG[��.�ӯœxdeIaK1_!����鿄��n�Ow�<*n�1Cv=�fd47�ɽx��=ܿs/NH�@k��o�u��J�5��' 0����:b�V��6k�0B���	���y�i��
i�t(�����!}�8��p�7�>�cS R��W���j" 0+1h�Sh���
���7����hφ���gY�Q���67��� �ե���P���0���V��J-3n�Q��8:�o��Ma/�����a47x��U)	�g~�^��?4��Z��@�RHM�F��*��R磵	(f�T���v�<�:��������~�����!"FJ��I}�\�x��-4���	�aZ��������I�5�+쀧y���8i�����?�z!0L:?E�����&^� �G���Hu�@
�TV�FcQ_x��a`>q���dxm��O��P�"?ݓ[�L����I�IW��~ȅܾ;��"2S-Ê�����U��1���bh�c?7
�6r:��ω���B)�gC�&ś�9P�%pۃ�-����b�7��z�>)$u���c+�y�[�WM}�-&qC�>��]/6�� \�ܬ~���<:��)v)i9z`��H_T4X,d[5E`��+��QkPs�xb#��jҸ�ɼ9�(�6�����������g�)l��D̰܅[b40ġ�Q$�%����ÏW�Wh�4A$�\|��3�}w���A�Bi�^¤�D����l�VK|��|�`��	��`����Q=��kG�4�v\�#�.:��H�wA?&�;������m|Ft�ǈ�$����z���ϱ�Z�����x��U�zbY�m��k8���?j1��FrP�z�	I&7���x$fGl.<�+����j)/U�G���O��K=������j�y�}R��-�EB�q2�����|N�-[c3�e��F�����ޱH`Ѱ� �m���2��S�.<���)�g��(I!�}�p�d�yx�p���	-L��f�����[D����v�.[��5�{u �9$��]�ɯ>�g�~�8�8!����Qi7-�	�X�o!�ZXb�H��_3����Uq���}������܎�uPk"�v���\~I��ԡ����M��'�r���;0��dg��>��v0�GS��8h�-�h1$U���. \�������Tݰ�<��v�{�h���fM6��0*u���l�X��!qy���Sf�5�d�o�UZ���,e�8�W�]6�b�����3�ʙ�a�PN}�/�Tb�3��9��,��ү�4?��ԡ���M�Zp��]�+m��Q�7�ۄȄ>-&9`>�D�I���@��#���V�Ċ�&k"��7X/�7�k�Cr~�)��k�Y!�O�@s���O))㷞����5>�k�[0$�M_oڪ�z�)���rNBG�S<mɈ�/|���GYE�\	�C|�9}�}�PP��o�L�9��#���}�v]T]d۵@Ap�0\2�g���Y�n.���z�sj۷��Xw��3O0�)���;>���YX�ɸ�Q���$;�{1��v8d��Z��x���Xؽ[Y%�A��V�-�����f�=*!AN���<}n��Hݷ��S;�DZ�	�\�$��T�"��R=��&<���"�C>c���mI����^"k�7�io��єVv3�ɨ$7���i׼?Ѥ���%7���`3�(��(�Q؅.��0�T���B�b��)i��Q:lc��&���<�6m
*�GZ[g.RB��Z쎠O����{�U�Q3� �{�����j���M��aS����l��d��uge��Þ�4�Q��D����o������Yp�%�pulε��2�xſܓ*.���z�IX\���@e*\�*�m090Ɉ�q"2�r}*�=\�X�-&�Y=�c��!|�w-ݮ�i����z$?�$)Y��)Q>f�	�:=��y�֗�Pny�f�@$��
�@H������/D(֎���Y�'�D2p�a�'(*������+�����q�O����i�q���:5|����B�B�zLß� 	4Ne�>Ӭ�Ϛ��Bk�d���;uF$[��e��z�W0��0��� ����͟��;d�%k_G
B�g:��o�59�j�\��hs���=;
�����|�����vE�Fŗ�b(T�(��ʼ#|���Yaqܼ� �媇`���2^����ɶI5AW�{��>L:�F�@��[�����,�`���W�p��i���~��d��!�c��jL�@��$|��\��l�R�W�y�S�&��X\�foR�d֋ƺVyh}a��Gxԉ�犇|OL*��[�S��.W����l��ep]o�����a	�A���T������?�WFFo�ͪ�?I���z�.b���*fu��JZ��7Ŗ9vr#��D���v������a`�A�Ro��Ӏ`�/C�������(����8�
������8
�c�Ӌ��n��W�{�����^S-E��ˎJ}�߹oH_?}���H�5j�jH���b��9hKq��ҏ�i�¡}R�`dV�M+���'޻`?�Z�?��B�k ����sx#��oH�0D��������hg����{���Yܼ�r�a�4Q��@�Ƚ��"�~�f�'����pwO��az��)����l�[���ioS�h2"��#��ԠI	���P�l�_�ߣ���� �8����.�j@{@�"��m��3�_C�h0a�{܂`^�~��\�Y�� ���X�#	(��>
�[��^x��Q;�8����O3���SɿaL�.B���V���N�`>8��k��5d��('v�G[q6�3^�A7�8���/9B����&�fH�O�{H���	vE]���,
���-�E�6�{��Ez0��J���h��ئh)����Zp|�W6.�4>@P&"YP�t㱆��ȋ��в����c�c�������R;��ӆ�Xvhu�yϺ��y�����Ɔ�S�aY�� $��B�@�֡��W�DT:�*#���C:����dA�ꇍJ}���Ebj�׸|T��14�"�`w��>ĝȔJfw�z�S�l��es��
i��P�"�rc)M�D�lY��&��R�W�x�$�~m%�J=&�vJ�	�q�������ݻ�
Offh1Q����;7w�;F�6%���M�C�.H��Ӌ��F���ӈ堏�5�������/�o�uۭ�*�(�#9Q�P�kK����h���"q���(�w����ř����ۻd��x��?��ȕu!�'Bf|N�4�c�n�� xe���۽Sg�q��~��2��|���x)�y���,���3F >�0��j�N((�,1�F��3Z�h��P�:t@�h@,V�E+If�OzQ/����@��h�H|����˿�'5䊫�W�ϫ .�k�A<�ځ���2���/3��9��|YH��"eE�p���pȡ����Yʘ9����>�\�Bݳ,�q��EǍ#N�ڪ�g0���94���.�3�X(ѽS��1���ߝwMB8|��R{9�ۤI�������Pp;�kC�'�Z�j[mUhA���4��]�]<v�A�薿x[U�	aZ��C Y�ؑq?h�˭�E�Q��C��-�I;�R�U�]�&٣��Zs�K��u�Z�]���w�
,q$�� F�[����!0N�u�Ƞ6~����a��)1��d�0��y�
ճvC�X��v�Y�"�J(�4A�'Σe莠07ۑq���q��wȃ�cþ֍5�f��4����,Ǡy�B�3�H��X��eA}$���:��z.*3.?���;�d7��^{���m�Z��o��#�N������b  �-���}ž�j/��?}�b��k�h�j�d�T���F�Ɖ�vH��b�v4��v�et��2�M\Gy�2A#������<xn�q�F�E�Mzm�U��k>I�	��#UJ]L����p&�~&�z��IFF\i9�gv/��z^Q����q����K$>��Ј:'*���ŧ�&s�)�����dz��otk��Rg'��'_��Eƅ+z���V�lN��a��b��>48㔔M��45�3oi{P��.��̨�J����V�\0��UD�%��jƚ)f/��'m*PsQ8�i��$��V&4��/%D��l{�M�4G�.T�Q4�v��	�rk-�S:�¥��a��������\�sx�Lȋ��	��%�zdOS����Sl��y�f�O=yk����im{?%��aɔ���;F>�d��n��:��xoKĺ44߫��иl�k�����{�7]�{��T(���?�E8�BX��|��N��P�gA��ѻ6�����#��L�8��h��׼T�H����
+dN�C�x��"#6���X���l��_��x�u��u.mm���LqP�� ���/J�����KM.O��]>��D������ �o* Ҳ����L}Z�|�k�)�ѡ/���?��?r���U��<��(6�+g,����u�	�J��¼������#��Nox�E��!a���,&��4���bܟ��M��y�ҊO.�P��톚��POx2qc��*�5ȴ��he�S7�QOyP�(�
_!\���}7٣#���Z�� [�!�>e�$�\ou`�*狖�(�o�"���.v�|�u�/����N�Ҏg�����0Y[��|����>�'�:3x�RZx�F�^B�灮��k�$�4�c���e)�5ۖB�9P�j������:��^Q��#���K<`���*��Y�b����dj��l���U�㛎�c��C���o�*�U�.�o�"�_YZd�.�DR[ �Rr�k��%A_����@���1����������}�g�~&O�C��fq���@�՗����� �[&������ ���YKm3E5��:�Pc�ȐM�!%Rm������K~D�-�2i���'���Nj�������G��N_���r��Y3�5�u��}N�K��=~X��r5�d�y���o�#��2L�T�,�2yʬ�0Z�´3��i�K:
��A�	Ϗ2��s�8j�Mv��-��-�mq:��M�|�us��HѬ F1ժ��&��~#9��{���87�G�	��Ԛ�W98��4e��ߴ��馊��ʷ�?���97d�p�6pHf�`�>�lV:k�v�Q�P1S��?��R��X6Ȝ.��0���8Ԋ�=��'`x�� �=�@��$-�5rS�ɐ�D��z����1G���"�%92���� ,~�D�h6��G9E�h �p�)"x���x����r�x<t�N���p)��?���]�K��5;�7"��G>r����ۼCE+ݷj�7|D\@��_Z����+:NP�s�,Q�?h�^��`�o��δ��2�L#�ur���>��b��l�꠼�L�2D��_:rF�6ˡ����;�9<w;w_��2��o�-[#Y�e�>�nt�7}}Q��dĳ^f"Dr2�S��F��i^���ɨ�~�Tn�DG8� �1��1�s�^�,ԐF�؅�Y:�0٨r���MunD�k:Ɂ�c���\W����72����H�%	��iX�ә�(w�fe�]���l&?}&�,У*3���%2@PպJt#�|6;�e�����╕Ȱ-6�fr®ؿcV+�����A��n�4d^��2;�+�ӝ��
�Ȃ�o*�_��K���}�ֲn�K�>Y�;-����Ѥe��c��fF}�._>�^#8^���3��p=�m�������\��y<���*-`�Y�a%�	u�NM�V���G��2��]�����;�{p����q����+��K����)�d��c�|��=P��ԭ���<�N������!�j�[��F�Ic�X\Y�h��������oU8꜖a��*����G F<��t���>��5�+=���V�;w�v��G_�(���^�yG�����q��t�{h�l��,��]�b� eh*�h]*�`���5"1�DI���/u�D�K!Q��r�N��o���p����Z� j�!�e!�ޣD[|�r)3a�����rk�i_��������dA�c�!�B�W��e o� y)��`��xݟ.�;4���H��_����"��bvp��PL�����(jy�dο���=i~Oh�[R�x������V�}q�1���q�e������Π�Z#�ꦯ��."�����|���&ZA�bPƇ� t�� ��*l�
-����5����.��99�j�?�݂��kցm�41Z��z�X��6� �`$*�u���j�a�%�W(�L���p�Ɏ�n�l��9u:�K��I��:��Ugn��`�0�'��5�[-�D��S��l.�AY<��- Uh���gZX��{�b���!��o5]�h�W�s���Tl������b&�N;�`Xˎ����l��*$~���/8[��Έ���� �N>���W�E�@�ӭ��c���VJIC�n��ˇ�SJ�
}�J?(I�^S��*�E����;,��$�G�������p�.���Z�� ��9�b�8U�5�~+�0(x��L3R�2x2F��|Ŋ������=���D�Pۈn��h�p�$�Bt��Mi�(�-_o��H�]z��o�mjQ^%�p����h�� ��5����;��c�QX�(��S,�L�C} U�E����%���q��=�a�`b!B�]��r�H����-��Y�3��T��^��	��^Y�fK����g]!){��-^{����!;��&Z`V��N�V��9�@�I����r��Ͷ�XgNS�����r����=�Y5�>n�q1#�/ZTj~������|*0���!�g�Z02�uD[5*U���t )_ J����i�7G1̝��l�!.�nX~WG ��ԛ+��ǹy�6�1�LS���.^/�˽��we�&�ƪ�T�P�b/��j3TGp����]� �W��03��7A��	�st����c3ʗ��Y���;&����s$�_o;�PcM褂i:�:i�j�� ��j�	]
ح�9��8ϼf�/4���Y���7F�&�,"'߱�0g�:��c��S�"<m�����T�7�Ʉ��5<oa��}��sґT3��C��H��$��,Y$��O�E�ݶ��t܏�<O��'p�D�����m�|��P�y����ը�Al���We\�&%l��� ���[B%���3g�x���W��,uj)���)1 ������_!�B��s�k�xȡu�(X��(�EE�AM0�^:�����)���<�C�O���8��m>�����UzY�	h�`��~Y�LZ\A:�����'d��n�C�/B�i4�o��a�hݝ�� �լ��Fu���;ܦ�V�(�l�gP|H"��=���W����%v���w�оgw�n��t��mZ�O��Å�ȫ�@�R�c�45�ng�*8�ǚ��p)A�04}��tf��c��ӕ���]�	ɳ5K�ѡܸ�E�=��4"�L}�����nO��_yG	��1�t^?F*_E{�]��y|�^e��n|�H�@n8�MLi<s�4X�(�G'h=ڏ�a��Ԟj��'����`Ȳ��q�%`��\ݹ����8��&�DB6�/�	ss���x��v$)������%F%��@V�u�J$�u�[ ��E0����A2������]�\�s��\��Zb[+��:�U12&��,�A���%�̏�T|-�� w�Ɯ4�E�P%Y�x�Dl!�Ph�k�U� <��cM�O�='`>}� �]���0Aze�����y1~߳P�F�X��E�`���Lzx���zZπ`M��kH���[�+�C����V����n,9��sx���r*U�k��
����-��z19b�4�����&�Ǌ���܁�iR!&�? "�&F]��<���W�zz탳=����K�E.�6g��I��&3��̠�A�,/ϡk�����8���Z$�G���2��u���T`�E��V+���s�ðK��*���p�0���4��d��\�S�VǦ�b�ʧ�6�H���0��b��g��Q↥O�TD`g���[�IuyTlh�{�{H��0q�Yoq��&�I��c�;o�e]ץ見uxP�.��>�\Y5�(��!w٫	��ufG�(�����>���W윾:>*t�[;�Y������@�	���{��i��0�q,%X�{,ǡ$PV߿
R�'.��Ś��Q�Ͻ6��<��P�
8 T�u3�u�����^� W^��.�������Nc"����%4[����=T��\��L���=�	6_R11�7�"ӵq�U))���;a�e+Q����]�`5 ���Nh��y0��̘؋����ٹ5Ѫ�
8�e���!T����
=��Կ3x�~�P4'���Vib�]i�m�1�����a��w�z!��Z_�������H�����?M,��oe�힙X~2��Ϧ��-�ҨO�����������Ĩ_��F��ʸ����Jᥒ�G���i�p�=������SFBI� S���b���.�1_��c�$Φo�`}0k�6D��o�Ic��Ƣ���^ߒS�&F}�g5~���K���*�0�$��dʧޛ�A�VQ06���;}F�N�TL_�����ˀSq(4�<�����)$�[�IrPay��j�E����-9���	����WRgo�'P���r*��
�
<PTѦl�ef�(⭤���jͣ�Ju1�O��SіN�ߜRB�����Ss�x4�#����\�~����ǒ
F���p+����g�J�OE+�=�#��'�p�(N
�[I Kӓ.a�hG6���3�$�i�0�G|�Ui�9W*�xV��)x�����H���{��k 	o!�kã����[��7��-$6FD�V�5�T�y��nʦH�rؽ�7)h�?:�2�Ȓ#�p�u����n塲p�j%	3�ˏ�i��(Y�p���wBESc��;� B~!�+���_Z�x|r<ӽ
� ��L!�&�m��h�(����ÿ:b� ��u0#�p˪���?@zJ>����(όF.�ą�\�����Q����r�����y�%|�A���w�{�&kV���*q�UB�u�������P�}DCtgn�4�?�jծ�w��.��2oE��W�0³���$t�,v�;ʬ��U86^6�^]�$���Cm���K�H-�I	%%���&��{ ��7"
�'M��?d�|��7&�?�0Yၧ��%����1y՚���"6���������Iֵ���Br�|I3̪�D��Z��e`k��8k�\���cp(&0%�\�P�X���Zí��8����!���Fj����>�
��(����
�A����曟��*���x�@+��׫�ģ+�<DB*g���K�A��}z��Z�3�TU���8.�z��@猙3b��k�~�(k���Ч��$�ӥ�򉴰����ʮ�R�ɐ.'�0(���p�$�'����3�t.�fڳ�\:7E x����&#j,��q<����m�	�X˼��_ou3�r6�9!�o�Si!˨V��N̻�'��<��ִ:�I=�m��C- \�n���h����܋�Et�G�]��ɮ��
�{�X;_�)8�Fp�E��O.K1Y���}�t"G��$a9�{�1�c�^��i��م�4ZE3�pt��'�<��-ƻ9N\��6��ދ�$��%U�KnA��$S<�&�m[Fm���~�M?K.��U�`|�����~p^�`y�5�h&�9|�w��������f=�e����z��z�X�R<��;��%A}��瀬���������j�ja(�m��,���^M�$"�$#ZFm��l��
e"˿�f��%��ݗ#bg�(���x0��g�h�>&D�pz&�Yhb�:�
/��y��uf��O�#*��R}�W��*2�	��qЁ�����| ok	hLs��R�����^��^�k5;��h��N�Š�4p�Wϖ��b{!�C��?��_z{ċ�~�W��}J�����J	�����:��>t�u��-�@r���i�~G�ڽ��\���8���!C�>� �;�S���sjM�uj�}�5i�p��ut`�;�ӥiN�	�=���{�������|�s]���>4���R�7}'�0��J���[�E�Ke�!7q�P�;�fD�?X�k{b�f��hl@{� {�F̒T/B�P7�!��	^n���LZ��_F�%���[��*�����*7��ca1!��&<<�誎Eڦ�j��a%8!-����y������ݲ"P�����ٖb���%a�:�n��rΖ��P�x{���&l52��0;$x�GY2����q��;�|/#;c�5O��͟�:����I���\�L{Wd��58*�5���~ՄۋPk��/$3={��9��t��D�y!��]�iZs��l%Zo�H~U�f�*�!�BL�J. Mǥ���y_B���3o�Y)MEM^����_�\�1n�W���&�k��Ls���cKx!�:6c�_�� �Ip�`L�}C���`萧VQ��%�XUά���l��қd��ȼol�i���ˢ�T\>���)1�-�����nJq
P��#�s]��Bo;�;��Oq`@z�'P�~�>7�V�w�<�7�"���g6�8�CA�H����3�jl_a��&L�i'���Df��0��cU�}�`���UydQ�P4�9�ҎD�Ŗ��)!7<Ɨv�{�p����f�tƪH�J3wf�%�Ԧ �_��-@��5���}�L@�'.#��sˠ��T��&g���2�k:$2��D�E��3И��cH>�ḵXF�bj] �7��R!�����ާ�n��;Ǔ�<���{3(���Y�d���� kď1���>n-�,�����Q�m��.�&��v��c$n �V^�\ȇ���5��ɠ�,����	�#e�A��ݗ�"^[Hh���(#Ƶ�2�+i�G�N�>� Q��B�+èV�DjUqW���蟽���%8�ӧ��/��<7e8��P�s=;[�#7jGӟk�7b��I�Ç�TV�$�D����������^������S�4��*!�4��|* ���c�[jkW;���v°����/�=�ع?����������c�x�k�R&������$r����@�� ۝�k���X����}�Q#9?t�F�V)n��ó��\#���� H#��,�G�Vå{��ݔDk�>�&�*";�yi���^	�~��˰b Q�;�H��zFމ GdHԭ���C��k�a��D� ����f2�Sk�>Hj`W�_����S �N��32����{0��eº���{�o;v�HYڶ�7,T"]<N+�'z�A�O��c�O��;Jp���\��ød�>N���;7p��i�*
�S�	���p��qbQm��GO&���q��+ZE�r�Ŝ%��u1�HFW��s�ߘ&��߳�ߎ$.h��O��ɟ$5�h�}<Gƽejkv� UW$���j��R� . Z�r�K5��l˺�z,S��?!������T0�V/):j��bB����~Ot�G�����⏶�R��}�2�����u!.d�ec���ǉ�~�(�L
�i��؛ph�\Ň�ϼXB�1�E��!��)�ʲh���$0X�8�n�g�l���L����S�A*������휧�Y����m7x��8t��x�;�40�rm{�g�k>v:��%�]=&h?{�~g9����k�s{�a5��:������l���氞̔��\�	
'> �nI�(1���k#��(D�3����6���=��qU��D��Ĳ-�y�A�9�����˩���<��G�ٞ֟��;Rfc���;UR��R�J1D�T��뙝��������A�|��d�-�3��~fz@��p��S��_.���f�K�����LM�)e���ˣLٝG#7��L��gY2J���R��7x�}��0\}a���'�����`x���5����U�FnnB��QLa0O��*,x�.#��{��@ty���:$C�}���
Y�ۡ��6j�W�Y����,�R��v��Bύَ�,�2�8~� ���L��\�*
��!w���QKS+�z�P�πjZ/Xt��V�4��N�`�y� 4u�������UNhv֥Ka�TY0�׎E�A�|��q�Tn+j|�R\mrK����FrG�F�4�vE� �Q�CY���d>J����mw�̙Q݃�t�#�$�]��>��ô��	r�4�[g���rl��!	�{(�����On/�KR�regV�VLT�XOkd�ٓ��(���4�E�q��b�m�SV<Z�FlcH�0xAS�����FP���|���sS�$��e���'��Tmk�R	�^x0����V-��*�lI�����999K�����Z�D�+�
o	��Uk����؊V鯂�R2s�X�C�KI����R��BвnH��7�ݔ�X��������Y�K���t�u�K�ʅ�]H73O.exhx.�ǿ�).�V��y��iL�x=6�Z	:	�߈�τ3�L ��t�[����1�=�dK��0��4������+ֳYZ�	��볏J��yt�uوp��=�@w%������&K;�]�c��90�����R<�����B��ؿ�H|F#q� ��X^h���h�J'�7ۥ�Y������ų�y��6X�x-����npr�����V�����u��_8���Ϊ1�O�<�N� �N��?c`I
\��
nM��*�LC���<,�ҷ���|�*���a�!���;f��Z�p
�~�6N��;۵/�zڃ���s��:\��C'�{w�55�ǯ�nWM�#�a 8����#��<�<�����-\�=�$�;������]0�a�Q�K�������p��'�����I��8}�m6�Y7f��a�m� y{ㅪ��&\'A�ɸ��.�J�/��q�aB�q���*u!@V�a&�xeڞ���[���6��j�vޢi���V�@�PNr��v�D/�?Y�˘���CZM��7�{�b�M<[�j�8zw?�^G9���U�[2�x�7o�hNq�b��i���&�����`��g�P��R� �x���M� X�T��bf�<�!�v���\�y(M��un�d0��T#B�����F��Y+dϥ3�@H�:Ѓ|���yW~l8���cg_b��B�m�B�$�w����O�Fu"P�5��{u�Yy���H��$��5(���edZ�,�S՝&��]Jf�VČ/ؕ`��N&��?�@�"_<�S �B�Ч�� -�����X�n[ J��}��?�`R��1�~Eqbvy�<��d�/��/A��Uk������3Y�S�Eܔ��J擫��p�e4��#�>�L��:����m��$uL��9�7E�43� N>1�*�#��=���V�IC������QD��-b͡�e�{�(�D�=ή�x��°z�?�!~О#dRWşu�Z؎��u�eD�}S�]��l��P�6��@ ��i�$��Gr*�Q�O���e��5�d���D���׻1<yp����L���f�5 G��V�Rb?P��Q$�/����R��&Ƿ۴Lk�A�����A�S��)��^[rD�9&�2g������K,ج�S7����z3y��������k����Am͓��8Y"�Q��۔0��`�x�O�F]��˳Q�0���T�����w�Y'`�Ո"�"�Q)�i�U���O�1�@�����duRzOGd;��g��D}�5u��#��~��r�'$�w:>��M"��b"�K��[l��N">+[N�j}Zϝ�9�Jx�K�{�8��pTg6�X�ϱ�L�;ɇM��J����+�����i�.�`n��Y�Y�ߐ�U��\f�qJYʅF�rS���,�ZzH 6���[��qE�\�t�Mr����V$+`�*�0���m�y�V�ǅ �@�����|��q�m���+L"\K�52��UƉ_�_a���E�㩨heX�*�+a�w*�M���	97���.n^q��"z p	[�m0]�G5�d���: W��J�,����d��}��槻o4�����1���Fâ���Wg��@oO�����?�E)y�c_�'���P�
)��I��lU>պ;8N�^V:���:4�/"����)U�B�t"�vwRwrƤP��y\�������%A;YYj8�W%�rE����G�n�.�/�l�C�b�w���Q�GGl�U���U	Oi�~uN����/�����r�s���F��#q�s�P��!��3����8��IB��,e�!��
{�\~%���.�׸�v�&"=�cUM��:<`�k�D,�4�/��O,qs$x���^�:c�����!�e�H9=Pַx8��R�Bւ�J��*�,��q�gw0��g2k>�2����U���z���k̹*��WZ\g���
�܏P�k�x}�*�~�`�S�/��|��xTC߳3�&���o���iC�#.&q�%Jz�Xyi�d��n�L�,��J՘�m����0\�2��AL���ݶ,��ѱ ���s��z̗�4	�� �r�vțb���{� �Mꙴ�R���p�nR�6��;��O�����ś&�lW��-T��9	_(W�;�*!�&-�j̛��g�M��~��=ו�Qs�(D�G4B��/�y�[�׉�?�1�&`Y}_����%���ie��P�����h�)�xHm�k۾�z��`QӚ����Nd������h��e�5�yY�sͻ��11�s�� �%��Q�����N�>²I�p�k=G�_��p0Y�w��Hb�to+$��lD~[2t�����+/^�s�m�fQ�?El���a� �\0�{!Ё;�F���ﰇͅ�OYUݢ�:�����/5��oK�m?ޙR��פ��P�adm��X�[ wm�^N҉��Vs���j����<�=jS{K�6b��m��;��*� c_���^�? v�9�%!7�6-]f�+b���_i>���ё��$'*q"Z�8k�Vc��S	�p�htZ��٠9{a���e*q�5��2�FL���q����A�΀EE˒G�}�8®�o���;���H�gُ��98�-%�͓0�z���N�c�z��ڔ��Zz͗bi���C�@�˛`���-07ۛ6[���qt��Ș�^���]_⮜
��מCp8�P &�:�uH�f�'���'��~�0���ln���;�=jH!����� SLd"�Kp'&���K�L��~���!O�ذ��ʘL�[�!zNt�+R�%��S��1a�R�޶�|�����If��W©<��B�#���$��]��?@��cc,t�2�a��s�����`K�_`QQqfQ�}e]'߀�"9�wX�&u3�-�K&j$ASgZ蟺�O����p4��,�z�\l�L��0�%1�7��u����~K��o���,��Dj��<���y$�Z]���y�J�|.mt7�~A����6+h�7��mĚ�)4���M�-�j���+�0��I�'4��%�@�YW�U���eι�P�����s˸�U
��oo��iꌑ�"#̸*&%��r�fԩ1/�S�y��=�Q��}s@��[��Q�e�q���X�p6�qwa�r��O�}��vg�y��<UJ>A�EJ���ݹ���-�a-��d��}�����r�#{E�{�<���x6�S��{�=�����?\�~�4S\α QrDR":45Ľ�u��;�����p��@��):�wg�c��_�s[w�5%��Ë��	���S$�w�����^9t9t��)�E����i$�sQ�1Y�Ouf���O��=�y��rC��?���웑B��p,��ѷ֐�Q�5��p$����Ȣ$���X����^��a�u鹦�R���>{�g�T����L_��:A��*JS�Z1�+��p<��=�%N�-�QZ+��vJ}�/Yw��IL��5�N��܉����W9��c@Ѓ':�+G�"y��i�sz�,h��].�k��鳷�x�Ǎ������ޚ������G��0xN�<��!��N������I�1�hD\���0��W�}��8��Lyޮ�n�j�-'SX����r@��I�w�C���T��'�l�p$����,s�����D�~m���6�Ӂ�Q��A���T�(,ªg.A��oъ���g��聾�ؕ�e����L� q����0�c4q*�5��4������@ݎt`}h��o�G�Xt*Ix_�ك��S#=�X6��eg����*RJ3�>!��k����i��#4FE��.}�簤����?�Ρ.?q���ہ�����|��H-��n��Q�+�TH��i}�u@��r�D�����k�]�8ä�=9}D���8w�a-�l�4� �0�Ԇf�������S��%}J���i��>�y0��6�"ci;{7�Ɵ�a���n�I,�d@ǤȦM_��jtqݦ9�E�[� 3�?���:�I�\H�]uxh���i#�t��
�`��Jb�T��P�R�b���ף�qY�K�%�!XM.?Io4�d��'�"�Z�N�J���K���/QM|�E�c��F��x
��3���ћ≟�}�j<T�ߠ%�?��ؖS�X����F�zy�������Ҭ2���s�++��񿛇.eGN��lt؆^xd��C1��2/��i}�ߧ6�+�����1��PA�2���I'�g ��IE���Y2�z�����#i[�uֻ�,�ʪ�M�g �<-��x���懣��|I���C��Fl��+7��W;츨zbm�~+���{�KIg}ER]ļ��l�=��G���U�"z�#�����SG��������G�ru�,v���IJ� �+:�� U�c{c�Is��ڹE�W�R	s^x�X���DWQ��ƴ]|��6+>�4[������G��zT����� �ҩ�m�}u�C�q#��8gt�]�;Ft��  m&�̚� �=u�(�l	Fl�,oJ�oy�L�D'����`��q�_����ts�ޫ�crd�ҦQ����h7�w;����!Kk'o��~T������! �Dd�� =����86�(�->e�PnAw�����E��%BK>���F8-&���V�V�����,7&R{l��9��6���-�`"���o
��<��秱���x2�S��Q�v���b�Z�
�+3�<6W,���W3Ja���
S�WݙB�7-�31�q�J]#h}�E��&3SO�mh^�`�_.bV���&ԣ���j�R��8�4��hl�g
���x<�n�H,�Ȟ��꼒�Ӑ�]ʹ�ؙj�P��5��f�z�^4�a/��/��F
�c�T������%����{7���)!T�z�)��� c?߷Qi�I�Y��d�b
��2Ԡc��I`�S�3�/.F��Lt�cA�8�_}��-����P�
2��:�puĊe3r�D# �]�M��g�f�[,"ʈ!��#����*c�i��Q��Pd\%�u�����4���KHZ�IO{��̿i��o���+�X�P:�2"[e�~ͩi���e5�3w�e��f��K�z�"���b�)�w��w�`���{24��,��N�7�!��6�Y���8cӑ�t
���']��rr��G�����K�x:�,����/���s�fVF�+�8������e%ƶ���U�#��|�Tu㘉2!=׈����<��-NOyI�"F=��P�R���>��-d:�&e���!�B�g^5��SG���,n��oЄ����)���EX����ѭ���΂9�p8�)9��3�!�G`��>7Mpd�l��Dd�[x����}0�|������͏��Ů]~��E��"A��$��`y�Hjȇ]�R����%<j_���QFJ����jY�4ZUk��
�f��3M�5� ���DDaG\������ƍ����J@�d+C�#�mپ!��( ���ڢ�fB ʋ K1�ho+�n,��U�Rė]gS��~��M�e�qI���8�#�񿈬���!���U���s��u�Q�ZdL0�8�YJ����E<R��=:�������Q=��A����&�V4�'!5xk��+�r�u�r>fB{n~e�t)�Іݑ�E��S���|5���Sq�#�J+�"HX����N��喰�5Z�7D�V;�}R�^�ұǱ�vV��U�.,?����.�a�ʶ8���V^cde�෬����!�s�����'I�ɟ�wVcy.���Ջ��)�Y`��r'D��æE5�ܛ�W������oWpW��(���Gy�Yi^�e�����:�ز��q9Ԡ�L���ͦ���AM�s�8�z�Y��ϊ�d$��x)A�������./�VŋS��Ό���S���Y��L'h1�ّ�tn0L�1$�E��v<o����=��dk�'���|vw�Ӑ`{E�=+��'�YB�/�N�d˂�N]�����I�\�0p<��P�'P%mn�/��+� '\� o���� �W)���v���%��}���k\�6MZ๔��]����v]r��������8����#��V�6P��Z@XSX�4��[�4�fm���(�K~�)qƨ#�bùǚ)S"���ܴEC�U������u�Ve-�Z9n�h��ⱴh�4�-�^ ɰ�tdh$Z��Dr�݉#26B����$�ȸ��%䙿�]���θ
Ml�傾}�X�ӕ�Fꫂ�s޴BԿ7ݺ'�U�k��ά���(�R�"�I�Ã�BGē�.�ep=���Bz�&<��F���[*3}�M�BW�k5KC�Ν���+$9Y�F �.T���0�B���NAN[�u&  ��AI�`��;���3Z��L�v�Y��5����%6�pC,�͊Â"�:�|�j��C#i����˥�̹�I�q��NO0��3}�]�lT&��n#`��}��f���V�	1l�ii�;�}�BU�Gڏ���uT$��&{��Yc!��v�L��VU\���]�z%�G'F��HI�c��K*��x-��t������V?�36��n3�m�v8G�Q�o�����yhs�Z��F4���\��Sj�+�����0ݽw�̨�v_|4�s�#�ң(��$&�p�k�����1w|���w�ћ�ɧ'k��|\g��^f�.��|у�4��Z⭊���7_����u*���� ��vFI[� �� 偞���m2H�-�^�������h�J}K2�v`�L�k���j3��lCڷ��՚-��+����F�S��R4#+����!s�R���yB���r1���?ۢ1*�tO�f)�X~.�B���HR�J�ӴM�L�����E�w T���e����Ȼ*�9/#�]e��Ut�F��	���qFy�-�>p(��+��fe�䎚���h1���d}0��<ɪO����	պK7&�Hp��8;�V,Moy��3�4�٢�?U��%�0�����x�~V�R`����.0���S�*����(�X�eț9����Zl���~�������j�ѤtnA�-�*P����a�p��Wpk�|��u͖3Gy���aeC�06���E�P��׈�sJ�����I�~~5"�]�_@Ǝ/����_[OW~T�ヘɿ������{ �= om�?�h��L�`~��2sqrU�j����U�P�Ӭ#���w��(Uhǻ���u��7TG��A^�;H�e6���˂vV��/��O��&�m-���5�CMg��@*�|pa�:p�oS|���
ɅW�i�Ü��J�"�U�z�C��%T!�@�����6Ň���3C��9 ��MD�^"W��W�}v�fz�G�㬹O�]-��Ч�nr�����T�yu�n��i$�,i2[L�>$F+�s�s`�و���Ϊ��(�-���b��`�:@������HQ���Kh�՝$�������$��v^��d�.�w�b�?֕��FEg.c�K�]1�aq�c��Gp�낵7g��ߺ��	�a 4�� [av�1*�Su\�7�0���@�}�ї���n��,
5=�0}=�(gV��9ڴ���Ө��5�|�nn@�N8%�F-�!S��%sk_Tşp�2Ȝ��r�޻�?��1��Μ�C�}a�F��B��4p���t Y�d�!�E��6uE����SEc��m�㾑�+�5��f����4�v�o}Y��.߲���!�)��k�0x
i|�y4��[۞�E���nkt	C�O�5��֮FY�xO4o(>�:�I[��QQ���0Ԙ��mxx�P�|�WF�cE�8�]��7�<�7ɵIo���1DPn���H�{���PT:1i@�R3G�G�g����%hn�1/�/rXPK1�
6Y����{�]��&=�����xj��>�^.�v�XZ�>kٔ6C��d  �V�[�gbPyS���;���B�zH���F��j�ɕ�s~��G���>Ml��S�Ⱦ#\+��k/6R<�m<���W��c.�k��������i�.ls+S,1{)AE������1��hׅI���(,K"�:B�4;�n��I'2��T[�]�����o�sޘJ�nc0����`Cp���JdÀ�y�{�5[���ٍ�"-�v���YINt�}��h�KVf�R�����iz��C�r�o�%/��Aᑝ��3bB�꜂K�&�Ŵ�Z�ZK��~l�:5����>P��DDj��[�<r�(�;�Yv3�A�੫a�S�Ò��w�ɟ�����{�a������2�y.�Q����ӡ��{ u�uC���[&K�����)�U���f��b�7����-��ɬZ��L�I��B��<�x2�GJ�e0,����=��)	kb�ǣR�xMeȮ�Mj]�[�i
wi{��3������������	8�:�b�;ty��*�E�ݲiN�6���*��w�6@����t�*Q�ܻO���44t����V.
���#'0��w�t��ʹ@���ޑ�����.�
9�^ڧ��u��r�Є-�GǑ�e��
I8�����wڛ}x$Q�c�fnz�;5�u�K�g_��R��>�&����rhA�J���+� ����x"�dT͟�7��\���ϙs<�B� 	� �̰�$\۫�`��1���q�7�
�Q-������������/�(l��9*���=s�0vw@0
�K@���8����5��V�z������v��*	�3~ZA��/���L����Bk�7���aj��i�O9y�����ڔh�Vȩ��ߩ��=�f7���s[�Ag+�Nc-�v��#D`���[:����gV2>�X��Nv�Ğl�;W��#o�7�٤�n��_�T����B@I�ȸ�ۯ�i�ɩ���\{����G��1C�0#I\��ū<(I��@O��T_�ȧ�j�8�G���
r�̟��>P����+�e(�_b���rcl�����j'��ˑ)q����pc�oNzP�f���.����r�����R���#
��<2K�ߓ��fW�nzq�Z̯�18��!�Z��&���o8�<aB�s䑖��d��	:�������fs�4�(՟('&���$b�ߑj���I5�D�nB̨��Eg���ykF�-��C��Y�j��m�$w� �r.�j��I��E��:��NW`�H�8�м���E�T
�<_��Am���2}�`�{����Bж�Cc}h�U4�- �dV,��kOy\Ԥ3��US������*��Oޮ��IL��>�{�%��	����ܻ��FhSj�]�m�ñ�5Ы��nY�l`2P�X�����hl��Ǘ�@!EcI^���b��!:�m]��L�c�c�m>�o]��`r�yb���p�O����Q՝ǔe�k�lv(�5�ʾp��Q���Y���sv@��};�4��!�x�^���_��]�wE��Opm� �����箅j������CZ�
�#��/��f��an�Z!U%@1�&��a��P�:F�{�y�)�&���Q�Qi{g����)��oG�{��ٚ�5�!3�4�vy ���b�q^?��$���b��STu���dym���,���z3�Aa��l�Ĭj���
b�![#"Ą�����9�� G��g��8�ob�?���x���!�o"�c�'zcF��'��kv��w{�4�E�X-~<4�755�K��_��<&�w3����|-� ��|2z4Ò�q��b���h��wz��N�9;x�KH��*4�:Sr��;V��z3�%��k���A��7�4�43��M���u�PiR+�MV�Pb?r�y�������w���Y*d�i�x�)2v��>�!�{]/��}m�z�/����.l6���9ւ|"��ه8Ҵ��8�(�p�IEƼ��sx��� ��}95"�j��h�AVtSF|)���d�S����[����d�����tsՇ���e	�Wt��w��_��B_�΂�������FX�b��ON�J��c�?��Q��·%^a�KC�(j'�	�=�"���t�Gϳ���	�AE�wz>�~����޵#:�����X�?�qv"����M/k���A����q}����1���FK���!��(�5��j�;�E�_:T�Z��t���������,YK�r/»�2J�	�d�ƭ��1�Q,忷�w嫺��7�,�H:��ҟJ���V��"�R��AҀ��������x\a���;��5��0?��w�EBׇ����]����v����݈�ص����xB���Gh�n�߳����3H�|�ď^'?�2��Ʀ��V���c��O.XW}�Y��M�^j�<0PѼrk�C<]�纛G�܉蘉���� ��,��V��9{ml:Ւ���ΐ�J5 -U���U�/��.��ST�d��V�d>s�Xb��BcDl���X��B0p�/�-�c<��
�G�J_�?�����D2�C����~����T6����n�Ɇ (9�3lp������d\bq|�n�V��hP����訠lH>�c�E먆_��i���iC l�6� ��Z�v�lܑ��&B��K�Ud!mt�S�h�)3HGG�]��?�`a~N�}%��ll`>S{j��;N0�5Z�χ�/D�ZΙ�Q�Tb�_0P�^��4��
���P<T*R���5�Ƅ(f|��My�q�����[��&j_>H�kД��$φk8SL<1���q�rA;"��B��,ݏ2��4׆�灪{X���7;}y��԰��C���77^'�:=[���`籶��4�#��#t���*��at��BI
�q��/�bx���"ge��bC#�`0�Ε�1��	i���%t�QZT��E�����g4lT����V�Rbo$3�W����I#�R��w5�\��Õ}B��ȭq����a�N�������|o��4y��n����%�I��N�Y
���J����W74��~�T����)}1)L
#������r!�o�GS��k)�AM8��
?��1A�$"��u&R>�EM����C�p(�ֈS���t$g��ʍ>|Ӣ����~��/�-J�d��J �"��`Ch�����7��Z�~�%�q쎨��˳~��ܧ�YL�K�_F�}��,�T�v�j�K9^�7�E��,�҈��d���6�&�m'eX���A�_r@Jx��}��(�����tBT��cχ"��9Ԗ�b���ݣ�,.V/!"5�����.���pY�];��S�3j��|�/M�TN�ot�o����6ìd�WG�#}��Q4�"®�I��2�=45PX�_���؆��'�&������%R�^��� LF�㔜�
뾻���غ�3�.ɩ��/����i���t��ޥCcG4g�+���yD<e��'�Vؘ�\��	��!�h�gϽ� �?y��Q���� ���z#����ڵ-��7:�Z�EL�JY�ș.�o	}>�g�p%τ-Uض9�Z�X�����V�E� O/XL�{`2X��G����c�S����e��(�H:ց��-fn	�~d��O�Q���~F�K3!6y�+���u4po��o'�*KhdN՛y��ސe�A]���6]
�L4u�����7��d�{?����bF<e`-w�=K��i�l)aZ���.U����8�0s.��z���.���y���	��%_vfv�dW�����7�	;��R�/ƹ�]p���y�F|�Gǋ<_.b�������K$��r�U�lՏ��?7X�����Ɋ0m�B�	�5�r���)�$Z�i]0=��v�8�L���o�W�mCrތ!���y��A�8�$D�s�6��͊�v��;O�^%�[�Yy��8�1��N5������r��,U��a$O"��*��������`��G����VT�n⠛�vnX�^F�G��̶z1�|�8 AÞ�X��a�e�?�H|���/w��G�y#%�۾dCu7O@�^����Z���$q��G�H���e����1B&b�{M��M�9�{h?k�Ч6�E����)lS�`��x[&(��$�ۋ�<>/�#q���l��������G��Rq�Ɉn)�����#��A��(IE��=`_���!�mnTr����B���� �m����w:?�m���&K�G<(E~���D��U����-_���Z��4��|G�u0q� *t��U�h�����3���y�֝edx3���R!��7�� �3���Rͪ�Ft�-�{��냤��e�ſܤ����;I��3�u ��9���!JC�uNJE@[�{�)���|b%!*��{pYb#���Z7���/OVX:l|�Q�� v�*��-A���wW����9Ierz?j���ڸ)ޟ9on栁w6*4���gO�WM�<��B\�߬� �"I�p�;��F����Ȩt� �lH�:��ݡ��fu��!e�dOl��0g�b6�W��x��g�H���B����C ʠ�V������$��\�u3z�6��l��B\���Z��#7�\X~x�wS�>;�."�Nu.��[�D�Ġ� "�MʅA�7�_x�#Tg���[����]MW*LsE��Â*G��F.�v�}��d��f�)�S�J^�v�f��O�i�uI�e��[��B:1� <��(�����0+=2�,]�֝��I臺�e;4�������ʻR��f�yi�+Z��ee%t�!r��X�c�R����G�kΥ���%�\�h��	�yR."B��^���۶�z{Vv��Ŗ�N��w�N+���`PY�b>�αc�K�m�i�#f[�8V�Þ*PT�����h媤t���X�� �.ˢGGv/�1�.a����s6��el���V�0�J>AAv%�-{�I�8D���a齺A�A���ׅ�]]�?2�g��t��~G�j�ۚ55|�Ù��4.tG�N�#7U���$�L�i|#^0���G'���hO<���B�n�i�.!'�I�}S&@����6r("ڭ��������J+�nCOx�UBJ�R"�J�� -�8�R9�f ��t�ӆ%*�Ra���-��)��rRh�����Lt�s��wp�q�t\� =V��j����@!����q��-�R�`&��g0��g~V���<���U�:��Q���jC^���^�s �\h�[I,�̂UF��p~�}g.��%d���|�x�F��0��6�;.!-�:KߥNWSi��鼊��#- T����!~ͽCc�tr�	��^Ao�\�<,ʲ��ܿ��'Q.vT���� >����4���H�j���R8�=�v C�ɸ0�98���k*�h�O�n�U��M�ڵ�����f	�a�� >6�tڼ��
���EA�G<\{{j��g�
�'��v���r���Y�FyB�&�VTȕT3S�h,�F٧�S���#�}=�
.w����E����������|�r�H&}'%�3�pN�d�'��x4v��W-����A���\R���K֊5�W�p"`־&���g��3 E< 0�b�K��t�Q�F�0RA3���K����6�S��ؠ]�tQ��}מ%��s�B�F�;��#�!���:��T�r�4���cHy�Ȩ�SG�F��H�a��I5?ג�O\���栤��jP������jG
G��y��Y'���:;4�=5ʗڢz�5_R9=���k�ݝw)�R�Ɓ�%ZsiV*W4Z�N�h����"����JE�i����G�=b��yڽ���p-I��u�4�~�X�!]M���(��zWj>C�z�P���WUv|���b�&Q�.۹��3P��
�����͟�!����
����g��SͲM�%�awu/wt�Q>���qI*k�L�7ᰮm$s}���`�|/��`��j�z��C��8��4���WS�����0>>z$VkڹM�������Q�w���|�Ť/0��.��.��p��h��,���&|m��1vJ!��d]���Th�NZ*n�H�/O������X���D��,9��m�eT�����Ԑ��� �my�z5#@?{�`KUcU��fU/�ʓ����D̅ŤdǲS/���ϒ�+(�nu0�M�٨�):ͯ'��+	� �^�i������k�g���P&h���y��0] ��a���C�t�M��\�Ƿ߳�2׽�������2��8X"t������{-�=�5�S�|EӘ�9ɲ�WyY��-�_8�����Hv��Mv��6�V�����W�z��ײ�r��_,XI��Y_�GjGZ�
��Z���>��{�yb�g�Nԁ�]�}�Jj�1�t�s���wC�)�X7�,~����T�QOr���o����B���C��2R��GT��G���_��7�W����^���0���P��� +�ִ��b���L�4@�r���A&��0��b�D�Z����bM3U�"�>"
�H�o�����X5T�����-}	�5,_����$��3��UY Gl%Y���=5Y:>;���_~R�&~}�T�:�K�_�Wkl�F��0�yn�**7t�@�o��*u����h���,tI\b��(���_��t�04
�'w�^�g�����}��#�����Lr+5ę�S��;˸�*х�́\%�։�ns�Y�^|)uF-hwը�/d��oį9��QpE��
��o���#���S�$K��~���|�<G!w�5�Jq
걼����� �����ϋ�s��J_MK胐�U���J�������/�M���:��)G(�������Q�X���w�6i�,!{��0����H��d��w�r�KbX�װ�&'ӳI���u.u]����W]�g,�)2��[�L"ˀ5:8�Pְ�/쉔~�ENx��v���f���8�Chۯa=C�Å�8��_����n�a@)��DM��Y��ļG��:���������C��pQu錎�]�׫Z���|_�[�+�
X�WnG�KF�F����u� 6k`�����fT���m��Ia�B3ͻ12��z:2��M����Ȳl�?�}�m��Y�=�1b���e�(��s�����a:�!�Z0;��,�7x�UV|D�|ش��jV��Dz�Wd?̤��T8�7�?ʶv�h8�F}�UN ���sORh~�@'ء"����2*4E6�����y��34�E$���j�?�� �v`;"[�P��shO_���H��C��9����s�-X���Z��M����D3�RoJ1B���sIP�1����c��,�)�%�Bs�8`�#r;�ݲ�	l3��R,u�H�0!�wpP.�o�pK
q�*��@Q���h�	�� ����ЪeX,�n{���Y-��]6(�䣔M�x��QON�ޏ,�=ZB�+U�(6�̊�2_/k7e���"��j�6�Q�W�-�9q�- ���]�Tn�~�_A�E��mȎ��x�>����:�EFUf ~����>ByU��_�l���+�=��T=r���������:cO�'9��?G=Mŧ��K@���	ͷ�=���#��,����{q`)v�'r5����Y�B��.T|��`)d��ю=�ͰZN.��**��_Y)ө5C��ŏ{(�Y�?�uZTɼ�:d���J�S!�o�`	N�E4]�U}t�515�w9.��Y,��=��Ig�NZd�*S@i�w)�������)�G :a\��)Z�[���n�����H���Lk�o�(f�䋆R/*dQ)�O�ߍ#	�[eF^A���MY� �f�C��؉�����\��Z-�e�\����1�-Hn]��s���_��!Bdv�Vlj~^��Q�)�d��g�D��ޯޗ�Y�7I�7�b�{>���ן���/��y�w� ���94?ٍ�E��U�رi�K��1�ε��ՠ�'2a��=&��Q�cPk*�.�R)��
�3���U�����.Ã�ϹM�u	q"��=��]�z�x&~&6b?��)B��5�-�#�3���TZ���Q��5C��P���2��w�����dN�ZXMBH6�c�Ν�mݠ�� �>ޞ�T!6� �%T}�t��D�F�w3�uo ���C�2r���̅ۯue�� �!,�����*c��t\N�5��hK���ɪ��o���R��c�Q��vd3��S:�v*\/��_��)*��Dg�s���8���͍y�F#K#.-Z�]d�0��݉WCv��8�=0nql)����#��5+`�[cťH�Q�q�L���\1PPi�d6y�邡�e[��xݮrdA��s4�Vhm�^&�D�Rua�>=�Rօ���Pl	�@����@7*Eʟ��"V:�S�A8>9����Y�3d�ۓ��G�V3d&sI��~�
M[���T7��}��m&:�`�.���9֖W7ş��;�?�!Cޘe���yAS�e#�V��Gi���^��\bi��]K�pn��df�i�=��n]x��2"a/A�� �s�4f~��)���Fϗ�Gӯ����?<<�=&6=ԯ��uК]���(��Ǻ�;�|B�}0�/LK4�X��,r��}�����.��N��S�/1�J�?]uoʣ��)o!��~;3�y������lU�8esqX.��;:%L�lZ1���%~��o.|W�*�>r����n7��3d����tB64��	t�c7T̒��aidc/�TF�H�X��f����e��Y��Ю�n�E�����i�^v�)ȁ$�(2�-���?�l����L�.�O�%q���.����,�>�ɷ�_"W�s7�p�M"��e/\И���?1G��4	�1Lb���܌������9	��ٵN
�<)o�8�bŨ�&�E�G�Q�7V�X���7<AVo�ZA��Yžg�h�x�.<��$����F�ћ6������i��>n�>���8�qj�͜�dUEW^M}���m^�C�\�\�i���Ϋ<�2�����O�������s�F��$0dtfؑ�<��ۮ$l,Y�;����"��P����u��G4����Q�Xy�$�L��Y)�����jb@)�~˩����G܅҉�4�.�H�����:�^�|A�9^42QGFm?��� ��ݙ���t����&�R���M,�!:�+��S"q�󑳯>˧��n�r�#��Є��'iԠ^ftT�Z���D��:Q�8�Ȩ��V�*�N���'�pBZ�Ԩ4�oұ�E�e�W-�5h���h6�wT5ӄ�{���S��������:�����S���U�-ɝm	*��Z� ����%�94�"��'o�8�Pp����)��<�����;fV KG'q�@�!	~|N����W��A&��s�.�sz#�#Խ�I���H��5	�kw���,�[��t\ޘ`���i�أ|�Ŭ��,����!>��ܬݛ�
��;�`��_G�	c"H,�+0 �(�mR�s��@�oP���<�Vi�0V�L��_^T�=�[;����6K��������$�Ũ����@4�(��/R{5��n\�8�@�<�V*@;�(%�Eʻ2�X&Ķ��9���`(�s�|"��-(XV#>�)�X&���������׺Ӽ!�(l��\p��ū6h��������j$��R#��N�x��*|: �mȓ�ٌ[~`\�or�ϡT���T�'s��oF�KV�}�L�S��k�}9ܑGQ,���\镡�~b�-6��-�����CV$x/X����ɖ��;@���ѵ���bl5A�|7[9���"B��׺U�M� [���d@�oIs�����nyvo��5�dT�6�/q�NB`����WӶ�LE��b��԰u��e�f^ZQi�T�:Pd���K�ؿ ��,������?�Q�f�TJh��6N��h�&�*(����&��c�B�qĐ�ZM���WQ��f��@O�f;"�}ʣ�h�m��4�mHLp�� b�ͮ�&���vEfU�z�X_a�ޮ�'�i!X��1�������`�6^��LāF�݅��"7�_/�=A�]A�#mLB��J�'e#:%j����Iy���u�d��5�eU&��@27p�
��a�t��&��b���k���8�w�KUQj˙[tH�;�.sFK�� ,4�e1|��3p�W�����~����Pl���
ʫ�A�a�tl��F�(@´M9բlc]������ؽ���i�$58�AT9��yD�O����w��m0���eR��Od��"T2b�����a�!�ʈ����w��k3��V�Q�&
���0���Spvs���{�m�?�S2�<�6'�J����B�sG�\������gbC'B�$*��Y��6g�K/�6�q"���}Sa)X(��<}o�8�gv�tZ�K���zc5&�3h�9e]�2������J��9�jy(i%a�lӃE2c`΀?k����!��q���m�1>T	����g��46���	�6���w6���1�F{��rͅޓD��/��v�E�=kuS���#�EX��4� ������|���O���TZ�b�r�`z<ܖ� �/ېF�n`�:Q�KK8a�T�ˣ�	��k� �,l=���Ö��#�~�E�sO�܈��2��/bw"^��i8b�EJ= O�L3�����_��'C���1��:�c��n0��g� Ԥ���,������,3ձ��~�-	�����[�����u��B���w�R���K$�l��/W�ӈ\�"җI�.
��}76)�.��js����3�,Z��1>�RE�,��꿍$�ZJ�e��x⅔�=psc���\j�'��o�.vT���m�D���9�ړv��^�� 0�9�%-SY8'.�X��9����<�pK��@���~A����<�D�}����},�j�y�i�sUh�����
g���&��|��x�ƾ����}g�a�cD�� �NY"hfnJgH�(�3V�?�F?3�Q_����c����]�u=���>+�N��R��e�ɂ��s�L�#�3Xo��,�B�7S�Hn��oT�&�˲�G+v@�H�&�k<Կ�9��
'�)�lV�b9�B+B]LFX�5�a7��U�ݳ�:ru�\ټf�4�i�|��T�z�ˣ�����{�Or����ڲ�)<�x������;^�!H��.9vA2���n��X�oi�hH��s���sN�u�Z@e���\]��}�Ciƻ�]�I7 ��O2�`9�e�h�߄�^�<K��JS>9D
�t�̺���X�\� P����A�4��.��S��9)�X�1���.�q�A�(����T��ނ�|B�D��%�4E��ɿ8P�R�}0Xd�>o-3�³u��S#o>���2�����|�f���. A5�Z�9�cr|p����:���]��j>���m�r]V���R)'���N3���n���`vGM��Ȑrx{��u9��3UͰk��6����s�M�Pk�G0��H�j�Yr��K����3f�9�f��7���� ��a1�"&������:��	�)�|/���HR��[���ľ+����*��'��\��d��jr�i�X�Al���A�Ia�+��]Sƴ�:t��-zه��E� 
�5��t{}����n��8��/������N���64��S��u��칌C�L{�/��%ԡ !�:����M�Zx}C����-�&0}�pZ���ۯ� i;�g��TO�0�$y�r�^��%-��l����(��AE��hY���"��8����FJ4Ra�|xk\�[�6��4��������g� �4J8���� <�L��a��c�A}hJ�*�$��o�;��:%�s��u6]l��;=���T�C� ���Cc�w������ISV�r�pvH�=��c���c'x��M�����R�P<��~��YS�/��SB��J�k�Ͼ�'��Mhʡ��J�e�q�&\�QE��u�̽����]	��H@�Eҩ�
�t�S�3���Գ;��~��=i]��Z�%�G���8.�f,�o��ڎޏi⺔�#|�M��9�@C��|���h������Ixe!>P�-G�5�bai����o�a冣� ��pu��:���RDw��*�ˡ�>	�4�:n�&�H�H,��xkɼk�m;U�}����?O���lʁ1�8zf�^�_��f�FD
/�qT'�� ��.D��s$�]��._�Q-�Cl-�;~$�������¥6!J���`Ma6��������+C����P���½�a>������^�@d�}0�K&�.�"a���n]�}��U��D�]D��ۮ��?	&;�MTEm��E�4��/�'  T&�2��r^�f���#)VTk���+ʭ�x��x�׉ a��D`R���0�9�,�k�ة��3R��y��=��C���t�Ղ��@Y�<��':�����+��hJF`�B�� )��N�1�w�">e��;��L���b$��ʚ������^���b�3�:�,À@�h-��_^�:v��\YU��~� ��m��2�]��`M��0����Z`ޅ�k2�dZ\������}�	�t\�Z@�=�(7y�~��9��9�~1 8��輸'x��SG��͓��2mt�Q��?���PwnQ��Ooy%$��F֝�c<AFƀ��� Y������;հ����J$�[�n�'��C���D��萌�;Ű�g~'�_�Cmw��l0M����'[b
��b��7.�W��+�T����5s���1+�
��6I�ԍw��Z;k��M��GGÛ���ܪ?�;��)��JneaY�z~��]�lZ��m�ÀN�:�y�䖞+���<-����%����n[֯�a��_	�0�'�8���,�̹�0��*�"��fȍ��P��`F<�O3��1�Q��Q-�UsRaJ��i[r��-e��]|wο�ݎZ�8臑�Q�~�0���Ĵ_�W�o��&�}���
��fr�H�N	�Ҝ@o�|�Bϱ��m<�T���7/�Х�_c��1�Xd��8I-�K�<�۪;6a
 �@T�B-Qȯs^�pon(�_����j�u�Yֲ�J5�Mz��1�X�,�����S���Ț��<���SL���78������d2c���Ϣ��(����O��H��SvWh(�I�=�[�Yffܯu��
�œ�~���C�����_t#�������w�e�6��jJ%1����N�� J��N#��'�ݗ�Lq�LL5j���_pD��J����x�WHI�?��E$2_��e�anȸgR�i�2J������5/�wcr���u�OK���6A;��5�<���o�wy�����Pʾ#�Q�+��BL$����߶#�(N
'���y共a.�@9[��]������8���!����p!��B��@t���dԡ2x���h1)Uڷ=�q�Xo�v{]�!�&V�%;sK��6��%6���~��X��f�?	�CZ�'���(��Iԓ�0^J�(H����� ,��f�7\i�!d׎,Da��V3�c4�8�K(����b�y3�
��N�Fp_�X�«�+���Y�~noŲ�YƤ��)RF���)�#�S��j�!`���\��s7s����r��k���+x�TĎscK�Ӄj�������'�/�>Y���-����T���Y��Ƥ¯��;�1�.6_	 q_���nE|�E��:�?
��͈�->�����,�[^�~�榷�Y���S8�^*7�xd]�: L�?q�UCO�k����u�.DOIA�󕆻6��>�;!aG��ݬ�g���y�22T0("I?RZB�0� 	��/�Ey�}�Ks�th�x�`�8�|D�|sC쀾��rT}�@z����ht"ȣ�?$7�ϥ͓E�; Gx�
�T��ΆX�/����D���K��R�^�t�`��w��A�\.�x��~A�zs�{	��(���h�5ߎ�`I-�&��o\�e�?ua�EsT��K��Cm�6p�V�]㺆�w�QK1cnM�x�o��o��t*�
ijU5�V6M�M�jƤ� $*;2��_���ye�����+,ښ�Р���"�:wM@������v�=|_��+�k<���u�ۅX�e]�s8�焢���oJ� �x#���sp
��^��L�Y�mH����D\3Λ�t�k�����$*Ǧ2Τ,7��'9P]yU�Kc9b����A� �9�3#��������WV��IVz�t|.+lyL��̈���I	)��P"�m�b 2�A�{N���H+��?��������K�RB���!::D��)i��\	�D�J���@�[��sF"��̰�)w�=禳i���5&�_L�,B�7q̷b�BP�	"M�2q÷�Ũ���_,R� ��B6�#=�di����p�`�>Nf�t�\�Dܲ*'�
@*^x���zd�%QZ��T���?Jw�P�P`�+S�yXo�Ye�/h-c`M�"��Q��_|LxrY�(��t���N��D��%�$o�`�f��ĭc1�c?��Ӳ��}��MO/���1�/˪�����^�xV)����bqca0ʓ`�M��1u��_����y8T`{��;�-�� ��«B�ҘE2z!��n�y��_j���']u&��ʨ��ݦ��TZ8�?95�f�z�6"��-��L]V#��f
���@�p�t��B�I��!����Fҧ�T�E>G1���*v���j�R����{�������Y"��`>��������Y�`������	o��f@�
���ٟk
�*sd���,GX�d�8�h�I��#@f\�n=��d�
�i)����?m�=~V9�׽3����a�_����	����=��o_"hWF(�,#���Kni�T��yٵh"g����$YZe�����k�]�L �`:¯�7��b���i:7O��,/T�����r���@8��p�U�Y�~!k���J����-#K	��w�6��@��dtS�Q�H�dX�h����_�42ة�A����pֻ���q���a?��9\����B�/�/��y�/l�BMX��Qp������]�^n4g9�\WR%�)Ze��F?5�k�#7��`+G��H���p!�OE>�]H=��>�7i���65�q)8ǭ9=V"��ؼ�	:M�V����$p_?�t>�݌+�QL���}�#�.9Lg��E�`^��zp�
H�=a}�hŒF�Uo�դi�֋�!���eq���%�U�[��v-�z�)S>A����5 rF��,g�e����7ҬO��$vAj:���)Ց��Ju���>P��:��&b�f� V�LS�A�+�U�00���$��c��F>| F��9o��5��D�Y�Sc�y��U\�tb�^���iz���+��U֨:��C�������w�	� �jM4w��ͿP*�`I��q�#��'���k,��%M�C�7�B�����V�S~لY����Jy/��JD��P}��T$�s�j0F��5!ō��]jB�v�����cptvL@_����'��I}K�����@��l�>˔E�'3k�����޹���o�&c��+�͎��eu�8� ��|IH���z}�~��(��<���H���Ϥ�խ|i:c���TH=yJ�c�U������(�nFsL��6���}���9�gJ�H�?v�cK2�u[�X-�!ff^�[��h���[H��^V�`^��Q�I��G�/���C��]�VW{�ϓ���(B�(��S����,�x�,Z��3����U9�UB�3�e�����<$б1P@m�O�B�S�y�������e���[�V�?�P�$!��V)��$lDS�rY`�QL?�K�3I�>V�q��+����Te���pS;� 1l��tj Z�S�6������B�c2p_����]��Nq�6��!-�u�W���.�T��B��x�R9JC�
�x�z��8$V����YC��`]5�Hb�%��*�ǌ6Lc���e������(d-ڥ޼�$q{�LPxu��IM�po��T��*z׆i��c�:r~sC�"��`�<�T˝ם��lH��]�[=��JQ���QF[[��#���R���=7(ct�.����>�>�Q��S��> ���ʻB�.r �7*ȖP��c��?���>D:;�e���]�;����τڈ y �f�P�����W�&z�MR�C��[��,2�G ��"a��x�����N�0�]���/DnW:b�(�<`T����}���"� ~�6&�0	��;�d��{O֨�a�����@p8 ��|�H���6�`��/�΁���2��6����ِ���$5�`v3E�Czr��:_��y��6���ѡ�������MŐ��߇w	:^�fb�	J���X���)E�Mb�Ij��n�]Ţwﰳ�f2&�6HL�Y(�Q�E�A���"����˘�~��8%4E�8ei$"��5��_!�	�0��b�ϕ�cb��ƛ���E�$t���,'k��*��CL��\5۠�t~[9�Ͼ��dL����O���t�E��v��lP����OM�]��T~2����W6��u4Q��cR�U��9B�i���q�u��)�q����	U{��25��L|�Α�`�ì�ı���f�``^��{9��Ӵ���}����ˍ�W����l$ng���X�,8�16���j�9Sٟ�ʃa�GuĢء�X
e��D4���+F~�W�OǉT� /F�%�|f��X�w&Ŵ��p�}R>��Ô���D�_��v��.I�.N�	�7��׻|Ɣ~t©�6��ҽ�V�{���ߓ��Zx���PDċh��5(�X�d�r��l�@fR����b ��<���OT>K�BT��|:CT��)" ͦ����jRG�j:\5��j�"�㿃o��.��Ud����gvrΡ�NE@��4�o��-���X�3W�\�=(1�:lƻ�͕!e��������;�0�A�6@ΞZ���C��3J0c�[�l�8vOBX0}����ۇQ2<X�) \fCȐigR'�?x�X�������H�9Y�g�L�KSЩ�b�b��rp ����'hߠ�K��P����Q���h�U�w�MCZ��Fvs�\�/���k;�R�Y�$a$�t�;��G�xo��%�K!<Ji�Ly�ME�7��z촥�-c
�=���c�%X`L,��խ���\�ŀ����HBFM�n7��o������֗�sx%݊|Ḽ �� �uE�|��]}�*�i�o�ح�}�zo*�)���.*�3ݳA�1ȔR����(�YNm37K?�@��0�1�z�%���;��=Zo_�U��al^�J.C0�c�GW����U��Bt[{��	�}K�dK�������+;�|��2�	V���w˒e��f�����H���n6�D|�9�]t
֫NX�
�d���-)&�@H�8E�]1D4������1��$��4��N�ػ?E����
=k�6᪳�"�JS��K����@�9RӘ1+/���*&;\Q0�k(Ѳ���G}�+�y^��{j:��<�s~O���W����L�TV=:�� ͖]���.�������$�M!��>r3<QJ6�Nu²	x�gn��z#\8��r����gt� Fbu' _��仒�Z� Ek߄�y(FL9��?w��ܼ0��8��{.1䉔���{ƃ����ؘflõ����W*�;�E@Kƻ�]���=�eR�j�[���5]O�͑H�̤jD:�f 2�-��ũ���&�Aѫ'&������
|2UQhx����K��㰩<]!h�plV���$�dm#� h�%V
��p}��"?u;�cs�wA���A�'��p!�=�!6���e(l�"ϵ?��{��Nϙ9
�Q26��(:2)�@��� �ɖf�����U���t��z��zUB�[�ȹ��Sj�Iv�Bw���s����v�VR��ׄ�lT;��r{'}C�e��*,�.ӛ�_Vc�4W��+%g���F�-6�t����?d0|�d$%0�>q�_���KlM�����?�8�Y.R��F��6m���ʯ'����-�X����E�^���?�++�G�P[�=�EW|�8o��w��- �=/��"ꩆj�X�̸�l�t	�eG	���)8X1��uj�����K֮,GI�@���!��%�<�4mǍ_���Z��-dE��4��[`� {:�����;���;�I8,�4��1��)*Сu4�ΛHl�L�F"<���8��j���X3t��V��6�p���oXM�!i��g�S��՛Ś|���f�K�%��n�N׼�cZҨϙ7�����r�A�`��L�7��H.�Z�e��8�ou��h8�l��b���Mz�A�����n�,�ǁ���umU_�pdv|��<��g�#=�2�������I3��ۘ^����lM۴� _�Xv���ܩM����r����l9�M0�3m�aj�z�M��>ZZ����	����Pm�4�mn����D������q	���]��lGZy�2r��|�'o��=7���奎���6����r.f�=�"-�&�1�!�F+�1sGͰ��@��.��`wH��k��
�Z�u���@ڥy68�����8\'i�s��1Ec�Z�"v��E\�k/f��?���s��5n���{*���|Y��S��`�D�%>��j����	t�\Q��~Sr���F�7U�t�]n-�#�!̮D��a"Ѐ�=y�TO�8Ѷ�X�?G��fڿ�Q�Qv*D��w$������$"'�C�b�)e.�V` ���@������#���v��1��nD$��8��q��'k�$�D�	�op&$%���8"����w�O|~۲��c6~ԑ�D6Ɨ���Y�@W
Z�&�2��k��1�>�a�N�06ڶ{/��X�yh����՞�e��c���L �c��w-mi��'� f����te^��?F��ތZK^-�E�����&'k_��|b�)�eu��#bj(>:�T׊!��b�� (�d�$�Ǖ��}~�ǉ�M��^�+���k��M�}��w����,qF�0XA-xN9���C���2ݕ��s�7� �K2�IÃ�1�&�
pc2̦���KjI���0�3*C\>z���j�T-�A��:KU�ѥ�t��L��	]4CI�,F�Z��d�=�&�L����}���q��I�X&(�.7k�?K��!҇����1�*(lY!4R�GĢ�%j4���
��ئͱQ���7F�W���7�JO�X%,���� *,�H��7�j�cW� � 
���Oi���CJJ��X��z{(6Y� ��ƞJ�i�7��F���{����_�N�͊�E��k�w�i߳�CF
c�O
�o��w\�>�c�+^�7��	k�p�$��6��@���8]X�f�x�ŘFۮ��<���q2Ѭ:ߗ�y�9P*TM	9�bu�=Ԃ
q��F�
�F�T�!~��4�q㌀C��M�4�`ZS��s�+J�D�a�5�6�$�twu!j��U�9/-:��o%\��C��>��\X?jR�t���m�t~���(��od��W (��ٌ��ص�{ï:�B��ϙ��Hr���39��@�@��E�jmAu׊7N�����3?�C�=ggְ/Y�����P���k�aI9B_��7��mb�|MƜ=����Y�%GO�t��.�M<@M䳥O�=��g��v|�j�����"�t��A2m�x�-��ѿ�+;��Q�L&~����k=Ŕ�����ҋgH|o"�{t^�G�F�k.��sF��JT���S����U�Z8 ��?�
:�d�o�L"�z7��A;��١���`/��V�*ӗ�hb����'
G�Y�q�KSp�������p(N]��*/> ��(�fJ*�0on8|�ݜ�_�!73a�-��Y4����y`:۴$B)b)7�������;��9S�,�h$�TWf���]Ve"+M@qCf���q�n\N�Ԧ�?�H�gS&ǚP�67cﻤ�U.@�E���MlH��E/M����J�_���d�g�+���'V' vL�o�RǖG������TB�+M#8%���ţ���u@�EY!�w�uy�����}��خGD���q�I������z^���	#Y���#`l��Ζ�k�u���?�3�I�Fr��a�;^B�/P�г�~z8���I����
�� #���Յ��M�����=��Vm%h��Τ4�G�@�dK�E���(T��@V/җ|%�lh>�����H�ax*�j�ϱ�a��|��v[�S�;��Ed�PyµmF��g%�p�*D��!�
k>>���6�M����0�����LxsD�S{����&�o�Sy��K+�Z�nۥV��|ܫ�qS���e� J'�B%��7��Kx�	3�p>�=h�f��rVCo�)�kY��>� T�g��ޫp�sd�n*����b}�~>s��q}����c������qN9�7�P�ܜ�C�6�q��V�$�?�g��#B�V���ѻd�B�[����MnM�MlE�
�2�����;�h�]8�:BKz��D@@�ٴ!a�t�����SP�^��h��g+��i�:��0m�����󌞽f�1��S�og6�;��W�C��e�wT5�-�,�$��oV�h�ѧ�R���4���h>��e�af���+��_Al������L62�#�Я`S�3"*�1��q�������ϊ�9�UN>GZs����6��N���Y���y�^H�ޯ�H`	�5���@��"��*��8�v/���<�^�$��B��\0��y��G����W5������$��Mm�e�e�6CI�9�H�E�4��Ր��|�dG�����RF���b���b�N�i���@L�1�wB��~÷{� ��j�0��1s״�Mo����!�T�������j,�!b:�5V2�+?�����q�"b$�������`��U�V�������	����tr	gI�Z�ͨ�r0Qh�5l��p�����3޼�tA��|t��j�#+h0*~/��~42�u�%kx���c�&�-��X�����AjX#@!�*�G]��u�1�C�r��ks}B����2V�v܍�U����<�ǆ�a��0r�(��9��U~��
���Ϥ�S����缬���|��M��I�T�5W�� ���+�+�����k	�(u��iDxg�b���Z��6[s��c5����\��n�:.�98� ��g�d{ br��B!����S���Q���Ͽ�<�a�����I�	�A�+�pe\%��!�N�33�j_S��BsopZ 1�ѱZ���UW�LH?����(r�$�Q��k\�T28f~�l���K�����?��9�Y�w�����ļ��7���rl(5�D'ň;0��H�<�T|�sP-�p�U^3������aכf<�����'\RbЁ<�f%4���)��ec=`sMϱu�m8Mh�8i��Fb4��`��� Du�1�Ŵ0*�xhA�)���E�#X�We |&;j����]�z�</��&��_��q�z�Zg�O���A�j���Qѭ�)�5I	\Mj!�-�)����p,�2�*Y�n�z�(�N�WW��p�_�콂w���?x_�l�o��{�O�h���x��lEL�1��G�3���1	�op�K��<����Yb��?���R�l�;�7S��BQ%{*���gm_CK��}|s��P���m<0����/2�N��ʛ5�j�[��sIӈ�;U����'-�r]Ϛa���..���փ��s��_��!r��˻�~kY��1?"vdR�d�0���H)g �w�M�ɂny��ѝH����85~6`QF[���^J�Ql�"n�-�� 81@XX(��{ۀoÆ���04h��5	�z�͂Z.���h�e���2��\|���W0h.�L�Jx�|;vk����@l1��X�����=:G~�p����E�"�k�%�ȰPά������B���Cf�i��#Ps7�?�(����[���p�l��&�6{�n��k���ȍ��$�3���m���|j�;�r�G���D^ᘣ ��&B!�}-8@Οg�|����n��޹������=�a�x�?N3G�w>H��q9dA��������=%�š���VC�>!|1�57��F���͠�RS�%ף���q���oݻ���N�Zv �޻Vp���6	�p��I�vp&�� ]�$KE�������9�nb�7�! g5��4��N"qox5����N�xW;I	�M��l��-��V$�jf�+��[l)�~W�8wO�ĩ�{�扚��w���Ǿ����"���EÞ�ߚ"N��*�/g��u�����7u�N�Cb�=���;�6#������g�,��E\��1�R�j@і�����ŋbA�� ��pAY�c������L)����d&���t�=|�?<�Rg)D�T��2E0xt���ٯd��	���iT�M�RJ�r��4�g�{��Fy�������Rj�T�ɶCe��ld�>5naEW �r�U�g���=K�7됸l�k}�
tJ�@�	*0�i7D�[���]��UIܺ6���P��鸢?���X�G��H"B� �T�����U�'�O�O�0`[2o�T)R��*� ��\�̑ֆ��t��#,�un`��^�K�
��t��_,����~��n�d����Pts9��w2�9a~�*�d�7�ĸ�G�f\�ȁs��%�r�:�|T�^>I�aЈv�P�����Nc�i�jpN3��I���ts�} "��-/�$�>n�� h|�\�N����R�^&A��
� �&�Y��AgjpLN63\;�/��>ӹ���ީ(˙'�>�� /�z�v�opKJ���EQ���jX�zp��)>��ҸH6�#��8_IRp���n��nsvw/���8�I�� �~5WC5�Ԛ;�a/�6�+y��\���L�k�t*-��,��j^_[%ϥӅҐ�	��s�P��a�o�U��O)(��y*Ԁ�妷�&�V�ĳ�d�G8;%DT;A<"&�����:�Xܨp�ֿ�vI�K}��4�Y���<Q��������d�e^E��m�i�ֈ��*m%�>���oڂ���>VX����y*���&�i/�䬑�&@9�{I�\����w�E�LL,x�,������ d�I�H��N'��D�c���;��0.�@�2��80U?;���ji������-qAY�����[�5F�]��u��Z��,�GPX�t�"��O�^ L�RLf�u������Qel�s��(��e&R��ݙ�h(��f���F{�\c�0�~�mRxwDy��4����7��>�<G#�I��ᔰ�l����b��l˨���� .S�;�5,^lݘ�:f�8�����͠���E�,�A���I(����W�ӠJ����(e>sQ۱ �0�r�$>ȕ��l�gf�%3Q�ۚêc�s�j��=ٜ�T�9�$�ʑƁL�����1���R4Z�D /s��f%aZ}x�����Ǌ6w���G�˗���/\fǒɕ�ß��Y{{��*�z����&$�*nK����n�߅1T�L�'���#��`$����IU#��
�Y&�uW���\�JA[��Ǳ�p�����S%k�)	�rj�����o%��y�?C�v�G^m��׎�~(��N��x�e��F�dc�5��q�r�j	$>b~�H��jt�$�9H0����nG��PihD㭌f�ٰ��X����zi\�>ug��1����t��|�C��[=���Sp#��ת ��	�1�gK�+�x$�	p9n�Y����)�E`1�l.�x��k�bY�m��w�l`�`��I�sK�H���1$N����j���9��T���+��1w�W�=l�]n�ؠ(^z�]���W�`��}H1��c�p�w=r�q����׺��j
��YY��"�G6�qs�����-��
	_�H$�堙���]�Ǣhw����p�ݑV��Mb�F�CF�Wɋ]eR�J���SB9�X���-�.$�7����c^��1)Q�0C�U�ʓ~�fx^߆Z1QB
+Qތ�3\��J��BO|�6z�̙u�N����eZ6.�b�d���&���_Z�g Y�|��(~e�A�ǐZ�ֹeM���4��1���Jg�4Ӗ��-OV8�+�����,�2�&���7d����u���6ae"�
_5Io���S(bG�A\&�(�,,�Oх�bĂ��p�_}���3J��O�E��^�� m����*S�ƿ�E�)@�_7nA~�O��ˁʬ�'�R]��~�#c}�b�'�x�@rh�Tf����2�k2?}���٩�ZJ��۫(��� 0�a��{G�Է�R���f�� il�f�P���1�&B,	b�D1b��Zi��U��/'>o�׉$�[�?��Wj�)U��c��[���Ӷo�A��$-�]Hǔ�Ġ�n�2�>8I�fr|'d��a����G����]��5��A ${��l��Г]A4�su�OؚH�V.T�gh����Y~^�@�:__YK��k���9���rO�ĮU�h�L*L⤉Q��ml��G�s9�0�x$�����^���<)���mt����cړ�A��W�T��-铀x��~���`f+yU=���u�߰���Wƪ�W�j���8��۫�Zi���Jk�}URgu��N����*Šw=t�^Z&�w��z"��'����Z_�C����-3/�m��,Wd�|�����$����W����P�1��"�e��

v]��y�>F+�ݗ5{(��ˈ�@�����?@�Z�b-�*t�n5���j����
\�Qf�����[�_���M\���O��=X��!�]m�x^s�/��*O��s[�a�<)F>�r�U)X�&ڶ�*j�;R�}k�]�+V��`L$q5����_~P�T�}ku�}���6�G��9�r2�K�# Zlȇ�Ӳ geH�����m��k�UE]")�� �l���ӛ`ͭ�x�j^�����7��w����F��U�aWK�ۘ��x�w�w23����J�(<����Z��Ll���B�?�{��Q?��
�r�R���].��i@�AZL��*�C����
f�l��a��޽�t��x�z���hzYg��3g��D���}�:�E���F~�Y¿gi�
De	u��䝺��N7��!Uؒl���QQ�j���Wv�Y�nm���FQ�x��qq���3%��+Wh'�t����X��m���(���E �}��Hxԛ�R��Lzn7K(�׭0gi/�i�]�leCl�(U7$� G�37i�4��\�e��O�����2�?��k,��0�|��S����X'U�-ӕ�gn���F��ʲ��d����9���f��º�������۸O>x�b��8�Q1%"�������	��4�3+ӄU:��� �5�e�FH�3�ws��i��P�f����yC���|/�N��al�CG��ͬ���SW�j�*��,�/r�S��3��l�S�8�Y�l� �|����<y�מտ����]�*�b m���+�Z	`��ƈ�eU-{f��1�]f%��`��'���Xtʵ�[�o���& U_@�s�D5
n�@m�j�y�����ki��uS�P��W ��^��E#�Ne�8bl�e�F�<��x$��U��c���@�@A�(ˮtu:�^�@��X#H]궧a�#�d7[Z�%Z@�1,"Y��3��19+o�z�3�T(�Ql����_/V�c�o������5T/)��UNN2��F4c�Ӷ,�nt��������8���e�e���UL�t�x-������+��O�	M+���B�[Q�
`�؀j|g���+&�O?Ł����bj�;���e��T������C�8<z�l4Y�9uO��T��֣�"��y��S�x*�I@B��z���s�2���,�,�rJI�5?�r�ۍ�wM�93qɔN��g[�9 {RW�d�r5���F������ayct�c�c9��J��jM��#5�Y�l"7u��3�o=�* �uJ!qAr+��ʯ�v��=k~Żw��HV�_Ep@�qHH�Fׇ�m�d#����b�����P�S�~ct�{"�6⿠(�����C G��;���=�Oe�1�ߺ��I�J�E�ygΜ:��r�A V���"��r?�y�s�h�ߗ��WF(�KJ���j�߯5�#ίx�u 0+#,��7?'���E�I�{͈�#������Vg+�		�,��d�{<s�Ҟn�;���E8�h۝���"�jς&�aq�
�-��%Zf�a�ux t�i8,�Ff�تs�+؜��+�Ŕ?����Z<��kv	g�N6�7����[ŭ4���Z������JJb�å%Ѽ�l1���0�|ޫ �����A�Uk��P0Mc5�nÃ�.�F���7��CF���6 ���ʋ���f���q�{<��� ޴�덣=h��Kթ��^d��"�b���i�K�aa�p�s�wٵe��n��^
�4l�ɩ2��v2�O���T��}�@��RBI��Ԯ�uT2�$�<���8 JF�Gl-�fU8sϩ�*H��l�mc�Od4���Mh?h�0V�H���Hi�h��偳I�q�E��/N�J!�3;e��I��+DɅ��t2}.`q� s��W�|����k�ws�A���آ�N3���T��Sm���Ki� Ot��$U�uK{c0��3���sk�R�Y/q!��'I���������+w4%����F*��k�Y�DR,�.[���{8He����o�@s@;|��b��#RB��[*�ؽ�bwk䡕�L�kܼ��Lk9M��ŉ���ҡR���|��5c���ф@ܦUYG�м�f<�^�E~�Ec0114����o�CC�~ Gq�/E@k,��*b�VWSp�7��e�H .�qrP}o�<q\kk�*;3�����J�Î+1,1�$i�s�{o�C�F�C��f�[i��F���6}��ELS}��M�)~#н'&+�����j#Y����@�)LL�H)�L����n�{�a��)���ʅ��n�\�":����W\��a}k�i����J�k#7���%ߚ�!ׂ�_��V�m�/�-��Y������!ϭ�����u���Z:�s���p�����޻=+�1Y<2A3����sM���{�����t�5|���J9;�O�R׬+D�JL�a}��Nৣ���&b��!�����$:��2^/��r<I¢�)��{�N�7#%��k������pI�抅@1Y�=셅X�J]�8�T�S�1��ZT�?!�A⬾r�&�l��tyXN�V$�����֍�!��a)�\#�/��6�l���Fs�l�y·Mۈ�f{s��ݎc`��E�c�9b���L3!Pt�����KJ{�(ӻu�Q��>5���	@�S{!�<�����a\��v��t��oe�)��Y�oZ���������͂�+hzU��ܼ��@eѲ����]� F"@�^��R����m9�Y�w��I���m*
~ZwU_�lm?ʜ�m����y8��#���W��<8  4�5���%C
-O|_���ϙ����c;G���dݫ	A��x��qK�����E�鴟��/���d�[��J�隘��.X�kd	��(t��Q]��T��VGo���bW�H��{��T��~z�"A������N�w+��E�&(1�@
�1�	�e;�I,Z]N�c�3݁�[8^��; )!���G*0�sN�k|{�R��{�|��NR�%��HJ^EhqѵBۨ���F��k�U�7mŵO�B��!Ի�o�C|>�<P���(�u����'u`�	���b�fKq�����;�$��H�5��,ձ&_"~˱=�8��!D�f���֜��o��Շ���8Ɲ+�6�a�,�o��w))��`e��\Aқhe���|�찙��ڱC��D[��y;R	�5gY��jt��k��~*|��dyH�>�vGmA�X�g����
�Y���	���4���@:��O�i��X�� ��-�q�o�	5�V��q^�P�N�A�Gd���P�'4�\���J��҄��Ԣ�����3��8i�q7�L�k2*�d�\��
c��V<�߯{�Q�.ω�hh�<$�V��氋���V������H
���WV��M!�U�*����q��z� ��#PR�ԕ�煵�9@��Rjx3$�V�G��1F«�}��=[g4ё's�"��>��<BmH��|ĥ�*p}D ������o)W�U�6B���VD���Y1�+��(F�`�m�|�&�5�*��o�B�`$ ��LV�.z.\8($R�FD�����v@-�كO��Wy��4b�wo�$7�O����ݦ��2�N�[�j��%�F;��Ku`<Y0�������N6/��ϧ�HM]��8E�E��W���ڬ4F/del缾���"�k���&��W��C�wy��|��EU$�G�qu/����s [=�H�b��j5���;�� �1��� �C��ox�m��]mV��������w0��/��񢈫���S�Z�U'�8�?��y�fP���_����v�K��<]~7Kp�M�#��%ir�f�T�.}.|��z�a��ce`l�;���=������8de��$h�n ]�|�����:�Rm���.�c�, �F�^��z��D�@�ͯi�+j�=�Zi�C����Ǝ������=�v���T0.p����bh�T�D���s�2@��-��<�ϮC��a�.��~h�N])�ػ��ͭP���<��w�r��(g���1Q4�����CzS��)�~6A�����G���e�"��]Wp�A8�ǥ��>єt����>��L�=�d�I��Q�����ב隼I�n��@��[�g�뎗�=@v�~m�4�^a�ٿ~"yc0���Y�~��K�|Z� G��/�,�VtW�z�Y2����X�' ܫ�:HU١��f�&ͯ�����}�Eu��r�Wܘ��o3. ٱ�� �sm����;ï�ee��x��QF|��ؖ��QbS�%
��A���Fc�ֺ����k:�'K��2��b���NP�U.N]� ���[�_xe���������:Ez槯�g�:`~�0�=�K��4c�~�m�~�f�5K�bO��}��z�����y�pv��i<l$T�F$�{��t��P��8p>�S���m��؜S9��G�\����&�'YpF@E�nl�Q�p�+���UM��K��M�3��-W�Q+�Y�B�G!w�24UN7fw�����k�?��#bv~&�"}?�p�.	&P:�~���'�aHT
)K{�4Y�삫f��[1�u���UG���έ��x���X:�bo��| �B�)BY�Ҧ���)��%�R������ii����S�!�y��Zk��@��7p�jm6h����8º�m���lԓ������nU!�mV��u��d���|����e���Y�o3�D�\�>vcqM�d}閬/D����"j������E�J:{�1M�iO�$�?&
@e�����h��[�������إAK��C>���%��>�ww�'�KҊ;�whF�U-��XWB�/��'#o�}۷H��U���ْ������y�-��1M7��sx�Iud��p�I�Z�Y�p$!s�|L��c�F��6V��>&З �q�z�̌GN�RdP^[g�#��O�����hȻH�;2�7;i�NM�rA���8��}d�LE��zp�0j49���s��{�c8m˴)���NEP������"��x�F�m����t�OHw~@����$N�Z/˛O٢��Zox��F��0j�m�j��Q"��H�����7��#4 �J�L��9f��e�� x_�&JQĬ���y�=X��:ᩑ�N]0�����q�Y�F4���qz"3�a����8z\��ufDTb��Ф,eh�}��nk����&�/���&�O�ҜK;����)�������|	��A�v����A�d��UW��L���tD���tS�%4����#$��r?nA��7W�-���H�S ��X�e7A�N��[��7��9i�>=�e Җ\�O�K%l#:�=2�@�� w�J�H5�]�Ya<X<�&����D���)W�GpU��qg]Z'[u��[	����� ���m�a9�l�8�fR�ȍ/��u�=����)!�Y>��g�yuA&�A�����7#�qt�'�P��'0_pmqW=$��xΦt�B�b��'Y�U��{�K� J,�_����gG��:�'6[�g�S�5Qˣ��h�!0����b�n�8 zk��s2���R�
�,�k���@D]��\I�UA��o!��0@D�C���%�=�0��$��aO} Ib����[�h?|̺���nl������6b�ʁS���n�T�?�z�����!�[ ��,Hx�=���p��%0� ���0��*<
���TNx��5�7b^'@���aVܒ��q�y�������咒�m'N����0QUb�[8-]IS.ǋD�ij�[F�
��9k������z������_�!l�n��[�ܔNAp{nC*�t�d�{N��V�h��Ϥ�e����m³�pi$O�x�^��e�Y?���K"��bh�M����n�kS�ꕫ���2���F���A9����5��~��ܬ��RǬ��υ�~a��/�{��v�"��������JYD�1�;��C��@��_��S�T��������E<�(�8Q^V�5q��q�Ǉm-�־�3����`��bxrvH�w�3��,�!��:aV8B��C���BI�xE��RĞM��7���9pX/��X��Ếv9��D��_f�t'���*�������iӖ�,ӝ�2��8O�vM�b�K��j�� 8��p��{p+�c.�_r|���Mu���&g_J!>��h�A`/�P������`)ݙ�C(��ޢ�p<Ou��>��x�"�W�Q�+�D�48Y����bd�ǨWI4��N�T;�2��~�7��BJ(����W�f���T�0N	�=,ö<�#w��q���ߺ�6R�Ht�n��HvΣ姞_�3!�s9��j=�ā`}��7�)��a�O[��.^�i�tڪ�S>{Y�جS�kh6�,�ט�5�v��p[B��&�g��Ncs��ɽ**��-�@� ��n�Q9�*�!9:,�3����I+Θ�B�� nZ�K�v��g�+Kk��wy�CB��Gc�r�R����s�G}7�{R�x3TQ�<��&���,C�TuW�bł<�ʨ�(�9��7M��k~��{�%��-�iXu+r�u�_Q_��ᨺ�e�C���{���������� ���'��'�uN��z��H�ON���!�؏��
Z�^���.�Y�:���J��q�wp�̷��I��ѭt�����^��j<�k�䂙;��<�p��`9 ��������/L(C[x��}vk���x-��P�I�8	�}x+�Nq��|�O�JG��K8�V)��N����E���Iס��2�ħ6^��t�ɧ�36Rn� ����1�@56"�_W<l�HL�" �	/�^�X���Tn���h�U��uS���Ȝ8� �0������C�A�l��d�Ҟ1��K�x��i�
.�i�Q��t��3#����٦;xVDQQ�8\Y떰J���������'��뱧z�h9��� ���T��
��P�DAN�j��Q���X�ɂ�D^/��*[�P�*C-�&�J)Zy��	;n­��i]zj�`c�Anŀ��:��}�cP�*4
WC>Ds�UlL�z��Y߹�-p��6��|�s;��m-,����u#�g���|އAJ��t�!�'�z����[�-�Ü�0�@�E�wۡ8��[G#��]Qj7�2�������zI�f3�����u9�c�9�3���d��ހ��zv=Yt�C�KEnS�����2�����#al��&��*�a�v��ʤ�ġ�K\�����X�����$'H��Ի���.�'��@� h�@/�M$�y���(-x�E����ۦR6<��Ĝ�6�!嵯�Sb��e��v��LU�y6��Lũ�DV��,�ӎ�[��U z��	���lryl!��!	ؿ)ӽؑ&W�lV	kB����s/�U�=�u���]��^Xޅaf���|�<��\��t̽�㲰y�|pR@�ԟ��|��~��=���:�\�{���hG���j��ow�e#6h���'#VT�a&�	���v��6I�З�d}eXN`��;s�d������GEL�D���,�+����ňb��w���<�jX�1�0>��LaT�k�����G�ci�W1O%�m�Aܚ�a�����b�~�󩡺xI�b��~�ן�ThP�^tvѮ����ߤ��۷�P��Hyp�`m�?����X:ez�/�p�NDwCp�l �q���J�z��>*0}�
g���� ����x	��� �JG��1*K�Yf��'W��c�)t�x�7r�F�$9���dM4�I.��ҭ����T�Ōشb�����<�f�RсQ���Є.J���6�����7Y޲;�Sa�;|>?;��I�h(���;#7v�V#�F���BNўQL���g�J��U��m���8̐֙M������iIՔP� _�md�.�.*��=�������#��Qi��]h�/ 4I~Œ�R�;�VNaom��B�䝒r�����<�`�b�Y
��1t��br;C��O`��Y={F��΄���"�I���,�?`��+.���[5�䙇aʶY������Z��VF�2\�$�X��HT�^Rļ����(i��ݙ��l ���?w��:�%�-���]�����QG���%T��¡�z�
8i�Oe��M�Ո8��C��)�H3y�� ����e_�~�y���!�f�ۛ�ȣ&�l��A^�{��L;�<�gFf�jkLɖ�d����O��8�G��U�����[u������#߽j�0)I$x2��-����E���H3��x�e0RީRq�)A�j@�3@���E�!C�\ -��L7�s
�4e&i��DD���g
L8�^������EiC�\�x@c�m��.͓\��J�w��B�!���x㔣�,�W������b�
_�yq�lV�y�� V�V�*��߇�z�z�v=9U�'��x��k�`�t; 7��ѰSL�����b(��o�\�PU�Dݍ�e$�ny���	\ �	Y$q���B����vy<���=Vcqݟ4߼O[+�ӧ�s�8����-��TU�ƅ�����_��m7����Q���h�h5u/�Ƒ?��"5z�2�^)$F|��-�W�n��u��q���Ú�G��,��uu��D��e�zX�Q'FR�.tx���z�4Ճ݃��]�Û�q���\�Յ��P��f��9�@���NN�l[*�K-�����C0k�Y�ո*��I�?��=Ʃ~����?{��o�4�k��3T$t%tͯ��$zݟ���	h�Q)�
���h��K�QxWR�#����W~�(Wh��H�y����?>������{c���F8e&QM�O|!lނ��sKV�'��("���� ��G�T �wF�� h��q;��P�F�芮�P�72����^%lE�P�;U*ԫ���%"����F���l����eY�b�UI;�_�8	'��8"��)s��?�^g��
-c�?(�����R��	��O�[�:�A�x�7lO�"����~_�a��]��y�n����xAz�,�M�h� _R:� ������+� L�� Y����Q�8,� �g#���Ay��3Eɏ�J5
���)�$�.Vv�XM�����ФF���@�Q�ԡf�B�ɾI���|�i!��a��=G���b�x��&*/�:���&�}*|�1����R�����Z�?�Ǳ���������,�{�U��U_l�u^��К���$��t
�Y�֍��=̝��q�/ֵ�!.	�+��k�8�_�	�c� z5�#��5��rj%�)�����0nquB, ��MU`�@f�g�7D�w�(��7"�M*�tD�p?+_0D��u��������ρ�t�}�0L��%|�/�������KΦz��D���~���,"/�}��Q}Lz��uܢPG9�����wJ�ք�k�F�I�x� ����/@(��J$���A4��{�F=(L��E���9^�䙪��$j���΋t�(7�(pM.���1�J�p�g�M�W�� h��Ӄ�c�}Z�XF /�4�sl6��pF���.��[�A](�r���@d/D�zE����Ս�(1Ђ��7��d�)Z$�"�2Ԇ�P �}����w����FM�ج�'���ŝ��A����O	�,����y��
�f~�x�/����Q��+G�*�b=d�n6{�C����E��p��P��f����.�b�.BP�]�힓!d��������_�Ǖ�t��gXG�#Z�`�O����F�Z@-s-,I"[����O��oU$�
q�)��s����1��B�ڰnk#�a���؞����i]�^��.L4�ԓ���w�H*�t`c�� Y����c��7�Q�2�z������p����kw��On�FG�������ݔW��w�
uT�ڰ�fA�s�U����ں	'�� �re�$s�4�99&dy�ܺMl0A*V��2�M���8g	=RU��R�+�e�pG�N��3ۥ�H��2�(]�N	��B��%�Fg��
�L��"G�Iy�wE��MbPd��*�M7 �k�=���8������g�W˰��[��Yܐ�bU̜���4�l{]��z
���v���vW1��wgH́�*�����>�B��?h~�n����r�	hvf�Y�.~e��[��y�:E%~�����B���˾����O���6I"Y��&��k������0��lsL=�D撔�U���No#v��дI
�����ԈT�20��mx��MK0�aJ�V���S�#O6�_3WKAA�L?��:���5����n�L`�78�Xwٝ���J,0?i11��>��4�º
���BY+9cS��R�׼s�i���*;f�J�Z���jO�xQ�Nw!u����u����x���0]�=E��ݣj<�<��$�*�l��D�TC�Ґ�*U\i��ZJ�&�Z�>���@�i�f�(��o�~�AAF�J�	��Z)AY��O�$�	lo�Qf��#b��u
DEg�+��b�d}-րKbc�?4YD;u���j5Iw�$ж���ӭ��[�q�a��������5� e�
S�t~�*L�(T���z�vG��D�ۦ��;f��)�E��:��z����t���E߶<IcT�#^����stj�y����W��P��_�������Q�D<�����Y��M�+�9rf�g��b�~���i����z�d�W����M��q���F�/���Nf��bٺ��>P�V?�����)'����iB��ȫ�ya=��s�@�L/=�w�,Uw��%�Bi��u?�P�ů��1�6���� }3_y��[{2r̿�M�n^�W@� �=
?s�P��9g$x�RNVlf��F��0�eO�˰����Z��ڡ�c�g
���#z�Y�5h&Y�_‪N�㻦r�p͂^LG��c����O~��z]n�;S���d�|�G�$"��r2_F�T���J�����pF���5|�q�.Y�@�K��������������[z�3�Hi���0� A�5�.'��Q�Ȭࠋku�;݀�.v1�)Q�?�oq�5�~]��ڇ6kU�����;��t�&���UP����9���{W���ЁV�&��LW�l��7ER��y+� �u��M�0C�z) ��£~���tʥ@7$L� ��0��~��U��O�e x��)Ɠl�T����?V>C�o�`ZƓ
snz	��=/�L�/�p�B[��ʜ����t���E���e�kd��|<\��7�V98��2h�WTi ^��#�����׹@:��/��U�V#^ �;�h��=H<�}��;�Y��:��	�yV��aH� ���h'�ݸ��.	:����K��˔_�����Ny�)��6�ei��r��3#B"�̿DL�%�䄫���t���lu߈�C��l=wB!���>r�Hs������8��S�\%��r+��Q��	�9"/�M��<ܾhL ��7�+ξ�E9Cgh�.%��s���G(U�X>H�,UVMy"�%���/�Te)>pi +��Qx���\&�W��߸����C6��v}����P��8��[P9m����5���S#R�R����j���k��O�s(SU ��=�#�/��J����+p�,�� �Ⱦ��h��z��|��T�L����>0ߺ:-'s!���6�/b+*�F�la�E��A���/T�s��&���)��!\�w��ώ�q��w8�ćO{�:���+Y�y*�	uy�8�7I|õ�^���]�'�Z�G0wxȰs��a4Qy�ěJ$��
f�'�{"6Q��f����)�P�Px�������Jt�`���s�_�1�,ĝ�R�=��O2�˚S��Wo1��N�2c�����Wz9���c�`�(�.��v"8|G���"H$tқ�Ξ���*i@̺��@窧��`��4�n�P���>Q#�u~��(���w}Hn�
��������ui���aͻ�8��s�1U�����7sj�,d�
]O�cB烛4��'kN���q|�?�2e� ��xT���ز_4�,9C�z�ڝ��+,Q c��Z�xFi}~:��<0i���(8�~\���平�f{��	��5���L9^`g�a˷�n;?͵���@T}
Wh<ƶ=�����>�VX�+~���kØ���%�6�spfR���1R.6Dz�?�'�&Iw"͖\�ȁo�ҹ����{(ׂj��'�k˛#v�;�/�4O�E�Yq���
��U[ѽ	��2�m`��H��3��3��p�h<��Z�̗ǋb�zr�H�??�����Y�@|f�ױ%�	6Rx
�k7��JnѶ)�d�b�_!���͸q�ϨQ�{�3�� �̢m�_�t��� w�S/v�9#0X��CiT5'z��<�pY�w�Ϊ�g��ų����f\�0�C^gx�Va�(*Z8�{��={6���n5�\�O���:]�{j�/Aȣ�5;bs�$zl>�ɞ��[�.9@�JT=�DH�� �*��h��3a�7H���vO~����^E�����D���;$�s�_G���� ���|I�����O�g=w��Ͱt�ٴ�_�3��x�.cƙ�f��G���[�E���_� �̚�_ �� � c@��G�m7�>�3m����Y��d�n|k�Ϲ<�W�w���m�L�@��%�j��_����u�;`�=.|pR4b�^/�}��;a���X�2o�˿�~�oS�Aj�#,�6h�Vb�Dl����n�\�)Wb��X��ҢkZ����e�?Rܮv�ڤ��p-�����m�c念�|�j��2z(��c�N�_�d�.�E�-���ݡν���b�.�rǐj�[@��]�����,���l�EV)kR23��i�A/�	h�X�=~ef㜸0�k��X*��>�֩���"e��w�q�>��pN��w�T2nwB;�����=nJ$�q6"T8\��_��K�Qq�z�BV%�T1�-$j�WC��=���;�G�$��c�Ч�w� �d��i�mO����K�! �Կ-��J���ݹ1{�
�)���z
V��ω��ۄ�w��op�Yå"�.zy!͹��� ��ڹ\]�=^��l�c��D� Lqz�f�t�僒��}�r�:���@�_�~��"R���Vf��1K%�S�O2�aMrg���XQ^�h�����������#�a>z�GTLr`�^�8�O�2�eS�z��Q-�0ݓ��{l�Le���/�i�Z�?��� v�(�!r�OLY�?�MIN�����ݽ�d=�uvQ����	A��Sh@V�ĖߺZ���yI��!Ru��-�aCDc!����~�4��MY�2�'�	I����(��Y��zB�-1ѣ�g�N�����b?6M~�.��TkYS}!���i�fQ�)J�Dz�"o��k�Ҡ���������3-P��[���\��Q�����}��%��V���@8��6d=$�)k�sffT+�Lo�#O!.���$�}r�R{Z��Q�^=|N��K�P�@4k�v$�W`�W���U�-T-�4\]�ց�2@.w�dH6b���&���I�P&e�r�P�� ��־�_RGO�Z���<:�y��E>2~�N�j�d:�� �,�>�+�����y��uE\�w"f%��õ��>�>����Ny�iR��*�5��m5L�r%Ţ8��!��-G-��ɖW��L9 ǁ�l-�u���a?�|�r'55�R�7���3$˙=��ftJe�k��b�z-�+`J�
���"�s=CeW|ۤNT�̰��Ci{b�Rv_��cAXGۈ�P��D����3b/Mj�,�L��}����;�6"7�8\K�\�m0�������*����CS���E	�M�
P���t����(���#N[�X����.�$&���Os������K`΀�L��W�:��s���L�{��N:��\��8�w��73�W�j��V�u!<����q �d�2��r���C/qm�%�+��d�1,���2]���U�lK��-u�<%�থ�h�LPѮ�)� `]��J^e��c�C��QXk�>yn EmR�N�`���{��Mʠ5��;�䡻��j�f����?�SAc����ҫ�M���B�og�1�9���]���d�ݢݏ�'�,�#k�I�	�Vtl��@ R��ȡ�q���WDoP&�.�É�?4�Ɖ�nA��4�����,�;�0'���QÌ� ���D^41��\3������=��eFߊ���Ѭ�a�u֕�vW��9��d*�GE�����ֳT	9�ƤS|F��բ���H��Š���hp��g2Y-2���'G_��^,���3���W}���.e�'���པ�j�s[h�b�py	l��+"��(U��ډ���U�v ��9��[�=���/��V���e��r��UO��<q2����˩��r�6�7�4m�ܚj�:�gm5?�7x�\4�My�ؒNp���R�x	�P�M0hZQ�3/�����w��^A�����&	�a�����_R\j�����V�o��~��3���o���asB��b�b�<g�A��12�S~g�U��MP�x�?����5 &�ֆ� ?��o��t3���.���j�����ik�qas~)ܰ1�%�9.��>�8f�(�����dsҦqA'�:l�+��Y�m�5�&D��=�����rа�d��a�5�C+؝�AGx'�o7}�=>��Y��8�
��W��t�v�wޚ ���2� !ε�{?er^�snס�k+2*L�(��"}
����t�0����3Y��:��npp���+E0�e�ǟ|^&+B�����2I�������xe��X��qr�<�]0|��J�Բ���X+; ���*�ѥ��/���$~����Rf��0k�[ŚaJ�	�8x>I3���2�{��e*&xB���H����s+Aâ���iq�7P��;j��\���&��0&�lV�0i����B�=܈�$��a�ԕ$�6`��.v(?��
�±���<;��3�A��ĬΕ�S݆=&��R3v=��H+���C�3�us����I����C��0\��M�B���S�E|�-�~GB��'�2������P��d��\=�������U�#x�k�잆�>���r��}S���h����.>X�ɢ����� ��7嶏��;��C,l�|ܗ�g���(���EHK.�N�0O	��;D�J$9yh6�e��P��<z{{���4D�d��.��3�Dk����D�I �H���r�Q���"�����Ì��{J7����e�kl�*`����aXE����7 �U�a��U�	^�*a�ij^��6rFtĀO�A�:-Q�o�6��u�$\t�����Z&���e��$�4�&������s��EC۳���#�E�*r}5���Y$�O@�@aD� �4���.��ő�k>�
mԒ 4 ���m5��`��bZ'�{���GD]2KH �v��e�S��<��fݨ����D^�K�N%���:'���ӄp3�f`s�����v9ֵj�z�b#oSڍ�\��zF��9bƀ�%�Aݎ5Vp���j?���O�(8nޒ�	Ȁ�p�1DO' ��)b�#�� h��!�`�\���:<�S/��g�b+;��b�0ŷ&"Â�O̅��L﫯��+נ�(��Z���݆jZuv:R���=��:��M��g�� h��4�d=7
^�@���SE�{P�+0���5DJ{*�g���9�uYh�iJ�X>���ݸՀ��	������^�����;5�3��C���Mo���Y_�ޯ[�Ik�w��{��vփdZҧ���i�����!{�L@�rs��K�����2�w) J��3ײfC���/�4\[[�`r��!���by�_��ނ-��: �ұ}Z��\�ux�3�ws�m�]K�5����Ӥ=SM{��zE;iЊr��M��7��w�W^��f,_͹�k����F�ݠ?����Q�|�O��ab�)�?D�R��ۏHz۴EY�l.�"
-���=�ӎ;��o�^���͂@�׹��F��^�Q���#�.z�1U�$nꦜ�[4�2���t4���5�P`[D_���s�b�2d�@��gH��"���c�B(lȗe�*�����ִ���O�9!��4)�sC!sN���K��}�ܹ�T���*�L7�٥b���q���&��s*�+���,A�Ό���������7��?Cw�tt,k�{��9�&��C9B���h	p8�mL<�be��-K���xa�s6Wm-m:��(����<u�@়�{�wpܷ/C�ڲ�]F�q���R���k����.��Җf���!��}�|�#7�5�T�NĎ��$|�B�r�0y�Ӆ����H�x<2��L?֞�ɬ���=��E聝6ţZ{!�9ǉ���(f�DDk+E��&#��s��oi�kU=Ar%�C#��EO;h�M^�J}f.�3:0���9�yz��'so���6@���x�2U��c� W��U��7�b�j��4�2����"�����o/+UD�B<���,F/�zU;%zG���u�S�/�� �:ݤ<���,Mz�l�?qP���8�-r�����u����'%�,��8��@N_v`(�"��m<VyWE{_Z`/4#��[�Q���פֈ�@�G��e���/F���)�E���8��3V@{5(@�[�����T����<��E`�{�/��s�?l�xp�'x?t{�g�e_�5F��{�[��S`�U���I�Q���5�抺Y�K�<�zB�K��|��e��ɪ�NI��$Ҏ-�S��3�hC`T*R���nY���ƴS����W@�����I���6J�Ě�iK�YR���Oi�H4�m5.ﺬ-�l�����R[zc��*&�@�`S6I�H���?D�Ԓ=�mPs�%P�:�}�| 1qq��l:�]�v�s�=�Tv�i��EfE4����-�3�� ����9��3irWdXϟ�ǝ��Y����!��lEbbc7bCG��Y����_1�s��w�/=T�h^��g�ĥ�W�)M_|rf�kv���|d������֑\�K���Q�{LJAZ��n6)�	���C�ު��@�dL���~Eh�m5��-����������r��xJ���$:j# �e�-'E�t�ܧF�z�������J�H�l;�����!v+]�}Y�I�~s+�)|�t����D�x�/i8!=�!�ފ�yv�	b���涑q8֚{W�A�;;�"#�^�]ۀn��b|.�<PuU*�Rթ��zGI����"��$�$t.T9�á�]`6��E�������*�;�|0[�H�s^�{���*�)43^b�c{����|M�uNEN�ha�r ?EtL{L�<�-.`����Ӫj�?�H�%:�f��q�}Y�aCr��~�[Kbx�\�� ���(Dc(�,��Qó�9�Y�9V8��k��ꞟz��[g��x�(Ó�9�bs g�6�[#a��My�z�h���o�d�>�R�6����©=�1
��	�����AQ�� �W����|x�{�?�q,h�a�Ýف/�iC&p���ƣ�����_�n[��� ����� �}b3���X��n������z��v��+���]���C��	{&[q�7��f�ʁ`kp(����mQ�ֻ�3���#�w_,8����|��L��
�~�J����:n�.r���A��Y�y����H��O�Ʋ�3�����Li�^���̶�W�5�Tf��A���	��a��h�Z����o�y�Fe9��~P�׮�	�D>�<���,��Dg��t�6���N��W�(x(�E�'����w�$�H��VTqT���ܽ��i��i�@���K��2ލ�o�^-�����z2:S�?�|�eI��j�<}+�S'j���G��i+'��OG�9Z'�ufC�J6��D�?�Bĵ��`�&�w� 4�z^#�I�ሔ%h����0�0�u*R��t/�wP͚,Nԋ1��� � 
`ܐR���������0~	اK��	�Ҁ��-G�� '�8�L�`)%�c|I���B?ћ��jmߕ�E���bd��=?����ćq"aȞi8���Q�DT�c�l����$�H"���n��<���S�;���H��$u	rά*���㠳�䓫�煽�05�����Ñ��Fͥ��H&��j�L���;vp%!t.��Piy�l�'@�����&�(H����O۫�,J�ShNtr>~�ޑ"�M�Ci�n���p��3�E)-���O��O��I�Û6�p���݆�Ӵ��SYI�|��8��>�8��T�*P�d|)��Y)�(��Dz1�ce�'�i�Ip-�Y羋�5��9ȚM�7���\M6��� ���G���ЮbLUۖ�Pږ#�=���tE��b��8��'Ry=��
���8_���� c���$Bs<M�{�
9���b& �3P9e����W��=ʧ�K���x�Ʋ)U���7������4_��Ȗ���N_����}�[�)㫓��An��PZgR(�<ǳ�%��n �S��V�z[�'r#�1�0��*4l���'߯�s���Aw(�_J�X�Gv��,�\��g�t`���RpuX˅EG�0A��2�^����M�^3:�H�=��=�#�:^O}��7<2In�5���D���;VWm��N���3�9�.>�7I=z��X�n)�
đL0k�>Qݨ��������/����{l�D-Bb��p�_�u���M���0ʠ�X/�l�j�a�����,��.R�xG�:���?�ek� wuf�@�@�JJ��r ̀=x��h��Z+�"���>�`�XuE�)�"�R�ི���".Gނ:�Ai6|b�S�|�Qk�Ɋw�=R��K�K5���k[
Ӥ����9"�Ze~�,4T�����q1P+���2�sB�O���;X=��-OH0�4�?�+�yQ��8��H6R?�� ��`����-��0 �;�Th�Y����9�r&2�Z��䥐��a���M;'���qI
�@<�_����:d�$*J��0�r��I�ͱ��#,}�-�ߜ1PX��VN�9����\���W^ceV�Q�$B��Jb�L�s�ØOQu,b�]t��9�V��%�ne�[���I<IOUn�f`�1�Yb���ķ8z��"�O��1��x��"��Ж�X�(�K]ͬ�o���&mΫ;�(;VF�������P�'���ϭ_A8�L�1>�Y��DF��G/��ގ[��I5��z����Ǐ����Z���[U]���̫�v@?p�e��3�Mn�\ɽi9����_x��X PL�������{1��IE�o{��?��o�Q�Y�g�dw���a�)����l�o|�_1
�O�����|b`�![{�7v}6_���Q�gȓ�DVA��ig��W�j�:��rP~j�g�ěd�{m�L	\�-�xN+E�v�j���z�]b�E���Jį$����ZN"ɴZ(�.�����"Ь��[c�+���y���Q|��k�P���"����v���U�S����َ<x��+j]h|Gb#���=�2���Ӏ�wޮl�����s� ,�B�ͮ���E�d9Jb� P8V|����y�����=H� �U��??T��߃�hr ��[I�����q�]n�s��Ŕ�l�-�T���T�V~f�
��7S5�t�u���VI\�=-�+Bb|Z=������$�G�Q�%"��{�5u�T|��#�Ҁ���5���0�e��Xt�V`磀�ui��� �&|��=�>8���y{5�7#_����M����	㵹�b\�wS�h�0�7�~Wc=WٿIĿ�5[���ă�E�EO2Y($N��`}���^$�)O�@�ޘ��/�ҟ��M1��ܙ���דÏ���l#������$b�n�Op}��x�}�qe؊(}wb��?m���{���3#����,�\1$� =�x��3�D[�lU����6�G |֕����!�`8����1.g��_s�\t��^�fu4|hZʽ�"|;Ĳ����ؚ�b�lbg/����F�g��،�9;a��>���i��'Hc~�֛g�Se2��_,p󺖥A\�A�w�y�r�����j��9�SHx<�a���mOOR<���q�R�B]�g��H@�	&ʉk��B��������"�Œ���%�u�>qNyd9�wk�E��Oh
�8y�͌݉��]|lpUOn?�����H����-���I��d�\��\Z����`��Y�q9E���T��͸��y���ޕY�t"�E���3G���U��ᖰ�P@o��q[��r�D9a=.�f�}v#�f���?�LAb�xup	4HX~d��B��[!FR�r1(zٓ����B�m��
y��i?pa1�Yu;q,�k<Cw�L� H�Q���$�K�%��̡��OW��Y�S��f՗��*(�a]"]���<Н�ׄ]"�]��rG
�rT����Ůq�^����x[�Q\�]2RQ���Կeܥ��%"��>�z�~tؼOۺdǼ�}3Jpژ�Q�[Ju�������=_�}��~1�Z���!Y�w�͘�L�Q�.�O�^��z��d-��g��H��&���BS{Z��b�bC��\�E�f���?i�a�-���j�G��xʴ�8g+���҄�䑉����7[zMU��l�O��{ް�`�+]$��5��F��5y>��X0�X�L#�!w.�O�nf%(<�=$�z[ �Y>�z��k��;A�z�A5�w^QZvV��x�c�9	�_�͈J�-�����-<�ծz �(��f4(�>�x���H�r�?#ߒPҸ�eįޥ�xy�<<�yr�=J�����JN��M.{���[4�dV�G�s�Z0����o�+I{��h�n��Πg_.Z�G�U{P���Z�;���0���(M{9���$\��$�<Vhm$�:dE��ﱩ��ބQS�d�# ��}��%%_��$�\S�z�f�ԍ��_I#\�����P;�L��,�٦v�k�*Zq�����[5��&�3�1=~��U;Cis���eD#��+�]��S,>F�̪��N����k�%Eȣ�!�����:�y�C,b����������׆9����>�mI�75��~�4!	(���!�M2MNݥ����7b]�Q54�˒�\��su��c*Q^���g}�?+�
\c�Ҏ>ј*� �)p����0)`��(6zk����!G]P�����x���ڂ63�]��B&ճ�}8�qw�(�ݍ�峴���ʜ-�4�~��[�7����5�Fܖ��Q � �29)�KSr"M�SX����,��xm]�5���t+�bc��RE�3j^)l�h}�,�5A�z�2���/�������ĺ��v��'ņ>����F()3Ÿ�b�4�W
[��=�N���5�� D1�zS83q��p����V������������ihx��f��:K�>t`�� ��c`�EW_�x�j���4Tplᨹ��:A�p�J��D�q柬SP��������,�q�h
��Q��.�Z^�����la_���P�Tped]���H��ձ�[f�Jr�ŷЍg����m(�߽`�T�CZwt�ژ�ş�����2�3T؅�B�E�0\�ή9�ҘO�vd����M~�ݙ<�,^t��7|V�H���d����?f��k�$��j-.h;/B��8�Y�7G�T�܄���W�>�<��]��z���!�,��C�]�	ءs?��L� dхc�s\	��o6zB^�z�g����-�B�,�6����͙�%����3p?ϱ˙mFv�����v̸ω|���ǃ����]�B�A��Q����
���{w������	Pbi����{$�qRe-U�T{�&���U�3��X�����ۢ7���M�CD��nկ�
*�8�ZsU7� ����T�͛02�4V��l�;��������\� p��T`G�8V�Ԣ0�v� ���HCY=g�"�h�_�t��՚kpt������!�䛚���nE[ߝ'ԋf��+e��A�k����蜤�|/�)�G�h�{�t��w8�鉍SIm��mPsT!��J'����`����AR,��r���U$2�v�`�D���������	T�R+l�,|�w�2w<Rh����U_� �Ԣ��(�=k�^��=syҤ1�<U���H��?�N_�S��0ֆ��pY2���i�1?�7pei�F`*N�d�X�&�]
��T�Cxd�n��A�p���x3#Y�g1����8�abL0 C��F5͜t�NL�FV�\V�DO�>��tl�D���=��V��]��cb�i�]����M#פiW%�>���]LtPbi�v��tA���J�yc���8$T�A�^Cƕ)�����t�������v�馫,K'��)�o��v*��j��0�G�N�c���� >J1/$�f�7n+����o��kn�E�-i�[��>k�M��_�I�A�(�����<q�̂�>>g���y"x�E�<�.X.����SK��闱Ƈxmڮ���,�wQD���`�~��V콟�,#�����JJ�(�Mw#b4���qIN�2ы��q6@і�fYOss��Nm��DJ�	f�=}ʣ�i���T�w��t^��{��'y��w��#9�wd�b�3�wÔ�9���M����9�E��ɿ��-�3�Ϛ{j�����]�����M��o������Wd�?)	f�f��`��Y� �y�����V�C1��	��R!~9Y^i	WJ)m8�M�C#������T]F�S֧���U��U�狀�&5�E����:��K n�0�2��B̬ ���x�{O�P���|�TG��Z�n*q����J{�`P��)
� ��s���;@0� 1Aob�WIPbqr�0 ���^
\Q�q���=�E5�)�x�I�	�-���l�\�� �J���%���vO8�π�X�~k����� ��v̊լ��{�o|�v��sL�]Nyy-�u���+��ɹ�;�~�g��m-��M��3�[���Z<���ܒ Rd6�͇��3=�M[.���-�fUY�@!2���|��0"�[k���&�B*5�7�ɿ�����wk���ؒN�6�c���U���	��[-F�+04�:��QVj�'y��}+�ӈ)�c��x��L��џ�uI�=���4��]�>h$�(˘C��@���5Aqf�������V�e���\l)AX䙭�:)�|ؽ$��$X���<�Pb,L����TW������G~�ݽYxMv2�K�NL�ku�۶�?3v�4%4�47� =���*����*E$�����f�i��>{H�D��F�|U�����NHAwut�sW[�~����o��
.$4!�~B(�m]��N��y��K�]�n���H�O͏��@�1%ʥN�{�X�1�wg�rO��o9 %��S��L��t����:��+H�ƓIcM�����-̟�zp�Kۭ�wDmj>�8\DJ��b���r[B{?����&�}�w���L"S ���v�x��S u����8��Jp�ɦ���{�1��ذHt*��M���8o>�͢g-��i���{���#n�& Yt��V�6l���^�,�V�mԢ AMG�0�9�i0�{�ֻ�5f�N����]N���%���aw���c7�Sy�������l6A�~
��v'+��j[W�%Mb�$����х B��0*D�x�+�]D�ʉ��<\rOC�0��2��>��b�I�2WdM|=�A����^I�)ӏ;�1ms�b٪7�
�c��oY<H�c�cl�k�+�,J
f�L�k��yJ+MĈP}r��I$�/����`R����W�+���v�:>�_}%�c�Q��xP�_���N��#�6b��IO���F�	=;(�-���%E@�}��Q9GNZ������"�â�Ϋ5��_��X�ak�F�6��EWI��e�#A�p��"N9�t��͛G� ��F���8,F�7����Lvo��i��\?��%�U]�����
��P��V8{֡QU����L����v1��;��޷��S]���ފ��}�)up*�x6!AB��^L-8�oS8P�_��7��
ꨍ���L��z��_��+y��}[�#T�v��Z�(@lں�T�<l*��)�Y���RJ��e�JC.�(���"����׎�<e�߰.s歗]��?�q�b��'�<�r�N78+�'U�e땛N0�|_�
��0d-:��@���$�dd�e�A���V���7.��╸+1/�����-���t��_<Y�ъz���Py8t�¥��	d̿���s
�?SS��� gRҾ��ڰG8R��%_��n���O��K�ܫ�agmjU�/�%t{*�W&�%i�;T��}�d�0u�}�@�[�3�z�Q簼�ǽ�P��NɁ��Tmñ�ةG��
`���V#�ϱq�-Hi'x[)ߖ�v)	89l�W�<Yՠ��a¢d��@�ڛ��"XX���.�&�E���Q�ɕ��r�7��8��n��S@ !�!j�j>��%��&�!kP�J���J)�ϊ�-���+�x��}{ ���OJء�tgܐ��@vqmF�%���=�r�xJ�M���p%�M�~�P�]����)�`⤿>��;�P+,53W���m�SX�jMH�$28`_��Bo��pbX��Yr)E�_d��D��/1���ϲFz��+Q�)is�� �x�d���R�1��\��ǵ&Rݐ*�Fa_��$�\#.;�>c����0�h���̭t�8�;�3��ڦ^��l���?8��+�B�X��j������c�$Z<�J�oL�i����r������W�QF�'�������R�)=~�����D�i�Q~��&Aj2Sj_���OZKnc᠈�G,h�9��l��3�G�f���.2�i�}s;� ��?�74���GL�S��A.*��3�-FGR}��|#��=�-S��p��ꏿR��b,rENX�mR �$�R*����|��8�֐p�������O:��L)�$-�?��������n�ϭ�h	��+|5[������ �߈U<���)~�9�f�?7u��k��+��x̦��Т�f'�@R�~,_�����C��L+�Ɂ#1:�����ㅟT��m��'m֎��<��;�oʡ ���GŮ[����p���ΐd~�ÿ��[n��F�]g��[�瘜i8ˢ��Vv�hK�
���4َ�@e8� G>�ȝ���1�Df�5�*-}y������p�y�S�����/9*jiڰY�I��@ �&�H�g�F��^�7g-� vU�˸A��/�B�u\�w�۞��#��	7M9�.B6����[����j��/�r�C]�[CY��%��O؊���Y�f%��P��b��*nN��.BKl��3fY������0^��f�P��t���ߟ3�eC"��G@�����^Y�H�a��ؚ�U�`i��&�a�ˏ2�ښ/�3��T���}����h�����-�b�t�>�}����ס����П�%ۏ��hH��:*T�7�(���ьu��@bX����w���p�b�6 ��r�l �}(IO�9��|���Э�8|��Fp �i��v�u��34s�MZa����y��#xH�������a�S���K�i�V{�aid����Ay���̀�$5'?̧�!+�x	����{`��H���w�C��LIR� ���4�n0�>���r`���_�b8�J8@!<��I�`�wv����)����1��].��5��4�Mu�ό��t� xOma�갆�ʶ�&�l�"5�9�5���Wa�P��ݝ�c����b�dNs��l�wPe�F��S6��X{�H-���C��I'$��I"k���.k @$�s.3.��4�4�N��/�����#s�$М��`]E�NG��ϗgS(��5��&�+Fl����������
�eуj��-�!�;~$�3��S�OC`ʈ�1������ze��.�h�렆 b?�CX<3���mR?iJѵ�SoG�TQ&R�8�e��J˥/�5(��4ԧ����̎�Fg�[��uw�?���߆��C�<fvv��A�p�`4��q&c��ބ��hM
��	�0X�䒩�����ՌfC)Qk�o/*Y����3����3�u%����>L�6])�ǘF=�uhD�D�߾D[�`R��Ѭ�rX�Β����te�ʘ�0iZ 6+�J:ʻ9Ҙ3�T��W�\U���p�Lӱ��#n���Eua3�����WVǑ8���Jn�G[ׅ���a�A���sA���֠{&P�"{�G|���1�j�8�����������վƉh)Lː� ��F���I�(��>5��<(�������{�O)*�"\e��e��~��oX��q��_u^�0���mPdCË��\�}��X�d�>\Qs�����QDx��3���0#���i������޲���\��Ks���0�����������~Cǲ�q����V��\mz��P��~+�.s��hQqa�f������yW�3Tₒgn�`U��5.�;.�X����PΚMA;X��P����?_��Ú2%��m�ގ�������ժ��Bd����)��T=�Y-Z���uBۀ�3����D5\�O�*'�ɺ�^M\�*�<�R��ﻌ�-��Bm�}N�m,��@����t �I�c�>_<�
7�����+ܢp���Ν�AW�RL�ܤwNR�Q]]\��5P�p/�ɗ�]vf�i�	����](�9V��8�z ���Űf�")R�5�g?��?xb��z��l��b0��Ug�*�.mL�׵7����@&�nZ����Z���˽�6�מ���X��*bEs��O;�uj�eL=q�`֥�1�󤖳TڽBq��P��ங��,d{u�n46"�UpDiIz��  ��꟟���i���RL�Tם*�j�0^����a5�vU�|��J]��/����P�K��Ik�J���Lb�>)8bYo苏) l�Y��qyG��P/�ŗd��U5|���p����XwMC�������K�36>\V�5�K�-�أ��C���)C�]~	��[�����=��60�I"��F��L�	 ��7�%4�*ɼ�J�y|���o���]��Oy|p�S^���8z]��;�д��������;�dZ>��kg����iƖ5Ge�n�q����/^lb[UTXQBWr�U�k��B��-7�,+N�z�y0���HkC������6Ԗ���?�c_���4�B�"��NR���±��"��^e6������HTO��ɿ�]�m�-o�s]��2 ��A���7TE/����:a�sz��䗁�bv�����)+s1��M��/���v�]	���o�3때r}Hp��<������"����p��D6:V�l��Ʊn&�V�b6�0r� ܅I��H~�__i��,T�Q_����O�ʢ��*^nO{=����,v<�kTT�q����������Ƨ�d�ɓ F?�����-�$P���9N~��OG���f�~�Zd�j�ep��M5��*����s�	��Z�H<�n֛�Ri� �\�*D/�kR���p.r��~`�IE�Ѧ,��fqI������K���S
���8��<w5�}C���#�Ɓh��m�դ&'�l����jD�L{��y��!�@[?�56�<�H���Nw�(�x��:!�=�
]�
o\��wJ��<���Բ��;�fWX�G�̩�w7����\=�� 2��V��3�`�\�}G����!�5�j��'�L~|(�iYۗ{q����D��k݈�t)���R�� /f>,N��1�m�B���[�v!��訤%�0�%B#��P*�E�J3�����;�l�r���1݅oke�M��QT:��k��g�J
/	|�AS�fl��9aoE�[��f����t2�%��B.�zS�*h��1�Q*Eq}M(l�� t�����t�#wg��Ȑ�"� ��`��膕��P}��+6[+��>B0sBX�d/�`1��r&E��f��
�i-����W�,{<BuvD��s9��N��
u�}|溎��>���ۘ��{ퟴ(����tV�@A,4�eTr>ǖX5��G�
g�@������f�.E�g�. /0�[����ej�k� #�TT��N7��&i닩�'7 ��J��x��*2.����H�D�u9#���Z��c6�"wn&Mᣲ�����G?;k��Zc@��f��"P*�[�ï�=5!	��L��m�\�wVd;�v�r,��[�&���/�Jy���]gh.�'�p�fй��ɲ�2o�A����V��z&B���X�>8�'#��!7��C�2�z]	��v�����x����.6/�m-��5 ��v�7+aŴ�LŮXO����<`>t����}ZyS��eX@�:�Kc
�.���N�G�Ak���U)�rơf
�ʹSQ��e�B��}B��e?ǫD�,N�S�r�I`u��DI�	�G`���]hRƭ�-�6;m@v�?+��>��d�0/QhT֮%�N_=Y9#�:�u�����/Ce鎔,2�Q�Y�
�txFҳn{B��AV�0�񚭙�<��T*�)��>Z�?%T���Zԡ66�R&�pAu��%ǽ:���@�3Znxֳ�6?���@�fA���y
r�`���~��NWR1���=zE��r��-v��9�.-�ܲ���.q���k��XD���<�
��ͺ��BeIώD9w�3|�<����ӭÉ��Q��}&�s.SC�&���p�#�H�;���  FK��o���n�Y������dZ��b�S1Z��G�����N�Z��FS׺�
>kd �.��a��*�g{�V�5����v��fSy8|&?<`BT����5� �5$�3�'�܅Ν��,���3�-�t�he����G2%.��0��,�'Ln�΋���u;���<R�YRb��Ƈ��m;�4DQ w(\�M��z��_����A�5*6z�d�B��	�+�Qhm&H�J��!E��=� X��L�@%UFs)FsF�0�
K�����q&
���T���-tX`1�Ae9E��#�s3�i^vz� 'Ĉ�z/��+6�bmt�[�I��h���]~�<c�Bs=��{E��R��]��p�ۢ�;VU�|;�uW�	 �
'�DV��a�qẩaz�/L�YEֳm�b� Q��&��܀��6:NK�H��l�Q',2��yOҘ��|��^��xPq�:Y=́����"䁸5II�iS?o}���e.��І��k=����.�a�=��̮Kػ5�M�ʬ�ݍ+�ʋ
�j�q��hg����1�o&}��&0N�%��}����|y1��ё���ge�T�ui��6<ںNa�ɦ�J�!�a�e�3T������*�ĝˣq��4���Ў�����T�k%�7`�,�b�Ǐ
j��}u���$~���A�we沤p�I��r/����	3�ψ�VTŤ�U�D�5����D%�Ѧ;���:�Q��h��qO�Ŧ����ߵe�p�]�-��`���Ҡ3 @�}[����5E�A�S��D��v��+3�$e��,g�!{ɮ����;�xP$#���V�)����)��{�)8��Ӛ�w�6>t�<��|�;�����UTɨZ��j6G��Ɉ�QSa˥D�w"���^7�pŁ[�1!:������sP驻X,]O[�^gGmE"۽Ҧ�r&7ٲBTIhh��t��uV|?��znC������[@�����Y),m���'	�R�%�=</���a{iR�yU�H��&#Ɛj�]?j,c��L�R��o���M����&�I-(�NZ��)'��tKOT���kǢ�f?�s�y"_o^]|�8ɤ(�l� ���ص�_B���2�o�h����\
�Q��	�T�hwx��0�]�A �'#����$���=��Eֈ�W��؏�fl���e�/R�q&��l�"s MpKd��?B��4�!Z+ܻhܟOk�"��H
�69�j�o�.�?�?�Gp� �Reg�`v�>kdg@�{��Sa�{�4�fľ䔋Z���x9�`�J~����i&;X0�u�5��܂�O99�ee�0t�,��!5lx�}7�TI���s����{�zv"%8�9��w�n�E���H�qSp�8T�O�s�+� X�I�#��Q�B��W���iP^��>�����e"��T�V��!��0�n��p�/���4���J��Y��Q�j��6�r�E��y@�.�Po�m8��S�x�ͦ�!j�k�K����:r�x���5���v�,r?>�AV3)R�����b�P��S�e�|��߱d$�
x��-p?�q1�~��������v��!�����!�?^�ƭ<�%�SW<�퓜F
o�_�"j���Y �԰�{�L<E�ad;,��s�$ϩ��i,���ZU�w�i��>6�Ȑ�������7VrV�'"���m�e;r�	�Kڊo[;����<���<�	�gܷ�Zo6@ȞH�5!��[��;�L!6�hi��hL͌�a���Ý�0�Z4� b�����'��P�'{�B���1�^jn|��O;��R�f�����ַd�U"\�.G�ݲ!zX���pSc�W�C��S�b��	?>�!U#7b�m���܈�a�״f�r"i��U�R^�v]P	/PB�,.�7X8�������IJ���8v�u�m����vu�.A>�������j�a�㢄�	������dF��lp�@�D��k��p/Q&tk�Tn�N��^�X�t	��w�=��Ħ��yts�ϑNtjQS(�]N\ή�G˘�CBm�����"z=�a��iḻ����$z�0��D
��yj�5Qԙv}�ag�kRyj�\g�` mn`H@���X��`�"m����z�����r?M��������=45���#.���<����d=Mw�CȠ�ċk�,+y�����b��������Om��G���m�1^Yq�� dۈ�1��\)9��2��!�&������ ;�Ǿ�|���Ƈ������\ձW���a�w��%�u fnL���v�"�/�A��c4��P�6ʱ��X�z��_}�Y���C%椆+T�q�_mqgf^�Z�T��N�u��O><�� e0hrAAP�$[�H���=I:n{J�wä��ƨ0��H|$-���w��]�#+���+f��|�'��)6C�m6�F,�f���M��)��< Ǻ�h+�.����<�s�gC,W�3ك�N$6LLL�a�=�"b��l7��q�LA1_7��g,��P��kz�U�H�mU���Vht��K{���.*�N�8�T�A?@}Z����75�%�˿��w���^�s���ɛאK�N�@`�H�"(Y�a���!���еQ��$$�B��!�-/w�xM)��uw�[T��6C���gҘp^;%m �Al'��̞=f��p�C�X������}�QuV����v�[l�gFz������h����`�H��v�øOh^��#�b#W���fkr�������)�]��.ʖC�e�QRG��nU�v"�jT�(,Ԭ�\ʼ�� 8��ި:qM�n�u2� �Hs]*�gF��Xj���xW�ǑW���F{�:k�(+��W���+J5-�
\E���SnԪy������Ĉ�f]2���Cx���0;�?����sBy�T+'	��o]��;��A�dߓ�h��c@�O�F��.,�����	�������*��cd9�!��ލ��@?��`��Ϙ>,�ķ��^۪��M��2P$F�Rx���*���O��L�5��Ķ�u�xf���2>�K�sde���\"�/�[(v��	G�#@'biS�+Ǹ6����Ol����RY��j0-�՗����gExj�������֩����Td�)$��N�|�AW|�w��N]�w�|\@P�a�Q��ļ�C�U�b'w�g's��7D@���H�!��3���ok�`Ъ�|4�k��:�������2'��ްU�P*)���N=uF-U���j�PhD㲼˓H�\�x�B������b�^�$�$+�����Oa0F_P*�@'?�OɃ5e$HI��}t,�z�BK�r����:�nĕ��K僤G�I��r��[��[�M�P��'��v�{�ԇ�f����[�$��/�W� ]\��{*�����M%�����+�c�ȿ�x4Y�K���C�p�cC&������܉�0hXD����D5�βT��l|��i�!uQM�ߡ%�	7��"��N�0���������4*�Z���hR5�ChH�g����:\��疞�|�fN�I��n3�u�uؾ���f�O���W����Z���3��gUFo"<�Ux��?*�Ղw�<�>0��yqoěuG����E$���2ݣ�I� M����E��Snc撴���M翱k��hZ��X��3ɺ"��9��qN� ���,�KD��gnZ0��M�4��II?�b 'T�D�؃�PM$����XZ���d	���Ĵƶ�������A|�u.�}'��01db�-�䀕��!�V�
A�_�;J�e��a�	(��"ϓ1�'�̟��J��yVm�X�(��%����3bX~}}�2l�V���T��k��!%����m�����F.Q�%c�� չ1$�'���L� 8�+ݍ?��囂 �!Y��CnD��2�l���T1�W��NkY��~��������gÇOP�ssN؏S�m�6�W���х�Mr�r8FY��߆k��2W坦Y��ت��p����Ռ&'>�{�	�ֳ{GEP΍�RLJW�:�k��J��<;b���Y�;~օ,w`��������\7�
��L�b�-:W8u��>/O9���jŏ�)L"&Š<�Zm~��[�I�TK_��N��TGg��u ��|Rc�Ҕ:�O�o����_�8Y7��w�[��:u�.�伡6�Pp̄�@tS[-�-$cH�@;a�'0d�g�g1_�	�`��M-M?s���/��҇�D~܈S�"`�����b�3�m���N��A�������>�첵@/Ux~�f=E��A������ 9tq]:-
4,n\L5��
�K����!��َ0�9�P���[�H�Ў�~�3W39Q���b]3]��k̪-I���ځ�&��
FH�������Ұ���2��q�_�E�O��5�^�E�a��y��42�d�e�Lw1;����:^ݰ^�k��%�w�����i$�3���/����g���7',�*;s%���#)�9��Y���Xq��\@U�|�0�K8d�6ݔ��f���r)��=m��g���\V��0Y�8aa��~̉�����AV�����r�ڤ���<ʋ�"H��M�z�P7�ru�������@�Y��z6��f�7��h���K�C �C;��2w&xM��.����WŁ^on�i�֏�-�����:U?�cb�s��<j�vs�dZs _`�M�Xq���Y�>�或J^��(�;mB
�	�g�:9D��O�ʍ@P��^�ﭛ�n2Z�����2z}��L����IK�4F���RQ`��-N;�i1�W�"�ˮ�fCP�{r�\>ry�$o��jS��k����
�?��tyt �ev�d�4�U`��p%i�>�>��Ӎ��<��M�8���iUV��_����T͠Y��6-������g�HQ~���hpR�B��"4�P)0�i�m�!���P'x�����BDM׆R��b��}�������� �X�op��#@�l��J��<�͵V&e�.�Q�h:������h�fVcg#��Y��#s'^���^:[3�.�>�����_�Ԕa#h�}Δ�!0H3g}Eu&~��PZ�FI�nZz�`��'R�p���|�6�a'��&�v����2�װh��D{7?6(�6	�_򧆕Cܳ��k����59m�qJ�U[��(��:����F�VvI��5g	��K�3��K���ې�1>��"!��:�[�A��FɄ�*wa�*���ؒ��ʶp}"4��_�t�."��clNHD����j�W��6bB�?�<�"��@�� �C���V�l,/��Nýu��;��A\(�R�х���G!b��uG�m���g<����fQ����5Q����tg=��>`1睜���� 2&bGґ�FD~�"(2){���l0���M>p	�k�j��!���:�cӖ��������
�L���'�Z����}���|�e	�M�b�;m���~��{2	@����ǰ-m�����
J�u��n-s|t��»�����a}8d*�Q[�u��z#���*�TD�8���%҇�mƱ.���Y�<��?C'�P�No�WM�v+��	�,|��	~�(&!����J=	h��[9��_����D��T�P���a�ٺ�b59<��ǭ�*���T��k��lD0��1��������d������ W�d���B2S�]V��3��L@U��H.p���8���^�O���|O���c�����VbФ-�+y ?S��Z�&�PM0[��9�Čk� 뛾\��8�|�Z<��ў��� j��~�NTjeD{��.��ș�Ŝ�7��	��o�?؇Ou�A}�ݯ�� w����p�Y���M�
7�h�f~|��̂W��ǌ��tR�c�V0�a�7�F�|�/+��&�J+Փ=���`��6R:7�Юd�:���{�����T��h�S���K����Im�}ci��{F��B�bo�F�ܟF�	>l�`˭E�ST�vJ��UMk�dL�H!�In�¡Z8J^נB9����d� &�HD<�SSb|/�[)���b&�'�֯xZ��Z�aR� �j�eEDF����U_(K�<zD
�g� �$e���!Sa�@UR����M0��Y��R ��V�W-�(xo�3!����(��䴒������b,��P��U�R7�l<��z5�Q0ԯ{�<Ș_��k�o; `���xG�w~�D^���� �I@kbnL=�(��"t��݋�(3�DZ.�)�6$��M��cp��gXa�O!v���["�ͫ2@E�N���ڝ�)�QG�榩bD�z����;8xm�Cm��ퟑN?2`}�qͿ�F/2�똚�e��Y�L�k���Ɩ��V�p��$.Vry�:�<�h�m� e�L����M�Ǔ��u�I_FM �?����ީ,���E��p�K����oŃ�T��� @�UB����&��V#�:g5?oB;���e5�N*x
m}I�GTCc�9���~�����e��3�1l���~���<M�h��ٓ9��S&�IA)ͩ�(g��Ϣ��SU���c)�"Ii����h�8x�/�LlM�ŇBp�;+O�T>�̱��4:{�^k��j �435ϴ	\��!o5�w��}{6撶fn����6O��2��[y�z����g�*��|_I˕�/�i�lO|'Lc$J�N��vܖ�e�� ��@�j�,c+����Rդ
�]�c�Y����+��+���:��Q|������H�k���BMN~?\�s�^�i#C��P�%�A��4'!+r^�x��xˏ�<�,��}�ߛN����g)��v9��N�|@g�p�Rt����Pi�h8r���3B�*�er�.�g��������s�E��*���Dm#Ƨj� ����}ZuY�t̂�ɂ�߅������d�U?o%���6(bڎ�7`zn���d�5�AT���Q��i��zj�J�1����щ��A�6�b9^�	����u��&�Њ�r�����4���+T��Qg�q! �.��.'��&�c^�Cۀd�=���
���SI]��XD�~(���^bw!p��Ӭ�kZ�����U?���J�k	��vJ�hWv�0��J���o��?��T�{�����u`��q�h+$˳��5�)��XX�5�Qt�Ws¶V	��,5�
R���D���!3([��K�/۷���iU�l�]�H��^��M1�[0ޅ��L�ÂFP��*�AD^�����
�]�#8�Rɝ�}yA��)a�B��;k��ݎ?1M�0K;�D/��>��O�a�}Q o��^aМ%�����UAj�]ä:�R�p�fv\S��?�L� 2�����da7o�|>K�j&}Z�%�j]h���y@м�����Z��ɧcoSR�a����̂��Rڽ����j���ƛA �v����)~�[pV�G�ֲf�6�,�����Y��=�{Z�"D�5�^�"�;�y�zq�O�ܡ�.�D��MG}߮���)F�B	=Dn9z�F�Y�r���>T�F`�������J���+�� �I�!��ahj�F�f�᧜~��Yj�D��rg�iZQ�f���uQc����9S��m�'��[�B��/Q$�� �+�W�;���!�����s�I���T�P��H;��-ؽ�Dv+K0��3��L���˩������G��ػ�|��L�"��	�f��CVrS*,��B���[�xurG����߁4�X�z�b��(7�$�\5�q�Mʶ�h��iX>�|�4/�g�oB؍ŅZ�ޤEm�R
^lH��A�����Z�S��{��@�xl�[/5��00��v�@�Y�`L��\��Y_]�pދ�)��~�/���ˮ��
��U�\���wYWG,��JHg������v9�tTV��V�-+����O�S���(FE��qoރ V�¥�v�HUkP��'m?L���?�py��5'E(L�R65��D��G�P^2�6���B��{rr�H�;{�]����4�'�nrRG��Oi~aS�O��Ow�E���'
1�S�=�N�P�!�V)*B���f��*�#�`HM�~x����cf�:D�WV���<.1�:��}�À�}&:cˇ^N���A�iH����l�aNK��%�6T|�3���W9�:7;�J�j��P) d�9ٞ��������Q���r}N�6��U�ngF�Τr*�)�E�`�B�"�x���uK�,Pi*�彜���3�G�4,S��)�#���҂��l��<�E���<�õ������^ߙB����b#Q��P ?�p���'���䧙�"�����vK�S_�O��=L]����!�^���1��,
T�%�6�ɟ�v�!SR�Lŭ��� s����@����|p%�"����9���<ΨVZ\�v���sgZ�z�8����	@��k�%�a���mt�?���%2�jS�bnq��k������s�mL*j�2��I�lc�P�����������9�JH4�kq4 ٟ��S�	M�fl�����K�=G\r����T���NM�F�P�����92�eu���q�/5��&Z�K�W<$���=�f��kD١b	ׁ@���!������N��@нI}�#��'�τ[�e�͊���<Q��
�Y{;P��{�+l�C�:���`"��6n�����G��%���ɤ�n�8X����E����K�w�a:{
�߱v�E T�plN[��b�ힲ�8U��:;lD��[�&���J-Tn'K���^l�_v2�2O>���(�gQ�XPA� H���V�'��$��je�	�
*Å3�)�9��<Hrk��|�m/ .B��c�6���Ne���`�ѝ�y���<��E��x��}�'o���{d6㤷V�sznlL�L��Y�׷6�c��mH_��)�?�>0pЫ.܌�텻��z��n(��ƨ<w����h�d��66��鸥e�A=>)�ӆ`�����j���P$�B�$��_�
�-ٲ��B�%��$�����$�9�*�Q���;IϐD&-o��J�:���c��T�������[���%2��}��|�"� 3+v]��Ko��w%�7��L��Mu���n�`w&���&#7 ���w��q6��1�>�>���G�rU^D'��8����D��#'�W7Gx�jϧ����Z>��;�ySA��C
��><�<vi�gh�$�\g���T5(5�o��|�'N�
pDm�;;D�[�q�/[Q1Mf��l;GL�H���).yw{4�Q���/��H+`RH"�b��gmk��s13�`ci5��U(�·*M�����*0��C�Zx�Xշ�L?���cl3'�H�OX���DR�<��?�}-B�+�Q?%U�~�{�����4�9��'D�i�N���Ђ�oG�h'mW���2�F�D���>��oM}VY"�a�u,��$�3�X�����~������*��_(�E�Z�e51����끓��iiv��ΩF�Ep�?������"�Vh�z���׎O�/M*�am���K��6��&��8	2g��Ed+��Ϩ�lքn���h�/�G�F<ɐ kf��a�8[�x�(r�\޻��z�0>�1Y���CŜw?��{�ؘZ��?d�E)�s�N4�+�D��7��fgk?Ε�w��~+�B�拂�R��ߴ*����� G�q�Q��O���P�|v~��"�7�Q�/J����*g4�{v.����i������d�������A�p��+B��E�l�jS?��;�[pV�,�/x�U���
u,�Y�.�%?�ʄ5HC\A� -�U�Y�Op6 �_5U�Y�!o�$�{�%�"jȘ��i޲�4#���B�$�@A���=�l-be��;��k��ȣt��|�O��r��FeK�2��?,n���}S#$�9��j\��&B\�/��R�m�/�R��%�mtb\:�M�m�j�W�HV7�
c�y7ĕ$2���Ua����װ�:h� �fⲲV��א���L�x� ����ƥ�P�������B�qE_��V�\���t_J��vŧ0��Ѿ�i?x��z*hoa���1���5Rt���g�����ge�����ljJ��m��<̬�����o�N����.�����o��X�#9k�j,�)�E����u�K�Q
.�䒪�����>-뼠	�=��Lu�b�z�5��_蕟=���ŷ[m*^��XU��O(p��-����]C�Y7S0�-����#��)�X		=�D�.�g�e(�W����@�҈�;I�$ې��3��j<����`r*���/_�N���l*�E��b���z�қ9g����z|f����Z?�P�)|HX��7��wi�o��D��S)O��<�Μ���ƾ݈�|U�i��u g�ft��.�w<Cp�8�,�����Y���1��#�@�&�3~���$(���9������ �� �Ȅe�֗Z���/4#��.���Hb��L�����ү�3n��r�J�]�����D��=�X�-J��zb�� ���@`�>E_�<ɷĩ��H"�Y��i�\�>9/�[@T�k7q����]�6���OȞ�Z�9���3�3��I~NOf֬�p�j}$��<X�!�p._:ߪ�|P��0e�V"�����9w���՚#��Q1����b�:"+�(|s��j��ͻ�� �XwU�CL��"j��:|��v�c�zЧ����W�"��s�,5�%;C�U{�ㅴ?@�a?�X�}���f�{��y¥Ί4���b|]�.:�����>�9������m� rF�ޤɧ�N�T��4zܘj�@��Q��sE��4�(-R���q�����r =�sd��zE�z:R��#�� �r��s(H���Pa�H���0j���N6
'��*Ql?����\��~5�����>��;4�ڌ�j.�|P1�F�LHv�g��K� �-���~s�яڛ�3�C�H�-4k�7���Ջ�ì9UPYL����(��K������ `d�?��ڧ��ޓ3T� 9]���j���t�c�w#{`��`h�9X����P���Y�2�u�	ҟ_k��G݅���b������!&^������8)Lw�����߲,�Q5�:J]M$�1�nŎ�s���zB��H����?B�z�dϞ�� Xi�u�v�(�.����t:2)��֤'���>��)K4Mr�S��g1~��[��$�w�=�㽙ɄX�M�:�if<�K;��7<�����Z{o���R��dn�(�`�+�
���o ��௡�V���#PNu�E�/�������u���b�^��S?��>E�P�}V;D�b�1��6�����z,��H��&�=�ۮ0��Yh�{`�r��҅N��j� �
c�~����*ؒ�{ϝ�>Zj�1���#�qⅫK�g�Dz�݋���
�"�it�+i9���C٭mh���A�|�����\����IQ�gU�K���R����
�
w�%B���B��;n����v�c�Y��Y��Y c���5���Ѽ��o$7��3�(�oB�w���}��4*�M'�>3/S����lO�b|� c�"�?XS�e���'2T��p6b��0�A�"����oI[wٱ�v�I�ź.z�] �����<I%��������cYw.R�W����D~w"�ol��+:|7׊	!�O9�ngC���C��V���1e�6i��?a�3�8�żm ޱ}�J���������2������ǈ�e��j��ч2dk]�Ɇ5�$~8�"�� H��b�8WX�����&N3��n��sú�+ڠ?ђxR�B�M��E���5ۻGu�`��7��I:"F�H'�r��e���r��U���2����N;A��r��#�k��LSHP���#ƽ�/F�ɦ�9�����q��3j���r��=���A�kX]�i�UMȆ�RPb��/L<�5�8��)P�ZB�-w��ݺ�[k�����/�6-�#�����??	�o�M�.γ�#�dWX�^�]#� >�4x�C3�`��
�w�h�.��d5��T��4�E�aQ�'lE��_�����M_/ٜ�mA������J���Ը� �ư]����6�bWk�����/.�i����Xrl(K��8���3^�GN�]\��Y�O���4P����� �dC�'U��.�u�:��.D��?-
)6k:���nA��U����6<uAFc�;"�1[�2w�\��j��߀�7j��F�%a�1v!3��v(�0�E:#�z)����2_#�n�J��'��p��k��]_!�hlՐWe_8F,��z0��ﶾψ�����+,�)ݭ��Gcz������Ѥm���B��Q�;"�\/�#�g�o$֜���>��E�����Rq}蝡'P+T�-W!�D���e�7�]/�yj���K:�Pͻ�
��� ɢ�#VH�:��m������ni���!=�N1/ZX�i�ߣ���`V�K����s1@����x�����
��M��f��L˗��}$lCAՑ�v� �B{3�)�o1��P� ��`@�P����3�&�g���p2�Jc��:���~�ev���̄1� �sT�Aڡ�¼eI��	�o����S���נ���CVۂ��[bF���k2?��-)Xt��?��;;e<�Ϡ�Q9�у�KOt��R��P�m?z�X%���a4@�N�v��\�C�A����盙��.+Y��/|s��Hɻ6��Qw����T��Tba�W�D5F����������^h-	�h[KQ>�	�qf�&p"�:�Z?v!�|�B"��a'C�E����[��=TRg��M�Y��k�?L��L9ܙ#ڰp��+�K�0Rں�Y�S+��ik��ip�r�'(Wdߺy,�-c��Lp~��p�V��/u�P�q��a����wh!��W��b�W��+c4�Qny��G	�e�QÎ�'��t�9���f	YQ>[o��?�G���N�A�ʐ^-+���}ǎls!����A��.��b��X��zc+D��N�����T���FQ� K05��ƅ���Z��̺�axh�F�W��8�o�O�%�PT�y�������;���W����lk��3x*�iq	;���[B�>Ӭ�J'�DJ�t�O�$7��l,o�?�pO�}�
X�.��ơ���iV#�cO�:K�$��AX6t�\k܏��aY=ݕ䕦��؀��� ��8���N��"�2��=��Y��O�!`�{�D�����<#�.����dJ5��.����*�RG�K�M8�TI��r͏))�O��n����U���JU5(�X�<�P�[�����R�Q3^y��>=K��H��:�(y ��IAA"��Q.i�Y&O�� �>Dm.j�#�8?��Ω�ٵ���B�s� *�Y}ߛ*����\ �� �K�=�<��� ����8��~��������NgU�������n���9�d��A��F�뎆�۫�s�x�Z�U�ٹ��pN:9.Ăi
K�@�Ǒ��ZUmp6?ww��s�Kz4����K�=�*%kP�?�DXG�?N�&�����(A���@l@�Ʃb1&$zM��(�Nau���Ov���]���AB�P����}���T�֯�����#l�r��m���)��*4�;����Mp�w�%\�[6����Z:m'�Ȱ��
��@���"i]$G+r���\��2����.��{� ����%�*�,\t� W�e˫�C��ua�c(�YN�^í�`����'����"o44����6VP���#�4�fav��i�������S>]=�����N:~p�{sH�9SCA�\-j���	�9�����d7�Q�����.�=R���!
�P� �[�b�HA����C��89��F�����♪�������+�yp4����{�#E����m����x��0笱+�׃:8Z}��`��|�?�pX$�;�,QE�Kņ}� ��=�+�Z{J�S�,�N�--������.�R���SS�~����w�df]���>"��	S�O^z��Li��]Q�$��6��^��5C�Ƃ`D�M����]x�6#����C1�dE$��0��+�̩�-/0���-�Qe�3Ϛ�r�1_y��
���1���j�43����玲��e<lQ���9Zu���Gn����Q�N��K\�w(S��7��� ��(�q#o������z�K��;GB�RJ��/P��^Xs�B���9���l����x��lo(��e��K���=��=ә�V#U�qe�-���� \�y1�4�z&����0��p������ Z�c�Ĩ���PO�T���.�1N����`�n��h'=���J�C�V}Hy��U��r^S*��ә�2XMZs����'�,NB5+'�3#��p��k�J����l:2y1�v�W��;���$D�M���,�Y�e���Q1*5jfZ�v��5���w�E���ҩ�C�f��|\�6��C�mS��|�k~>�i����y|�CBW:3O��9�U��!��
#��ç�&�B	I�w��ר)n��1��m�r�ϙq�p�/�ԁ�Sd�78+D�{2�п�C��$�Pά��7��k��{�F���i���������E
˦Z�˨�0:&��=Dly��NSA��U��j�YC�25g�G>V�|s#[H�Nf�L�\%-����23l7U7��ݢ�v�}Y;�8�|m��6�&���w?wJ4VÙiB%q$���u��aM��O�A�eW��o�(����M�X�mf���?p_�Ԭ#f=?��L�K��2�A�Ԟ��AO�@�JS����o�Z[T��F�F��ɻ�4����G��A�yH��NԳ��dZ2��c���Kؠ���S��F�,��
�yäo�1SZM�uc�6f��n�����9��9"���<M8	��h��%�~�������ݻ�r
��Q*,�G�� &{���@��C��<F�Z�:-�o��?:��5�S<��_t��}S���ϔ*aw5�]��Ky��#�CZ�aф��p㈄A^}���y�Ԩ��i�+�С�);�ǫ�) �7/l"O,�B�S#����nȢ��j�<��Z^ֿ��b�0+LV��C}�G܏
�gb}�q)�BN��W�@����d?�� %	@ct�R榰�'?FE������1���H�`h?�s�9K�Eğ��Ћ�G��q�����-�@���c���PW�#ѱ5ma�y^M!�&�o�:!/lK��d�
�� �"��/��,��v�1{+���*�*�s�y�A���Fs4y�(�\��3h]8�X	�s���^bmu/�J	��dc6Ռ7jW�5���Dgs�����#D�ҜHM$[ʧ�7��UOs%���)g���$N2[��l��(R��گ���T��
r��$f6�Y�%r����"~��4�O�(7՚��)�w�i��o��I`"��ʣ<�1^	.��S�:�Ve�;���= ��a�̵`i���ڀ���J��C�]8�5''@A��N{z8���qcP��e�Ŗ���l�=.�܍x����W�m,�v�������Y�g!�mx�¯�)15[z���fr���%�)ܱ� �	(��Ż�\���=7\C|��a��H��d6}7F.�]ט��ޤ'��䢞r�&Z_ pJ��ǒ/K5�2��b\�*
B�S����<Q�2���
T��٪�N��)k�)���A�������K�tI9���~���� �qv k#��rO`��ƴ�����Ф����O55(8�@i�a*��I�DCF�	s;�¤a��p e�&t1.|yq�݀C#�cx�P��a-�������r��8��ط�`�Ӱ�������"E�$R�zs��f�Q<�s�iD���b�h��9�]M�(àD� ��6�����%����Q_�!���&�#l2?�Wn�RUn+��5�OΨg�>&�)�O�Oa��������DU�  ff#۶3�L�Wi�l]b�[)N�R+�Z�9��
�v��Y�S��?}�g�E���$�.�� �XMN5{���	��O�m�h^���A��gU��|�}�O_�����O�)���gn8��`�BP�ɤ���������������X���#k
뗷g�q��75��z�z�*J��e�m���4�EzG�*L�;l��>��1ٸ�}��0a��X�Q��C�>��E=琹�����&>r�f<���%&5�A*)T�������.����v��n/XEi?�zmKdgc�`��k�;�����<�̐PҜF�nr��K{�I|k�/J����g�5���u6s�A�g������i��ZoÙz(��-B�Ņ=ϑ>?Q�Х,�q���k:��Hhj����w�Ɨ���^.��Z��tE�s�]�E	��oux-^��oCZ��Ӆ��Zs ���<+��7��	.>v(�cQ�_ct��� �K@E�@�to�۲�)�u�v�J�<���E.?c].�Y��������s�[Pt��m��B�,�k�u�"��1~��S�>�WSn�#Zm���)��š�\����oC�ML�&��כ¾��\{)\��rŒ�Z��Y��Zzp�*H��>��F�$AM*N?��<D|��G3?]���J9�8��0�5��6L}�!<ӯwOh�^P�e�����> �����F���!��`#�\��5��}�ˣ62�sD���3��
a�A�_ �p���=֗vT�����5"���I������V��P�@�s�eN�*�&�h�TE��Ž��Z-����7ü���:Jv ê����g�i@̀Sz�ٚo&�GYD&4{�<��Vs�a�����!�boI{Gg� ��"vp����K���� ��KYb��p���ߦ��
�5�/��T0I�8n�=��K�y��C�1��b���VF�<���U��EN��S��B6{���){WD��7:G�ݢ���-0`�m~GK�/�٘D4/�fz��3�N�ze�8N>�:нZ̷���h�#�mb�`#�^���̝&��6O�d"b�^[�K���Ȍt��	EIl�&���$�����_9s0 ��0�#a&NZѿba�i `ɤ��	Ά?/��w��U�/8��W_y���EQ����S��?-��(��)Իw�]C�x[�؎��jv�*�gudCsҫ=1�ػT��i�S�"+�ի��l7ӠqU"r��9�=���Fy�s!kv����꾎��#ǖV�#��xl�V���ɤ���՝����v;�g(l&����fT�k�	�����;m�O/��=	�%�����H��q&��Z��/	�<�$��-/m�?�E�"����`>o��n�6�qM��]#u��O���j��X[=���,C4�c�r�o�yz��K�� +*�!_[`����l����
�P�*��()Y�,@h.����J��ݑ����F���BU�`R�S"Vcx����
��pڽQ\��l9R�<��J��u���H#�򣇖M���"�a��P|�K��{9�������PT¿�黚��iޝ��c��y&Q��,ʟ�A�)���t�:L�ZѺ)���(�OE�82O\��|£��n�0����� �y�>H�<U�S�YC���/о�j�Z�R�G��*��rt�1��Y�5J���cH�ly�?����{���y�֦F�ߓ�����j�����6���uKm	;i��!q@x��4:+β���)��K�6]I���8#N�ù���]P%�~A�v������"��z���u���2�;%��O���+��ؑ,1��;�����~q�ݑnk-.|?��|ei�j�
�� X��<��	����TO�G��@�>[���v�fF���\��O�D�Z���=����B=W'��%��� ���Ff�&U�=�\ys�XP*��AF�2&��ًTQ�ھ.8��q��X�\��?�씗��4j)�7�^�d,���#�ؙ�y�7�'�F�%�4m�jp�U9h+~:�yhU6�Д+jI��sK���7>r����2�Q�[�ldV�����-Dڛ��dǽJ���X礎/?w���CP���L��>0~NbQ,��Ϳ%�i�$������a�ݮ'��X�_�w(k�a7Ahb�Ӌ�^��p��;iZ������'�ȱ�-\K��7��TCּ�lbN��LU+=/�mʯ�x�Ĕx��:�<A�a��:��]�o�s�v��8�d��	��YUoxQ�\$�"=�r��*^��������ME���O���ra_S�Y���l���4�h�utR�^��7������፷8��J
ol�Q.�����VF}�\�.D[=���7�$rZr��Zj���ԥ��n��n�+O���^��I���)���N#@�"���ɻ�q��8���VL�� �F�H��%���:3� ,��|~�[$���Gt�8���A�Y�W�Q�'�p*:N��Q>�|�F/�k�,���1d�MEk�6o�������̮:���f88��%�j��fT���ѓW���H��2���=#[�#ne�}u�e�ս�^���I�p*:W��sy��+��@[�8��R�{��2K�3�]i&7pH��R���#A7tBU|�ҵߔV���xQM�udY�����f,*.��}��}u:ފ9d1s��Z ��r��r�1�;��"�5�T�o
�Go������~4*mG�!�@�;��n��K�و�����Z�×	�'�Vj�_��(nC��E�W���|��
oyw8ɜ���?�F1<����e����� ĹoUz�}h�ps��^���F��H0��Sd�`����-�!�yJ�F�2N�6/��t�B�x��8�C�Q�*���cIQ��Ń%b������ q��!��tk�>�������;b�`Q�CX��{�ƍ������2ζ|�	�ϔ,e�l��� �nW�T��G�,{�DKa�lZI��3�B��z��p�Y݋��C
6� !��y\4���1	&4E`�%��t�<��$�9GJ:/I�9~�8U�2��>.@���]��lڝ
��~.f��{��A���W�<X`�؉y��m�N͏sFQ~��[/�P���N,�=�)��/���V�ڗƦ=��p'�����o{�/��B�
#���wƞF,�-���j�7��6W��A&�`�?C�\���3�P�y�{�x]��Z��7�CU��QC�٥�2n4#-%C����`�՘���|��F�Рb��dX�sp}4(=d\iq�u�����]�M/��������9f���5��4�ϒ��5s�"�: 5�;x�_}���`ܮsz���!�|�a�l�跩PA�%V+��v��� ���c!e��׸���?�.��]ȡ2}� �̵{P�&w
��V#�0²�H��iu�n�iWT��K籀��*����~A�$��s��N�$-�&XY�x�t����M̓w}�������C̕k�y��1	���u����*��_<.|��4�����4�t�w�8<� Ms�^���w��*�-X����5ܙPf�� A��n�_�ݐ��E�t��cv>��'=��,ҍ�\ߺۜ˖�ſ�@\Y���W"��Vvz�Y�����u^�xm���'���&���N���2eO����c���йt�ўo�<�Ӑ��Gn[m��:�!����)N)��O����ˉu��s���.�˺�tjC`llZdA"a}<�pE���p� tV���	�`u>o{�Y3kN���A���*�4��I	evX ��ɭ]��к���Ѳ���j� |�&������y[/�et�P�1|��M�x�s����@��H��7ɟ�ʧ$�< iǢ�4nC%�6��5�^`�T�C����oj���a�;	��c��"~p������.F�z�̊����5�JI9n$ũ��D�OM��	����H���6���G!�}.���x�$���hr��P��?��B�� ]�[�Wd���WC�CG2�������^�B]O� �f6��#�)�3I�ɼ�nA�U�����i�L��n�Zظ��X	J��N�W�6�a�D���y+<\��g�[�xb|�n�K�b9��O����,570��Xy����������0R�WqUH!�F�qdN����Ɉ��~�(����(FR��;-4���ߋ��ES\S�OJ�-o#�Em,n��}]Wk[v]g��!l�(q���������o�nfYF���0n�ry
h6����>{�%�����
����~����U�q�k�-NIM �q��W��j�U�Ŀ;X@w���]���;.��ᇜ	��#�Zt�6��6>��������[ƫ�hZJˎ�
/#���/W�g�$Sg�T5��:�>8HV�ޒ���À����ԿI���v�Tћ)���T�ю�w�Ջ#�;p�`O�``r�6�}'�4:='
�oИ$N�Y㍶���2ֵ
GWj�"®;<��|��S6�Y�~�0����i����\���5�=Gk	����.KW�S5'�͈�E������8��]t�r19��S��)_���uOy_&@f������;�a� �n4w��b�ǀ����
v��"���R��.(�h�����sHv6==�tP�������\�~��C�{̈́��ae~YR�ei16����3�8��kT����-6"Q���TVtu�S@�K��~_�ˉ\���ǖ��E'Zq���v��j�!+��A~�RQ��@�̓GoD0���^X;++�ԯ�;Iţ:��y%�X����v�R|�|C��^С�[�HFY�j�-0��率�T��U+�{v#�j�@�|���u�}To�GR��ˍ2�)�W��X�S|��+�F�C䮳y�-��*�(���uJ���5�I�,?��"��Z�W��I���������Con4���6ѧ
)��W/�)��I�r�M�q����r$ۓq���+jP�A�6���dd�$<v'v��T��-}��ٴ��jbN����x�<�L��Z(���38��Qc���ح�2��?Y+���r�_n֌m[ѻ�.�c�?H4�-��{sFR��i���郍Ǩ�P��t�����JǨ��`�:_����_�Ih8�H�<����+��,��s=p;�>_�����he�ǈ�O��P������@�yǵ���4��HLk&����D��RS�����2,��n��/~������<z$v����Z�M���{����v:�6l��׎���L������=�p��ё�|Lhi�c}���e��ʆ�T�r�u���ջ��ɷ�V= |Fi�p_]�qxPm��6R��)�[ѿt�(�� mM|���.M����]����8���;$�ࡐ�i O~����Q���38�Se5�����\�nD�^���,���8� �|��o�O�&&���4p���a�d��
�Y��z�;�?��ݘ�.o��z��o��B7�y`���4H��3�"W� oِp�f���PEJ�]�7`�w�| ���>f��/Jĵ0g��RI?d6�i7�:x���6�
SE��[��}!@Z�� E�B����i.�V�6Z}!�@	/��R����yF7�L��}��`>���F����X�<�m]"/zBA�~�m� ��#Ge��+,��l)�ړԿB�tO�@�H@�:�w��E,&�;�2��H4�J�� ����N�F�.�V�jo/��;|6sf��C�l%o�1��w���2c71�������k?�!uН��C�$g\�+�Y�
�T�Q�5	���ߗ��bD�l9J����]k��=8uFkַ��$��W���ҍ�*vb$�z�H;��|k���q���3�?S��K�y	f��^�D��`n,�{�qe�	Θ��;�Uxx���O��pG���ҹ���#C%mOј�"x+q+v��98�v`U&����r�cF'�H+��S�i���>1<qwkÄ�' ���l�c+&J*��ꪩ��$d���yu``B��D-�� �1��3���ɗ7���c��B�QY�q^\� W���}V��	�|n�CfÑS���7���k�
�ZQg�[�A/�U��
��Q��q����kuF�f�����qL���L�T�S���qk�y[�\x��}L�*�Wޫ�
V.-��$���sE=��*��ڡU$��yY�X��D~u2nqK�ߠ��7า��M�t��(�V~G�j.��*���BiҪ<е���)1�@3��Q�@�(�2S�^����G	�)a���J���?"A��S�ߠ.u�j�{��0S�;U�x�v@�/�i��'#�Jz��ML���6�]�|Ή�W��,��2��y�5|LH�苎&�{~��%S,%�R`���Z"��_à³u���k�����v��#{/�NI�~2Ҋ�� I�����=�vEI�l�ѽj
�h�(s��EA��'�+Mr� f�zz�
Z14hG6�d���|?�������-F.�R�?pt��7ex�����<��7��,x��KA����"M��V	4,�������I�t������$��dY� 4 A�aVEt�t��B�ex�y/i�T��_���R΀��Y�CT����9e�?COn�)�2�v�Q+Q�e�+�7��(
!�Z��On"�,*o�,Sݗ
��OL�ΓY��fR��.�:������'_���۴	_�I�C�߅���6Ѻ���!T�e0F�VI8�}� [� �_�f�"�Q\Ea3̸�pu�Y�J�F�Ӄ�x��s���<ڷ�\sū>�U������L�I�޼�˺�/�@kc'^W.����)��ˋ$��JW~\�q��w��-!���l�NQ��s ��р�r���i]�8_x#�(m2f7�UDW�n�Z7�wڤ�m9�+vR��ew���·���+�=���Z�&�n@�u��-�@ϢX���gl�w<��A���o�v�ѹz���y�6y�|!I2���7W9ƽ��/|]z{�`�t����SJe��TCQ��H���U�o��C�Xw
J��@�2K�
\��e�sd�_d��R�.6��K���67U��%!"�면%;t�k K�N3BڽF���6�+3a��_��jP�#ȼ|��
靽ZJ�f_���=��
�����������rMˌ/H5N!a~���L0�I��hy&��ʷ,H�\�Z�Q['S�9��9x�ä��|S���=b�O�I�[�$�U/Y���;�&R!SOh���ʿ�\���\�݉����:	���ŕ�P�#��K��z<���k�hq%�M�훭����7Y�beIH�@-TN��)Jy�z�
��]�I��w�����֯��͌���0|�,y���@Մ��L����܎A3�t쇊�Sŉ`:)�H�Qr�|:[��I~���;�����H�{�b�x*�ډ��擇�W��]I���Z��J��h���ہ����♭{��Α��N���B�8t�%���tC(���d61q6xv=0ߗ!F�(#�ml�3�es�H J�S�1Z/���N�k�-�fV���/�Uin�OKX�������;�H�u�Bf����П�X	NRt�����p��cQ�Ur,ME�(N9�W?�,e�������-�L�V�	�b��Ef_�}��������6[��9.z=�ͥ?c��4H�C���5���.��c@P�34^�*��-Qf�>����/2/X��24n �n��@F}���)�M���ѿ�$��x�m�l��]<��c��j.��^[ް&Awy%_ˇP�>O��T}ږ͚�]o�~�@���ed8#�V��0>�͹'���3�l֚'�tM�B���]-���
����5A�m�N0�+/�	w�je����X�T�(�'o+Hbu�v���Y�� �'��F�y�6.=a��*��JD�X#��/�+�%��}���g��L`g��M�*˗^d��';O�/3<jJ��i���~��
��۬�	?j��j&{�4C�R�Z��RW�er��`����Q�.�=?s)Iځc��#�%F.ܒ��Xq��k����>vi�i�T3zH�ˉ�bz�>��i0����BZH#y�����rMׄ�È�ņ�h���f��,�W��
�s��'&��ƃb.H�#�Cxq]�����h]�yCX1`�3s@�V�*��B�R����9��S����:+c��Vw?�9z��x�[������ډ�.^���;�~�x˽ ���V.��ǻ�Z��"��4��k�^���|���ͽ�16"n��Q��DX�Z�|(��v�ʀt��A"&��v��MRs����y-���k����R=2l�T��C�x�0�'����3�k�7 ��Z���F U� ?�5����x�c�Cv�<%����R�v��'��=8�V�(\-,��A�5xZ<�>'�\M��YI(��Mv��5ou�\P Nr����-XI���9��T
[x�N��;�K�D�,UuG����&�"z�p���Yc4"��hK\
bU�Zr��X���.��0�/1}x�?��|��ʵGT"�%��:ܺ�&�4��12P�c�_k�D`}d�}ڊ]��ܢ�gU�Q�Ȓ�YC&�o�@@�d�>B���V�Y��@8x��rFl�z�Lf��LnNf���Nc�RVc+x�5����?����eu+�M��ΰ�/H���tN�,V���9�K�����6����|�n��Ӊ��6�8�QS�.��$=�0V�� nC�l�43���u��?���cs��RR����Bn3��4��y��~$�a��ڎґ �P�C��\��Oત^/:��0�jCp�.�7��rహ�9,J�}@6���T��y9����/���DvQ	�]L}>	�g�j�� ���a��N�95�lB�������h10?C�w&=iI��1��/������e.+���a�8vq� �����ć,l�Z�2�$���l.W$�'����	�Ű*@�N����x�f|��'d&]L��(c����r�52��I���a&�#Z�a�i޷=u�f7�!�}����n���d6�;>��Ft�՝�T���� ���~���D"a�x�M�����o�A�&s�>� @�CV�@|�)���9������F<)jAa;5�+'ǮTn���g:N��+���1Q�1~�-�bC)�r�0�2-�DJNR��uj�3�s�3����G����.�ܡb��s�%5@?k{�3��������r~�H�qG�I1!҃�),j�;l��X�rIVҧ���zȯW;�پ�Gu
����BN����������ܤ��)��n���ܹ8����j�U4��x���2��i���P��̮S����bn�������6�xt�қM��}��B=xg�H%�e����<.�c�'¯W��D�ɭ^Ȏ�X���T���{ �rʙW�]4��C �{�V�A�͢5�P%Z=�Be�D�&�i{%�&���P6��g�CKj�pP�q�G5��>Bx,��zf7mg�ز�Ͻ�4 �@&=ʨ�"����M�@|%p���$\�#`��0��/��	co^"kz���/�Qc�%��[F����d�D뻘�Dα�tSx�����Z2��=S� ��L�M�Ԇ<m
-0ɀ���RG�L��U�^�_�'�ey����B�+7��8�gjF��L���l-e.!�K���3J�s�e4�����ַ�+�>�z+�!Wl��
�9dW$Ux��s�M���>�0�K�ZC���fW���zP��S�˽/�XB���7�e��}�������KZFy�r�u(�บ�F���f��.Ч�� ��9q#��:H��v+.G��S�)����0�dp\e4ԝ��v�ֻd�?X��7��U<��~�t�$1�o�G�f e�E��Qr��	�y�a�Q�߰dhG�3�eb�(v}��B��c�H�ph��� 2�E�����_==�2cs�X��}���ݩ����D@0*���6E�p_nAcK���U��G3�p��%:]��"Yݱٱ/a�K���?��l��g~�$���Y!��(�8@��`���ؗL�7]���A�v}��ل�3��;�q�� ��vs�3[)�NzLV�zU:U��w�#����c���ez�5X���m�S��#F�D��O��9�F��,���R�Mh^�V*!�eN o�-���8�;ZA�˚ӥ��s*� [�]R1�O��y'��
M:����t`im��wI�]�+)rȡ�?�vK�p/�=ū��˷w��/����"�~6bg9!E�R�'����8b."��dw��8c7O�7\[��M􅼹�98/L�:gn02��أ�tnM��3س��_������R�*���p��k���gr�=��ųC~�]�z������vw�!��f��G�K�`S�E��?�ԭ�:����{����������$����E8�>j3�l:��.7ʟ���S��C�hy�HݿM���IP�YJ���J��6h k�}.��ۗ��'h(��[瓜�9|���_V����٪X�������!"}�llR�K;m�ސ?m�Х�N��Z�5��$� d�v7(Zum��Mȝ-�f�-+���_	F#tJ96I�˴0\s8&�殔R�6Rp��F���)�Pٯ�&$aؓێ���0��px�H�I#N1�ܲ
4�����Z#B���C�<:+�H%���|�ŦP!ծb�.�+I����e�/��b=��ݲ�K�v��?"~�(\�^9bU}f���}��^���j�m�.G��
g7!�T
�={��6���H����0b��[���X-�j�(�����T�gM�(�
��4���?��Z�_���W�:�>2�e:����!a\��=}�84R����� �[{��;f���}�xEFoր�����<4�2&��
bty��%��7��!�jٝH�Y��Y�u�0�7�9~Q�ZG_�y��:C�A�狪�8�-�Bufݢc���d#Ky5]#�~�l\��� h(:S�p~�� �Yղ��N��[׍�D��ŢF��� �f���1y���B�i]d/�"Qn�^���>�b�c������k����V`����D�D�^{~9�.���nRW�N�B����`�FI�o�*U���� ��S���Z�'Aͱ͠a���ɦb�HL�-�zK��d��J��Z؀���O��u &3{�GKj<��T�FO�t[�e�n(��g��i�Ϲ�@I��'�\/?9՞��ʺ�p�1�˥t�*R�>�"��}iq���,��6�^�ł1���[Iedv�+m��@\+�L;�~�����Z�+K�`�fL�O�����,��6oW�*[E��I��$�j������	��0A%�Rj������ˮ�S��;}�kk�TҽF�\������@��`ŭ̅��#�9��o��A��\���k ���lRR����h
��l�O/";��3�A��F���R��~f��4��^�5�#/q�����XS�T�)d��!@�����u�K��ڧh������E�q�a��b�:Ƥ 9�+�Үw��eè���:[*��M��M�D�X~3���$ɢ �p.�qnd�����Rw1�E�#�8ʒm����� �$�h�%
U*���a�^���d���3���������W$2���{`~,r��`�_��h�;��;#{`a�O~���n�٭�k&���Z�E�t����ҳn��`_Y������]�1|n*D���*[(��K�S�'L��a�D(�|��L����Vx������%�.p�Y���|����x]<�_��W#`r�]�Ns'�Y~�o�n}�f�d@ �2"*���$�%�����c�I^Wg*��:]���J�e>:`�b����?�=�[�py��C!z����m�}(��QFI�3&>���߉���T�<�cPd�J��c��MVe���m;&g�gځb.Ŕ���Ka� ��@���b�Þ}1�� ��V��'�*���#�'ox��_�+��m��O�K�k�X`��!���l�`y�? O;dL���^=_���[��cd�\��09�KZ�(�@�t�ûr]s����`�t՗�o�,oե'�@�7&f�S/��]E���8*T���%cNŴ���T�d#V̺D|�ÙG�y,�-�Շ�7�)E/�}:MRG��p�؂H��ڕ�)�~���qL��0M:��̏���X��[b��g��@��U-����3_f3i��k��]4�_�#�[��ˣY���Z������DǨ7���W*V/�i
���~2[��,1Lя�mοm%%��`~�6��S��O��
s�3ḏ�}tO�j���ʮ���>���e���^�P
e���D	<���Gג�<�[���E�����Q��ǝ��VPA�~�J��{�2,���F?c�!�pt�E���"��U���)�_�7�P|���ȉ���uCk	�z��*�W�ᫍ5M;hpmk���2�5���}v��u��0k�G��1/��?V��fd�e5
�.g2��{������m�v�q���A��+��)	��i��%���96�������PF����1�.;��E�,A��jH���s�!&�D� �����M�3����e�f�����P:�>X�j��:���h�
�ӣ�'�wH|[��c�����9�W�\�a�VJ2�B� D�0Z	��j�����Z���Ԕ��ZF�<�m���ܯ�Ԡ�^~[@�F8�����|�ݕ}P�'��et��4����W����~�N�U�,T‥�'�v���*�������َ_�D
P�?%���]�Ā���y���Q��X`';{�ˤc���]P0�>����ۘD�]§�T��K�罎o��x����.V`p5�͚Jj6��an���7l�%�9ae���GQ�.��4V��`����ɫzA7�c���]��^�NH%Z��A{`�5rls�r����n+˕�Fù�
���B�Y���j��V�ps�E8�����G������4��[_�\��v�v�����@kCoR��ۭ4��}:�B�"�c�r�<5�A����w��ا���P=�<�;��~�i�t�XȮ��OEƏP|#��OEw7@B�B�),�܍*бxݝ���vČߥ6�`���.{��\bߑ@��!Z��%����礭�(��\�V��m%C�M�-~gO"gt�Nj��ݍ5���B�W�)�����>��n:R�#�<7���~������w~��<�򋧟 �<�!����uK`�B�E�3:@c1��ɲ��q��7s�X��[|�P�/�}@����6��J_h7q@����0Gy�����p����+���b�TI3�ׇ���= M!x��e���>z�{q�(��+*�3�0O�q��E��WX�NI^|�y�l��`��)vpf�5�⟘�ՓpXBۖ�`�G���M����i�h���������@;Af�PbJ�85Ut_1c��gf���3?"�����^��^�q��������`��V'�?{�;��@@�a�+,�P�2ؠ�;Îy�U�8gG�f�e٠�VC���b�\�#��hp6�{�����P�Tc��O��[EZ�A�v��shb��~�E��N?�,�w;��9�����t�T����x�uEQ(R�>�Q�e͇�^H�Z��	�[Um�ϯ � �����&��$]\�q�9��М�lXe��BW~�F�J�it���*�1��^�gTc`K��X��4��*��=6l ����Q�l�R���Ƨ�H�����륌��A���E�o���J8L��N麎�
}	�^�n�^��}�P��L�|��ݧ儫0V�pi�	g.���crwȶ5���؇Ǐvi�˛j��T�N&��`i�2�œXÊ�K�D�8@`~Q|>��ߊ/f���6<���80��˦Ե\0�6-�"�����cd(0(���R�]xd#�q��Xfr�J�����zT ��^iD�t�/�	��o_9aD����Q�N��߆��INʵ%�;.��{�ӽE�"���n�3�TI�ʑ#�qX���?���+�m�j-E�V��n��9)��KR�\�?� �?����I��	m]���7#`����=�?��M�*@G��p�1n�� T�T�,�\��K�in�1~��+>޸����`��xfa4@�F*�'6���T�P;	�RDi�d�H��@�Ҙ�(+N��N�bM�ܛ���^԰�VK4dށ�����dB��q���no0yx�A������A�t*���!��*xɴ�;�"f�-��ʓ-X<�>I��˝ '
O�}\P�RR^�|k<�VU\ �x��lU��5�p���Hyr ���Xc�7�d�o�VT���4ZR���ȁ��0? �;��K����e/a�L�S���t�H�jiF����4-Vw��(v�,�k����Y1�$��g1Y��<s�Fт����/i��`(4�{�P;�-l�6�u,��E�ј�K�S�읕���P��H#�=T'U�@��`���{ɕ��h��p�^���n4��ƾ��'1�����	?��]q�s{ѹ7B���	�\��bd\�N�Z#�r; D?��s�ܐ���D%�'kn�NH/�a9xt]92�r0�DT5/�����f��u��]��3S�df���y�n��S�� ��h���ҠI�q�����GJ��k"9޸mH�\]��RIa`8����e��j-N�JV�nw;����9���X���2��eg��%�W�|��D��1l�'1�⩲��<�׉�}"id_P�����j�m�u~$��>�(}(�*��*���i����e����T�O����#��n�m �G=�O#�g�^��%.'�M�A�&*�D��tB�b�}����Έj�v@���*#O=��� ��ػ��·l0�Y�VL��C7�m�b����	Tz7i�V�;!*y�Z@'J,�;�l�	��0��'>�� |��k�F�{2�40�݁D�e�K���jA�q�a���;%O5 �14!�d5?J"��d�{�ٕ�%i��ؾjt'tJ"�,��G#}�sO�?�iB˪d�a�k��(�~�bB�J�+�C��wa�?d�3�@0��\�䄼	C�T&l�8G4;h��7��LA�f碍�Rt�.uұan�GT��C��bIVg�>"�t]��%H���4���9�|�A5	�)��K9��v�m�����	-��9'�#(�KL��E����h_<��8�j!g7ܸ�Ê� k.Oϴׯ�ܒ�"����|�/��b(ipĲ`��MW��~�Iv��t�9|+)��P5�R�=H�&�9����+Jxޮ���E�5ı�B �A��kً�`�'�\frv��9,�(ve%�C�ji�+�"�4�:��t�)+IU�ϑR�+�s�c��$@���9��ܬ�@G���/����8�gZ̊�aμ3��j�*���4|�`TK�j��˯G7�z{��R�KxD�|j�\��l��{_���7�So�i�K@<=`V�^C��Cdb���A��<"7��t��m:��k��7҆���M؉K��ӈZ�1�m�U�нPm�Z���>[DU�ցv��J�ݭ,�zhxI�X9�U�W6ܨ�2"?,DB-5*�ϔ\DS8(8�x��ew�mH8c�_�v�v�"�����5������+�t��R�p�y�f�.ݲu�����脡����ӂ��v�[�T�J�N�/:���zҭ�������L>�8�b�QL�01��	�`��; �#E� m��Ǝ"�ݚ�����mL�E�Վ�ern<ř�-)���;�똭n|Y��
�p�y���3�+��p�׏Eg�|�6pu���n�l��J �|V(�S�X'^��|�lu�^9��1��}=_�c��M��蒓G��9y��g���o�� ���`���H&��L��\�2��ANpmy�,#�_�JR��pu{�Y����宅�sp��~�g��������`.�b�x�N5Yƞi�a��g�G6��b(v����Dw�өb� %�����3�"a:�����k5�!Y2�����'@��Z��M�o	�
K����:P����c��A�!��96)3�NF]�-����}�7K�ecY�Ƌl�G$U���^BG�+�I�����('݊;�M{%�X�|F�veZ�ʡ��'��L�s�ڨ����ux����;���/V:@ҷ1����ovY�����ZQ8w��X�z5Al-�<��3�����}��EfEJ�<h��N�@q;��ɮ�]'�&Y��o�R;�ޯ$L*�)����
��V�/վ�Q�H,p�Np��/>��ܕ���� <b��84�1�q:�d�%�d�46��|Q�s��7�`��q����7�&�p@\�����u1�<ۼ�|U#;^���V�5���#�8���h	F�!e��s��|	o����NL�T8w7HT-o=�Ɍ��S`>P�}\�]q���;U��w���̧����HQ	硚~����6�����
��,gW��݌�/W���=�x�������y;S�G A�*11zh�w/@@��j�Sw΀�z(���z�sN@��-����</m�0����zS��4��D���]�d��`aA����1�M��1D�aM�[A���i(�6g(\��ɣyOM�zȲ���ӈ��ݣt���	�c���)دD�پC�f��j�}'k��}1X"�j����&�EA[;�T�&E�QzB
���7���H���k�v~ك��PK	-a�eN��c��U����Ԛ�T�`�	�]�������l�8g)����>�=Ԩ�]1a�r�,�CH-���#u{̏6�]���x�\{�
"*h2��aP/��Inz��晣��v>����Q�	r�s���6
��)y�I��?�UX�G=,G@�ؠa�Fk˿�8&��ɣ��)6��@��:
vX;HI������t����̨#νQM?���ܸ�N/�����\�Ӭ[�o9ZiǨ�M��,��T��z�)�淳t9�S�;��UO�
� �1ByJ���º�'{
��CY�����u�MJ^��X��Ć�#�K��>�H@|!��Pm���7�f����"�t~:�fB���}T�2/�-�+�J������p%s4��GA�t��bu44�!���5����I�T�wkz�_�_�ɻtЉ�n�2�-�^�o�'�>�p>�<��(�kr�O�F!��&���O���;��X��q�v��D�Ҝ�-�]�pЗ��S��!K��h�� �W�4���vdn����O��^� ���p�Q����+��2����WF8$�a�1;G7B]�[PF������B֩v!���� ����/��Y�M�V�ԡ?iL���0���|M�Wr^]C�*%#�k�paBJH�}�v����@�TW�&JGo���]�)s��#i6�Y,���ףս�dpg��M�oP�-c��p����L�in�T^��DX�����&g�5��?���e�K���"�k���7�����
H�` �}��ptE�V?���և��J�`/h`��<�758D(���ޑ���(�s8x=���6P�<t�T�LK�S� ��U��o��&%d�3�e�� \+�a2�͒]�0�#�T����c����֖R]��m���s�7�,|��?�D��M;�xk�%�&Da>��B,o:!�:����!dX,�kYD��.v5�r쩢L.��`��Z�7>=9�@��js�'���[�V̓#h��k<�L���G�� !>�[qu-�Y`%i-�9��r����$g+ɶ�5o�O8���o�p�OK��~2*���'��BUÈ�Dщo�N�Dщk�~�Z�;�9��8�o
"�Fi���(��F}"i���Fᥩi�c��y~��6{��$�ԉRB�\.�tvL���#�V,��LM��fA��,�$Z���< >���r��e�;4��<)��9����Q+�wɵ���W.e�q����{��P��֣��Q�R�,�u�Ҹ򁀺�,:?>������_TV����v����R�X�3E�èH��*z&�T�I���Q&�h�H��v3�2w��b2��D��Ś�V�H��dNS�����iDF\s�Y$++F�=#��Β���Y�Y[�λ�b���ß0b�.��\�h��,:QL@%��b��o�3�6�h����f��|�O-Zᶮ��a;PK�ca���D���gܩ.x�&���]|��\p� �N�sW�jQ�|2�I&
�U��2I�q�#�����K�PjM�s
�Ӱg����s��iu���x�S.����~���:�B	�����_!��[�Z�=�'v*�i��g!��+�^�֧F���-���D�dDw����k�q��pok>igީ�a�	8�P�0FMA�����5���b�^�tt^�P���� ��B�|��';��Z4}�T��\?'���<�پ{2R�����+qg��6�c���9B;�d�}�k�yh�Î�ifo)�� #��y72l@��8�:h�X�Z�=ZHj3:���.��	��h�,�����0�
(fH�:'p��>y��qŊؽ�����*!4�=2����K���69�ҷ�X*Qfq5yi�w*̆A�����f�{�2�J�1��O1'A;�k׮���S���������"������8Uw��X�#�ֵ�0�Aĺ����i�8)~�ht��p�Հa�C��`�G�w	�xL9 {S0~�|u���w;�X�w�X��ܵj5�[�3�26�����X�qݍ宧���T�l�3}�5���Z�0\տ��#���AZ5J��J�»!�&Fpl.���y5YT'�:^�,d9�^c�q,��kL*b^�ƱAr��q���1���6��D+��堂�*�ٖ9ީ��[3Z����j���i9*�-m����ck���՝��eB^@jk�l�,gx^&�9�3�E��Zac0�e�)h�Q�M�sڗ��0M�#0� 88�M�l�\�_���(`�)T̂Hl�fv�wq�g��8EP��z�zV��~�n��K��<�>d� o�Ț�_%SÆ�ZͲ	.,��if��E��B4��0��lG804��N���˴��zM�p��l��c��Li��F�D�a��v������ngf.���J|��3~�B^R��o��m�Z�N�F���+|�4=�5�St}+6�i�˶[�V/'M�嵙G����WϷy;�6���> ~�l��M®��v���(z�o)��H��KA��B8}��O�v�G�B��b���
�V�x4�$�2��+ u,�e@��?��S��g��WV}����`l�DI�Da���{�
��Ǟ�/FB�}�Gzꑓ:�g�n��fdF	`g�h_�)z�D��ė[���.۸��l<K���v�eb�Z�~��9SxQ��E��M����1+��:��e���"-�cO�G&�W,��կ��Zf��Y�9S��;t::�A���|��ZG�FR�o � ��k���5;�h"{R��mf�ɿ�O��^ú���uo�E�W�1�"�z��@eKh�b�($rxkq�P��'Ν;׊����a�,�g�X� �~Ɣ4��&���ʰ%�s�*	��dM�M{�Җҥ�{�O�1����hEh���>Ġ;��*6�9��V��v� ���Ѻ?v�+o���ةsξ�R��֖�g20�jS���$����Ђk��uc8�͵r��[�Y�%a{%#�n�˓�I�$�lC�9���K ���`��qAO��1.q�x���)��ۙX��A$b�{�=2��Vl����w|���D���/whL0�hD�g)d7��!��lX�|�]�Z%Gmkw͍�IG���<3m
�J�Z!q��nM����3���'�k����	'�d_#���xF�NY�E2OW��Z)�uq�?3���>�{*.S첮�n� K�Nd�i<qt���w�{f̹���!>!����:F¡#�ɤ!"J��5�5�,.m���y;C���_��5��<��pډT�������L�,zǙߤc�^�|���3�%k7��QS����D�78!M�my���H��WR�j�6����y@�4�/��śM�Jp�zw��m�YXA�!�'#i��~��dz\��B����i�-����D�*���$�>eRc�{����^�7�$�c��@���YߦlL�G�!�Ff~��ut�z��ٟ�з�ǿ�ah�2`�[?�s1Em�0��X4�\���)�I��!�3(�1�q7���wp
�y��]M]^���B�z� j�a��m.�/�A���to6]��*��zu|����N^��g:Gq�:҅���W@�T�0^��7�d=�2}�@��	�j��ch�l��V�>[�/�D~����.�� �&$�^f�=��n"��5�����M�	�Q����X��k�b��y�L�!�{�OT+�V'�Z���
��~zJA��G��,�����02��	���@���L�싐����e�_hL�����0ϯ|�����[9l�n����%�� O���*3�]*��#"%f�ɕ�F4W�GE�}#]Y/-1E�dC�;+�֡��'��Is���"��@_b��pl��G�����"��'�hM��}Dt�^�O�-�j�nzؑ����8W8:Ð�=�U��}����r�M���C��x��M9�j*Z'N�0���� uB�MKaĆM���XZv)l�1�@��<��E�w��"K��[4%��cY���\JM�K�G���Xʴ�޺�h�m{T�qf�E9vu��mF���{�]�.���̚��2l�&	ݭ{O7��6QUr�l�c�b��i|Yl�z�Pu���۱�Ѝ�w=�B�bUD��G���T������t4q��!ܭ�BU���&"�m�Y-!�Y���L��<���6��Ȩ+1$�,�H{ ^�zY����`�w��ך�����4"��E��8�;��j��p�H��jg�\��!h���Y�iJ�݁M;�y��	�PӴ{��ZI��4rZ7�PP���):�}��<� 劉e6����ޢ�}�{KԿ��8 ����sf9�.q���G�S���q�x�ñ�q�����~>G��W����'N���|#��4��k\~I�pmaCR-aDP)�����x�誌r��ʓ<�Li���CN��w�﯒���,�T���R����~ؒ)n�G_�@T*r4�0���c��[��N���Ѡ�xw���'��	�K(3��g�
x�E ��_�?j�Q���t_�:K,�ůа�a����#�?z����Ųu����Cd�9k��^�%�񸀌7��L|��� �7�O�n�\��Q�,SE��_���aI�X��Q�|�Z	9`���c-ݕ�|��Ef]�qX�Fu��Z�z�.�y6Vj�JGc�V�;�)�"�W�{�
"��u��w��(=��Sq�>7\�K�'TD�6[��Up!��E5$H���q)c���A��п��z*  �d#jnr�hw�&��$��g`t�%�|�M\v����d�D�3�P�T�^Ua+��-��<CwL�5<�#�
� (\�u�����6}�I������N^Ϝ�O�d�}���v��xlFt���_(�0�r��i_X�ϗ�D�V���������h��ON�=iNr��+7H*��M�hP5)�����t���r/g�s�Os�F���q/Ѱ��<���é��		�!�* ��;�T|�U�������_�GhfX��d@�����TI#a~m/���5OLM�C��5 �)M	Z�'�g/�Utp�\� �������	 �C\+%�Dؠ-�D4�|�$�q�PKc���{�s� �q�j|b@������2���xzt)��!A��8��Z	������P'������\o�c+�G����qf��1������no��$zZ�>H;�7��uP�������I`��p� m�ShH�؎^��&*���Cp����@>b�A���$��"�GC�h+	�L�_C��R���ۅ*x�o�3��Ѡ��껖2;��av�F����N�%+�(��ZD)}t�)�p�6�>X��ҷaHhV���&��H#��y F�@e!��/��E+���K��ya� Rxd-�-F ��T�
pzS0I���8���?���ѝ59���u�F��eJC�5�s��K0��H���` �*26�"7�����A���:l�ТIz5�#��`,��kބ�\5���ʿ+�^�	�#������"M2�Ml�mP7��#��r�aY,d�9�}F*�=J�حۘw3]�|�D��:�C# �_-L��l�$~����)�8P�_��9���"!�E�+�#�(�ucY�	QY[�����}�p�w���1�\ka��yp6g��sѼ�%%q��Xw�q�M��ϐ0�D��? �s�O_ZR��{�T
��E�]E'�+-�řږ�}@��n��ntH����^�-ڞ�T��92�.f�V�w5�[��-���^�*�[�'�$U�ɺ��Fu/	�TO4�����h�EQ�xü�(�f���=_�Bp@�.����A&R>����צ ��-�F�N���01�\�$��?��(���Pls�t��Ag.�VYUm`i@�W�_�l����'�Dč�<�!�����.�lM��^��	'Dޱ�ŗ`-�^`�V��]j�!Z����ǁ��.�`}|�3� @���x�����<���|�ю<a � ��u^�3��@��}�8r��?}�}��QmɄ���:g5��X?������K���zzBc'���ڲ��+�eO�B��z�e�}*Y��(CEk� v�����H��-/��4n�_w)��'�ǛtM<ߒ
j5� ��|6�ӑ�qO�~X�l�Fٍx�y��o��)*a(��}<m�p2J�n��"�����D*��e.�'ZjF�t�����
�b/���0�z�3��?^�A	��fL�D��jI�b�,!U#�zZ'ʍ8ڧia@��А�G;e��熖�2�c(9�t��i�݄� ���$q�>�ũ\|�
!-�2��%¾�̯��G��S8{���H	�1�3Q��I�k
+��Ó��l�O���h�+�s�s�쳏�栀K��?G�����Y��T�����#�����&	x�����«/��8(ӡW�;nF�����i�q����D]��X3)I���f-�|��]I��7�2oj~N�k���+̐���ծ����l 1�ȑ��i������cx��t�J�в᥌��*��$7����P����%��b���_=?HE��1������.׈X�a{�A�zIdl�ߡ� �� ��2E�L����*���%�����[4y�LZ����-�>T��:y�h.{?,��Ŏ⽙<08k��$ʟ�G�|[�H#��n�- ~Y����Έ`I$G��șz���<?Xʒ$�zXB��K�0�&����t�Eg�
T7`�L1��F4�P���8�O���Y�n\��d��_q	9�(�QOOy���6�2U�� W0�E�E�� ���!�3�QەQ�iԂ���SW�dIE�3�kEQc뷻ѷ�� �uD�hH-V'!s���Bs[R<R�����zӇ��1���/�*��(�ѽh�|�����Pi,h�V�s�)��~�80g!A��8��b���;�7�v�Lj�YJ��A����bD�,�S{����N�Yz����#�K�򽇬��}i��9����?gC���B�������W�����T��M��#���40n$�A-E��+�i1��1c��<��zb�+�9	IF�WN�'��^|�6ORc�<ߙ��EW,�A�g+�����~�N��G�CG�w��K�c���Obw|gL�4PA�M2c�SڛЌ��e��L���g�?[9��2"�9��]=1�7�֨��:)HŅ�Pl���֩,����|��������ؼ��U?yH��w��O,Թ����� w�Λ6~�6��������I��h|�B�I<1�QΝ���1��Dk�@�#V5�ښ�G��B4w�a#7�G�~)���������8'jX �� ��S�	BIi+���Mt�{`^�̒���������?���t�Y���0pN��9P߇K`�_[��p<�>4�5+��f,�h���m�׎�2�����M�M�kN�W� 8�։�|��/ӓ��Nw�:���1�?��!]����M����]�����/�� �X^��2C�Or��3Q�6�Q�~�s���.���h"�3���|qTt�௙#质�; �}N��EUǸߊç�i�ҕ����-��͐ݒ�u�r�q��SD���;�������&����4q�-(��eV%����ú��e��QMq�g�&���:Qɨ0��Heen(*�kQ$�'���{(�O�>Ns�M��ej���Ή�lhŵ.�i��Ȳ)ߌ�'\~���Cr?w���B�8+Gk�?�?&���j�M���g��HQ!|����'�P�'@��;/<��ը���V��k�B�2�;�w��x�g`5�#��B�=��B���>;�D�ξh��&�8"i_tj�b^�t��i	��a��ʴC�`'~0G�ﯳ)[G*� IP�AS��"C�H����t/�bw>/��zJ��z�Yc��D���烕G�e��c4�_����A�bX�.,޼���'�$�!�@@��[�MM�i�T���1��Q���>�c��)�8���"�鍻�T�LO�����ک<��e�А�R���~���y`�=���1/��z��u[���#"�m�Z׀�e��L��E�4M޿�vяZ�J�2�Ѳ [|�n�|ؠ�h��L �壏�>�7���pll"��.�~�>���Pv��Ie���ϯ~^�TT�!Zx�F%B�ʢ�B��}M�=����/����]�qUJ��`��7��7�^Sp�FE��<Ss�9&v�1���.ˏ�l!�͹jdm���!�^(Ëk�'���>�3)o���Jw�W$����-��7^<���ѐ�K���=~$�GGB"x��,�e�-Q��ee��>�_xB���M2p�Ѐ���D$��r�pZ�T$ƥq�g�iY,��>'I�(&�u��xW�9�M\ZUFWc���]�ގ�4��-�N��Ʊ,9j?>ې+�V��:����c \,=��ݸ�{��a�`/(�o�3���ܝ>T�����tbݹ~�"���M_9�2<�B6Ң���F��,?��d�I�L}�w��Y�0�v�� "А�v�eN;�p��ط<��5W��w�����$}˟ސ0�����o�n N�5����<T��=H�ϸ&�=�H���C�hv&$��F�I����RD��۱�ذ	NenD��3oY��]�7���$��0j �*v�yͮ�굽e����I�1�3KЀېY��ZL9�<�|;���1KAT2���e��ro�۰����h��a&�"J��a��sl%�o36>�iĮ�BVHpGTO;3S3���y�_�,�Q���UQgA0�<X/��d���"0�iޅN�(�;lܔ�yY`ݫ�H��vԄ���������NҁG�h�Pȇ�[^-~��R�c&y.TI��?����zX��̇D�7Æ�x0-)�./^^A�u�5��E���T�b�*h��ۍ8˸�U%�����r ��}�X������t�j�5A09�d�����/�ͦۃ}�K�R�C�ɀ�ͮ�t'���m��f|��K�D_���IP�t����@�f0��ޝ|�`k�K����k���}�2uctCf�n9�o���=�n'��nЬ�Z��M���a��Y�Vғh<���c���M��b�C���Yu�{��@:���[�Yh��k"*����8�#�9���@�51���R�D����Χ�ړ௘�$C��p5�Q���� ���5���mbĠ+;�$t�0(��q���֘�4.lK$�����Q?O�.D�*�|f�=�5�vq*oY�=H�醰qT�|�b� �T!��c�h�̂Z-�Ff`�ܾH'UᲦ������?������`A^�Ux��&�6�9���~c+�+C��O�>��C �x`�����7y:��왛�P���A'xY��("��b���\��XG� J,���Ulr��}���Q�d�|�|y5֚}_��o��T�f-R-��&���� �7�C(� Tz/�ݐ�� a��z������C�%�q��b|�p&��iWO7��h��h����9�:n�Y���Ƨ����Ȍ{F��%�u_z���$���VgOyX�Q2���i��ܬ��j�B-I�UG����&@�3�*�L�ܘ@D����J>�@�ЂQ(@
��Cɟ4�*/3u�>Е}�jH5A�)��3s`�l�~�>q���@I.N�~�t-6�T?�����>�`+�AQ�r�c�N,�8�5�Ywjx�?K�˾Ҝl�ˬTQ%�G�~9���Z!dpu{�
��5ɮ��&$�E�M	�h�o[��g�߷��6��nk�v�Z��?[�p���d���3(w��v�Y�a{�
r~�𵪡�"h&8i���Eiďmsi�V˖���;K[�=��x�O?�}���aTbx���;Fau�Oc�5����2���1�,����ј7�$�t3�i�7x�7�6�>��]���ڱ-�7G0Z�A������WA����-�k�Q 0����E9�sD���;LOVRq��V:�_�$y���z`^���e6�����@;U��@�&x� �������	`2��*j�L�A�R�bĨ�;)�*o��ՠKb�b��Z�v�AձFu��oi�힫�UkO>�O`6�������_��,tP_�0�tD�Ԏ��-�rǩ�I�!@��'j���x;�7.�|K��˹�4߆�yZ�fёn����a�v���T���j�-�c�7ò�ZĜ
�I[b��w�:]��x^]������x�L����E)2���db�8���F3)�(hTJ��e^��!��D7���*��/�]�Dl;�	ve�,+�b"�ęˉ����<x�I�k�����&�a8�+k�"A*�˟�����Ƒ�q���M|�9}�]��[Ӄ�e95<�B�����(vv�x����	��8h�.R�1 ���.��ȥ��'3�čBC��Y`������5T���F�^H��M���W�]!"R�����	+F�RWM;��܎U��gkx��p�u�R�G��z�x;���ϡ��?4)�i���BdtZu�B��2�����F������G�1cݑ=A7�ON��+�~|�U��e">�l�B5���ρ(����+Uz���ea��)�jDY(Ƒ��J���9Ƅ�Ih��׾���Y=��O,-�\�+�"��s���%�so|8�1� � ��f�%�RI�CjDM���2��#��1�T&�-�uf���[x��?�E��p	��{�a5p{��=����骬F�F��:�u�#��Cqג����ԥA���m�%�����2�_�}zv,4���muT=8����1b���j��:Q�,B�<?��0���j�_�.��s�p���D}5t���)��r��9-�NMb�g(k�� "_��QWO��<��ׁ�{�Ho.�h��c,��	D����goB��U�I��я�5f���	�X`���ō������}��K�����.��b y8�)c�c���̶%f�� .����V�R奷�(�G�~�i�/vQ_�w7��7��N����fS�:W�9���N���������WA�>4�g�j���Q0OUf��ƹ�"���BgP��JL*2�ub�^���V;����]�B����@V�A�[Ȏ�Z{�H��zZJ�P�6�̔M�����#�ap����˯ �l���b]�T��F_Xa9�PƁ��&H�s�5ܰm|�.���u�g���+F�v��ˤ�Ҫ�P�)~����AJ���YG*�/��8�� ���1e? ��G��� ���B��E^����)�,�z�l��*� e���PN03��N�J��kZs�V�׋�d�:�ںLw���]8�g����ZaG�����h+��`���
�~,vF�Q=(������}���RѼ��S�"R1��ƃD~�_^&�2�`N�� rae�X�Im���8�@d���F�<�
g�Z�uG�1��+��ԭM96���%if��2���H�U�]'�5��%S���0F2=c�Ag&�/�H'a�0��0�����e߿Q��N��CN��.f�¿t�����9�R7��k+W��T�a	��;��M��u�a[h9��v�$[v�O�㚍O����"��ew$���z9�<�q�X��ɔ�|6df�1���I��L�Pn��=�Vr:������e^[�NS$L #=�J��x�5�Vz�p׌���gw�����<�e~k �G�bW ~��&8*P?k�%�_�}�ДSGi������iE����
��#)|�>�/��&�������(UMd� ^n�V���i���.*������Ymd����/u�У��l%�W�}��j;��u�����_��=gHB�#��<Ϩ����*��Ű{���I6��vB���d?�WB���9�X,>1"�?�(+Jl>V�c$E���朡�ٽ?>�w��
YW<-6dr;
�8:f�GP�������yP�]��8����v����$���e��'�z;��85c��*��#B�6���Β�K/=��Eh�zz�<\+m�S7��~!3L�X�1E�nd�<�lwxg��.v@�%����-2Y��\:��x��ޖ��(ǜ�d�r���~=wO�~}�-�Z���M�P1��L��*��ヶlr溚�57�3n};��4�$0���P��K'��ǁ�ʃoJ�}M����vV�� Vr-����a6y�𮖓o:w���!�>�T���9D�A�\ak�*8�M2mV?L͆1�#�A�f���>G3�[�T�gz ��6�Y	����?6҆\g5|K�(��b�e�89DF�;�ִ���%����=�d+�j!�7����BrXo��L3��oz���.�?�(��D��\��n,����\o���,F�DD�= ��5�i��&�Чx^���W��v����I�ʡ��/��U�ge� �? �gR��Ύ��V���\,��za?�q1H���茍]H�.;)�ٲ�P=�����2�s�4�njO�����x��~�R�p��My�s�L_�[9�9D$�)$��5N�\�rҎĦ4�MO�?��n�^G>'+����r�+4��bD̉J"yn������﹪���������QxE���ַn/}����p#d�"�Mf'�g�/�'t6~#�FX�,̼׉��k��g�f=���ČM��R�Fuh���`
�͊�4�0KZXU!���q6Шi���3eQ�NƢ0ּ m��ȇ�H�}��|���${�9�i�Lm ��εC�s�S��<�1� ��� �psN�������>xb�72v�1��II
��6��,M�tn���]�47��}��/[��ZM�G\Լ(����x�v���b��S���_ao~�zʟd�F��©� 4���o2�t�X����}~O#�S}�	w(]Ck�UE7	V����f@�^���t&<v�/�u��C֙L�k���뱑Շ%����q!#��!�s�������+��'���Aj7KƧ�AU��E��'�BeH�e��*�#�#z�ɫ�(L�m�H���P�sw�Ӽ/f!��Lj[?ie�Dx�~=�{b3dGD��]���HJ�b 09X���>����M�����'ҩ� .��V4j�����ǑЇ��� ��8D�<����*=����z/��]�
��������p����ƿ1U�r��sF�շ�i�8L�/��RP��u�/��C; m��/�2���1d�T�wV�*oY�(�ب)���*�r�0�ü%[H.�p�L�T�����3���8��r�����ɍ�E�߾cų(�
.^��G���;�p�qDT�ǣ^3�z|��B4�eC�.?��
�+�@]��.p�ɫ'v��h�bQ�b�-���7�p�0HkPl��g�$Y��CpO'��x�/��5_����^?�Z7�����w�簚Dy!�b��M���]Φ= $�u����,�;g��9UZb��o�⢿���V,� + ��u�%)l�#QT�pɡd/�C�^���
���Z��-�������@F��d��ְ�\Qd�ÎM�2 G����&�9sT�?'?xM(6Rң/�b�&���Ny���L�ۖ�VtK&�0�@��%+{F&�|�λ	��\��$�b�o��ߔ�+�@��ڵ?��D��יv����-�[_�<�UW�i���E��M�% �����j��������^�t�V˱D��۠�e�2���������h���H�ޔj�x��Nh��,m�f��]��	�l��é�֌�E�pL>�p\_���45�Y���%�"�z_�lI�	Ⱥ��$ �r�����w�.;����1����Z�S�U�h]9�ɻ�ev1�{��]6S��x ���R�kP�OX	-�_4`��
�ܣ�����r����� y#��V�q�H-Ur��<%��-�/�>�Q�M(���˼�_�/5�z��l�n��%�\�UZ�s�e�M���:��mz(j���,����=S�㺑R�MV�H(i�����������::j�8��'J���u��W�	aYD�*
ɨ�q_��q:َ�G�&KO:�Oc�s=��k�4 �"1�`�w�8�1�L\Y�	H3��t%\8̡�H}�k[â`"�σ�u�:�O=؉ R}�ݔ�3G(-keF�G�8�57�]YF#�G���l�;P�Q�o��#w���mUi����蔵P$8�9F����������-��8Ͽ���@4��/���N��)��H�����$$�m+�x��%�r@\W�d0��U��bp[E�cEL��
��6�k@�b�y�_�g�G\޲H��ț3-���(�?�ȃ�q�J��P�rU�@˝��D��}+)�<A1�^�=�q��\�q�e9]3�x Tup�A���~s��v���5���h��F\��sq�0kw�����k��ږB�u� '�K ����9c���j��X)�b�j�i�=P���-�����c���"��@Gh��SфA��Mj}@���ԕd?�!{Ë����:*���"�~xZ+iKbh4�}��5p=m��Rtl�I	U揟�I�g�}{��9�B�s�ă�GznL��L��֚y�v�t	M�g�Cmu�����\�X��-?7t2Hr� ����y\!s�՗���~�s�a=A�@q"H#��=�y����?,G-I�0�����%H��'��?�fd~��~կǤ�{�C4-��m^�0�J��� �;�62ˊ�����tV�ﺗ���&	�t�jh��ظ���I��6/!FQ:�n�
O5�7	��j+J&�������C��bgT\:�W3��*�K9����{mj4�$�kE��K�o��>����>�.n;&%4Ϫ���9�n`RI�>j;�O�P�U����@c��r!�y�ӅYt�U��&cz���"$A�������Xk���p�4PU0G�^�s3!^�&���e��f�㹳�U�"wLڗ��ȃ��O��r�hUEQ˰�s������&�b��|,��梼I�C1qc?|�����NJ8?G�6���T��6��˺������@���;��[f�������H�_���.�yU�/Җ�Y-~]g���uX<F� M�
�I�cd3m_o�z���n�tΣ_~p����6j�{��쇯F��1:(� ��RlP���x��,��C�"�<,�&d��J�C*��Ӄ�?������Zbʾ���ik��O��L���^��>���}6�i}h�X��Ъ�-��0V��<�����#1���q	ÁG�{S&���ڙ5>p3��8���^L=��$,ȓ�Cqw���?)���]Mw�D0�=_�sR�`ae����#�$�输,(ʝ�RH}��Q^��wu�yP�e���'=v�;]{L�� ���R��݆v7�r9}���a�ź����|�]V��$���@��I��!�,El�5�^ ��y��B_N	�+��X�g��Q)�O�d��C�$ɕ�i�U�s���L�$�R�o�үdE�6Ƿ�e���}j,G�$��8��Y��/�I�k�Y�G�Q�^rMH&o�<��Lc�r��i賻ҭ}t�$ϓeEŊW %�/�i}WU��~��\=��n��f���5�>c%egh�ѡޚ{k��ѽ��M��q�>���R۲�.�K�^*���Nk��:͠"b�ῳkQ�N�y�0晃�/x�QBi����!c(v����t9���L������7�KS��+��g#DL��ʀ�}�j���hA0���ɯ'��&8���v�$�ˬ�
��%!��!*i���,�TxV���:#��_�Uy(
I��G-
�#��)�)HQ�Q#T
Ø{��ˬ��ϴ�G�~���{���hi�gVߕ�'�.�(�[Z
����%����\8K7:��K�֟�X?%ĥӠDG/��5���ӷ�q�wZ�?�S�@DK q<�U;0ȡ�33�]ո|	k����H��5�00"���xr��T� �Ff�b��.�=��o�́��p��n����ؒBՐ����B�7<���J�/�(�҃��;��G�]v�w��� �A���Y�U����ޖa�w	Ű�\�x{4� j� ^D�ZdN8�M�_��Hړϩ+���x��-`:?���w��t��IU��X���8��:�6�i�8)Ԡ)�Ѷ��!��} �r�� ��와�w�G��될E� �k��h��z��O	�x�a>L�vMd��7�:��'�h���V�x��3YX��HF�l���� �Zq"
�Cy;NI�Uwq�ж�����ϭ�$i3����E�E8M�%�x>���S���(֐r�(����[m⟿)��X��!�M�y_��.!�RI��F�';��˲�&<�\��ٯd�}��3̖T�� �C���wQ�@���?�x�$�ǩ�j_h�����o�a1��_p�Q��-�x`��Z T�f�c��[�r1 :�Z���SԢ7M˴�aO6d���]�������',�g��`U��tzz���e�-�t]�%���?��������x���F�I=�V>^����`7��ݯM��|���w�R�1.4Rb6`w9����������}D��Fq�*k�:[^��,)�Yc�a�==�dbG���|s���U���׻qCP�9k�R��t��p,�˭���$ׂE�QH2:�Aɝ�E�9�dc���z�`�?z��]���,�)��߯���?!OV�._�dg�`*���V\@��}�*J!H{�UP�W��,Fⓛ�l9[�%�KQycfP�Oc�d9.�_�l��9@�_-O1.�~�z�����UҤqMH��w���[:��j�i��Hi��% ]
:HH�b��`���SEZ�Ë��w��	`gMu���뺎/$�̥7������P���p��ĕU�h5�#��\9���zK�0z�ddyc���;t�=�_���r����+��?^gw�m�kF$�λ�"r&\��1�ߋc�*��d��������q.�	\�ک�k3W�f�0߹kM�E_:3��TYc��Xg��C��;��ٌ\�m����
r�2[�Κ5Z�o�/��\���̘a�>�I�[I�� fXIm�q�e�j����q.>g%y�>[fP���.Â���jI���<ʶ�o	�7�=&���n>j�siZe^�3�	�G�x�y�_���0�@zōî�=y�u?ź�
'z[�$ )�z�`���� !���*��gLPG��'�|,����Ei��_/�\��X��2���"�2ŋ���p�(����E9�V9�}�͊MC�=�Bѱ�}"��Ta(`�l� ��6uߔtAbn)gS�&�	[q�r�)v��ꌆ���qfg?tUî3a8�����lYl�A�@�]YT=�$�c]����tu;xTOܙ�6bK)	=ӌ�H�O���B���;']��\-�%��6�&(�ql����Cs�9��&-��9�d���5fqq���NĩK��*Q��1A~��ܱ�9����U�a��О��z}_��<x`c���b�]\"8�v��}v��{�{4�2�
�6�G��+}��S�#�UE(�fa/s�����b֕K�pg��.�y~K;��o9��=a;��R����1,�z�*H
-I�:w*R�q�]K�cR$6�P�W�Z��f��K{�l�<���X�n��D��Pm�*oZ,zu+�C��y�'�9+�cY��)ަ/�"�ZPg��r/���׉^*�������8z�F�P�)���'�?W�p�y�ZJ��|��z����¶��2k��J�K�$F���4}7�@�Fäc�nw=�7Z�=m��ۢ�~�
e�����M�Jq��^��Er��Bkb*s�'��TfB�MSQ�~KjS^�����2L�}�: ��0�hû�m�g(� �u{�G���|�;!�B��������|ͅ��W��h���U���r0G�����*���Q�c��1+Բ��97,�Åݓ�o��u/wM����m)+�*�m�c��;�mTWŀ��Mo��i��Z�U��B��|��j:z�f7֛bK=c�H;�vX�
�z8<��򲺗���ix�M3�?�A�~%�Ɛ��l�ã>ckvITNɛ]j@�P~_�"��8�$
icQ����T�#e?��3�+'����yl=ʉU�k��p�s��u�UA	�|^rg=!ߙ͂L�z�P�[����A�,��þ�hu�[�w|}����_fN����!'�j��q@�E3����ʹ��I�����p��蛰5G��m�M�Y@�1hKH�x�w�kq�F�Jߧ���x�A��Y�S[������ȸ.��(�F��F�ɬGF@����1�~F~N�yS�p�)S���c�t���y۝!Y�*u,^N��qZl%o�k�ݡ05�9�ē��S�)���_|�r�� ��;�7�,���>h{߷)*��bMP���֤Cf�z#&���Z�x�C�*��b�(Z�H��Y�v�}�UX�_Y��F6MW�S0���L��hv��XU�uz�ϖ�'�q��n������q�W�|����>ر�(QS�Wz˨A��T(�qX�aϹq�aQe���9EӮl�6M{G���O���-�T�Pe&8�6uh�|�D ���-j�C[���XX��U	=,�nK6�Z�
�î`{��CY��֏ث�K^7m�H�A�h�CzģZ��/�>�1J��yT���f����o�b1��]Hp$�9��e�!��0k��ͣV���/+�K=�9�鵸��%�v����4����E��H��GL��}���4�:�h%����xw���}{r'�Q;����Ï^��"�)�����<���=WA�EęT�j�a��Zё ���ĜoWJv�ų=����w̀��%�L����<��w�͊ŀ���̘���ԫ&)+�oW��::��=�'1��U؅�at��(\���i�kB��3TE��"��֐�&��������1��:;|��/؏v��)�����g�j2��UJ��^���:P�f!��`y����X��g�	3ar_1f�&��Uz�y�U[��1�jBL�F�1�W�l�9}]Y ��(� 	�ؼW�U<P��')��H�Ȓr:�W*Ax��PT�:g�|��8 �|-F.!0S-�.�~԰f���$Ý�췌��m��Gni�7$�8�j���t����A�d������$W(g�K��/8�R������G=%��ٖŴ:��W#�I$$��ڿ"{�U��9d��P;\��>����� u�E�������c���RkT�7�	v�s6c_۟��K���_@���@P�.P3��@�
���g�ַ�RD���wس	(h>���q|������M�?:b��m5n�J��c�^1��?[.��d����%������L�@��#��7@.t�;�8��+��*��)�*�,�LFz�ݧ���l!���=� ������y����84���穻���L�[��N������f-�h_,D�I"3j�\��;�!�]"��Ŏ0����ԗ��z5�c6f�J���o��D�`~C�����9�ӺȪ�s��|!-\ݢ�����0�+ɶ�k�_�5*g��� �	�@��8�<�K�*a��T'��>p��9s[M'7P��nc�����;�i��<=c����v��T�_M�p�I���=�2��߇~���;h�T�NM;y��8�)p��K��4	�ǃ� ���yM���VZ��8�b�<��U'xSc4=}�M���K�q/ݰF���^���i�j�I62}4�kPG�'��O��:⎋���&�փpcUT�&���=���^�S�����Ij�&�Ҕ�:������>�"��M˹�����_�J_'pD�5�|U��l:OO ���w�'jk�eZ�I����,^M{�0�*����]᥃�
.M}���qہ�ME�aώ��꠾ݮ �69ME�c��L���s�ot�i�J���`�(]�ޗ�Tڞ��>~�]�M4���S�B�
TsH��6@��sCf�4��=��͸�Ӿ�[���:���q*>۪�	8����S-�i7{�O#���D\��J#k0:�.��U�-E���Z;˘k�B��E�{��%�7����Y�W�Q"a��l疸[��JT�O-��r����7쮓@��3��r8oB:����u�#��'�@B<�g��)���ز�ʌ�]Q$���Fo����>YˤǔM\CDOk�I��F.f~��6]����b&������P�DC���8��;���P]��26��Q�J���C]�t\ns�h�m ��&�o�{s����4���H#d��瞩�G�b���ӣ��F���%�j�X ��a��'�C]H�(��ޤKN	�+I����V�)먼\�ZG�s%0�&�Z�'*�7��Vķ��ɂ��n*��^6i�pZ�_��FR��.pٳ�L(Ik�d�����ʖNE���8�f��R��^����H��QVRG���)K�w#jm��l�"��J#�� �\݀葲�-�U�ğ�i��8:ݔޙ��}�~tz�{2cL��� 6�h��W�B�]k�:��a�XΝZ��s�T�;X�W+���G�a?�iQu4�Q�j���qp���l\��&^����H�u�����]'E �܌�Ӽ���D���͕a`Z[�[l,\'h"!x>�x��O��Ł�H3��/��=��ɛx����-Q��!V��[5��z�Mv�ٵ:>�ٙ��0��0`��qh��%����w�~W{��6�1���;R=d� &K�C&.qW{�sQ��j�eS��2�b�F��
�(MhA���_Bs��!��v.�G08�d-����a�������8gF+�
't6?o���j�C;����� K�ܟ�4B�m�OL'2����Fj%�l��J���m���������K6�Rr�p��1<,sy�#�L	M�sn���s�R�L��H|�)�ߏd��Ta2������|���(~7YG�p�-�.�PˎG���B����������8�����n+�.ZH��lГJ�(��v0!@��_%@Q���Iyi���D1��#:���)Ӄol�!;o�)k�9���9h�����|C6R��@��I!I�z��Ć&�Dq�����O�z�n[]K΢�I��w��vQ{^!+�Q��������5b,4v��]P��3I[��Ei����B�xJ/��}v�W�$}�7��F������'�j�`������e�V��2�Y2�����*�&D
*��@9�\qI���1����8��������o����M�	��U���&k���C�C�U�A��h�������x�.Ə���v�)?�!�!�U!ފ�/���R���b�ËU�ݶ�<��a�=v��j�#���u�y@���˒����hь���t�n%�FA��:����J�N���^�ח�3#R��.Jp�.J"I��b,
]��ѭ���FEA��I�a�贎�X�����z��/A[�Y�m��1�J�D�z�J7�v�ɛT��bho�c\��(
!]wg�l�yӓ0ٝO�����f�I�a�&P��݁_��n�ǜsY�ޑ�zKr��Z��pV�+�b�
A��5�K+ޝ��7K�#,,S�,�_��{,1�+@G��Ts�Zaa����FGW~�m}#��<p=�ۊ�ye�C�&M� $�ש�m%KSۧ�TD�\@��;�� �̂�!*d'�{����P߹F�f#2_7�-F[�7.]� �B�~)�Tiϖ�����$���b�)��B���2�,,�z�Mfqr<��0��
�־=UI����9�(��t��\ye���`����{/ku΍�</�ȉ�L��$h�f�IV�'���y�Ħ��*�o�+�/ }H�n��8��qB�m���w�y��|���(%oC@Ttn�`LZ�p{�~S��D*�W�dƗ��\f��~7�ԑ8 ��F�:�^�2ڼ��;�,���H�,����7@�-��VS5U���uϐ`�	/xΘ=�TDl����c�$��t<~3��L���i���u�#;�N{"C	��K��B3s�`�9�d�/X�f���{�-��	M|��$LrS��ͻ���V�o�3��h�fļT�V�-����P�3D;�,�	}~�.j:f�a��z�#~�&��B�^��mj����U���KV�L���h���ƿt��7�u�D�s	�В��r�����o܍RŦ��X����+����r|6��f}Jes����-5���l���3VL�Ubf��9@�H�q�X$7��Ȓ���n���5߀CZT��O��P8�r�t�,�^��\�U0�ϱ̩E	�[wEjإz�1Q\�҆��F1�*��pY՗��*��#=�%~9�)�-?��RM��핳G�$f����s�/<�_5w<�]�������m�;�VJ�d�t�[U�=��_��	?�ί����=7�x���*q���{�٘�CčY�i���=Ė<��Ȯ�!���U������q<E)�]��*��gs�����HdFl����@٤�q\@2E�2 ��d�������v�B�W��_�^�e�Y��;����8�>Q3~P��J9=0�-z���͂r�ȡS����:,�!����δ�K��'��K����w_�%�H�j�$kw�p*L|)�ѹ�xU�&�B¥f�6��R�f��[|��8��>U��(�N�|���3�!Rq˖e��H�߯�� �����1�ǀ2�Q�֣ғꡁ6u�mT��K��z6�CtS�I �磏��Q����s��W�J܅���?L;�LN��Q�@��^�8�x�P7rݼY*ߕ��ʴy�����c�/�P�m����"�Đ���1��j��X*=oK�rڻ	��zw���]WL܃��3n	�ڰ�d�u~���H�X���R�⾖��·��M�yIh;���oLG���y7�V[�
ОUiM6|�N6bv�l������ϗ�.BZ����6n]�D=R�Wm���X#aK���D;�r�����0M��͠���t�ϒ��V7D)��<�4�i���4�*���c�U�쥿r�D
Q?�-�W�M�ֽ�3y��Bt����d�3��װߠ�G&�7�~;ю��,r���8�2p�YUnZQ.)�3H��&\�L��q;J��9C2V^,V�ӁX#�8+�?+�'#���?�L���ګ�¹��{f�6-Ê����>��G�Ҥb���{�]O�I�@�\�OkwN��Y\a�5���9@��Ɂ?��q~B>1�\�(�'u-� �Ӏ��A�0���ɦ*�r6��ŵxJ"��{�f�k�yf�!o�Q�7YM�U8��pk�H$V��<��@��P=�w�4�@�&
�<BA�Z����Չ�����΋�4�Qc@erNa�{���d��z�6�mlE�H����x���hf�
��,�~+��+U,��z;>���=7޶23SQ�r�ıa�! �a�v�U�%�`�=K�{��L��r�w� XʅJC��1'*��u+�I"���I\�������W�P�N��27�t. t��iU��[�'��i��S����}y����S���I¥�
�Ur����Z��m�E�8)a��~#`�m9U��	nx\ &��#`��q#-�"%��J�+�2֍m���r�t�@�l<˔Gq�6d_�⾟$LX��Á�F�Z9�A�lW� ��Zx���� ��BB9G��)�\qļL�
um��X�Zՙ��_
�7�x!\p�Ùj��^���G |��z���um�m̌$��;�6*�@2��'z�o�)��[���J*%�w֦�*>q��A�H�ҵ��~4ϟ����E���CA���-�6f�.��˒�weΖ/4S��X����􈀂��p7��C��g��r¨�R"��[Q����z�=��m�Kf�#�\Eԭ�v0�V����.훓��Y��B���a���Zts�N��ǔ�+��
!%��?=Ob1T�H�:X�̨�+�!��	�pH@KNY�zh/��A���W��L�Vc��ǫ �\�֮k�ܮ_,� ����
�l�� 7�x!tU�C�YjY����h�S᎝'�1H���Yw5�XlT(��#�G�-��x�eA�[B`��x��s�D���h�J�o�8��Ɉ42�@@��R�YO�xM4u���{m~�,�p���B!����U>I�׆?��5��!�1��G�*@$5$�ԃz"��P�(`聝����WpL�Ni\F�Fq4���tf�� ^�g\"�
1+^rlp�|�x��^(p�nd+���U�(��h��{-K��U����@�}��?�k���=�����={X' ��`��L�s��"��ϥ�"�p{��P��s_e�F�D�<J7jC����q>�q�C�5����
n�	�HxY���$�l=����s�H���|&�W�,\�Hb��)2r�_N�ŭ��zt���9,�m�\xtɟi?a
#�͊���!����h	 @�{��jn����%�#G�]��C1�o��Q��^�[�x"�u�T[�A����M����nG�KD����kw�s��j��DR�(i��0�.��bU������j��X?���:����#3�X�!xh,'��?l�s��D+i
�=��]��Hdzx�� �IK-�ia�/y��Hq���u�0�;,�;�9Q����<�(��/��ή��3"�_	�	Vu�w���h�Y���s�A�<�����r�����Y�����x��R��s�A�4Py��W
Y�Q�_��׌?x�hy;\�� ��%wjwl�]�v��S�3i� �������<,����x� �2@e� �Ê!�'���T'���Ǟzzq�|�]�	͉��,�f���U:�d>m�73aDn��\�������wD�ü�ſ���y�	x������X��T�5E��T�p���ji(�H|�f��p���	K�u5?Ιv��F�f]'�"D���G^�(R曕��0\�ѣb���L)��p��]�4Iݿ�U�ӧ\�5�0��|�Dv���b�R@�o�r&�
Z%~"Q�]�滹̼��U�[`D�!��cb)oU���t8�ڤ��F�N��-���*f�(�"ot�����xp�dH{��MR�O���#��Py4���;*\�(iz& �!�,�E�t�eC����������A���c8���Q��8&��lu`�S�BH�*z"Al�(h���Ģ8��}9���U�]C��t���X����W�z�(��uq�gn��x;��9H�0�`k��n}��<C�$[��E,��D4Ch��N��o�7[�O�9cܕ�"��N�k!8Ѣeh$dJ��g�s��ZC?z�c<�ذ.��G+K����RL;_�)�?(k��gc�9]���n����L�-�@��*��:ߧbB���\��+E_PZ��Ǝ��[nI��=��%�#�A�ytY*��>��(��V�d�	U����fa�!J�]Y��C�Oɘ4���څeh��R�5%�"C�_�8(r��P7'b�@c���oE#ߛ��l����������8�>�� 
�^�e�� ���"�)�>�X�,|J�T:�����hT�%�=]�W��-��AI��X�v8H�4[�u@��\$JIᴱp+!RN(xv�ǲv�bP�s~�Ȃ��;�f�:9e��\��߅Y�WB�>���|�CSF(�wBY��і��^�=ӆ���	�
�O����CJ�S����>�L-3o$�0�Ǐ��iǤf�^a�PN2��ڢi-�i'g�-Y�]�n<�xv��0�CW�+e�(l�۱���%x=,���q`V	G��*�d����W��R��IF��x@�Xqg�P�EgH���c�z��.E ���c��޿��g�^�}Gl���_"��9C���w[�T��p��j�ǏKZ~E����O8��|08��I������"�j��-Bf՟<��ʯs�QA?��(�Sکi�%�$?A�ekK��h��`Z
2�p�^�w}�/�Y9�/��ٸ�۰��ii/�'�`w��$'��>�l<�W��-QP�K�x�g1]�7˦w�I�;_t���Β�ջ"�_�B��I���/�!ᝍZ~ԍ+m��4�V�P^Gi�nw^<D�?��c���}��Ә[���|�f�����._Ad�0��Y��Pl��uVO9��R&/�iA��lڥ�fS�ӳ�d%���E��Pxʂs%1��\QIÞ��!�(��cK�9lYM��	Gs���I�{�Ҽ���Hy�]Ȃ���?X,l�n5�U٨T|p^���z���`L��?�UZ+U�R�g��*YS�ҽ��K�{6����LJ�����';=�D��q��E9�S3iY�q�(���.����[�)�h��&�t����3����d5P�2(��f,��5J�RY�Y����0�:��h��|5�4�_�ø�E�- �~�s�z�q��7!�aM�i[�{b%�A�[�8��	�r���m�Vm�Wd�/��iK �����z ��x.Rq���%
=`�֐Ʒ��}����4͏�ے?	W�ݨ��(��a��S�% �[P����s�����h��&nO�q5ʎ� p�w�ZY�e��xУPF3�+�m���yuo��n��戉|���+=�zE�7;v�iq���!Q����n+%~f ?]����1T<�2��P�i�'�����{����g��*wU�����q����U3�vc�oo��-x����e�F�u�hg�#��A��.f�5���2RQ
gR���m�%���<Z��_	\垳*��/^@ȉv0�ԷS�A���v97Q����n4�ϩ���ΖY�lr���!������K�<#�w�Q&��w��/#�]�G״[U{�aŴ;�39V���`�� n����h�fD�}�`���Ƀ�����m���&j5��R�p:X�p�%eH�+�V�\?s�3��{��A����Q�mM�bI�ӻv��	����A(i����?�rvwN�J��O�R����4M� �8�@�?�D؇hK��;r�e|�F���s,�ʟY��ަ_��תJ7藈ʵ�3,}�-{�I����rc��`	����M�O�2[8QY��T7���%�
��@e�m|�]!	�~��/;����Pc�o^��C��_T����Z�$�`U*�^�T�1�e��{)�vw�2�J&�:ºdD{Y��a�-:�..Z��0g�w[j�(E�2@b{p���,أD'��r�+�6F*���|�vV�� �mh>�ë�$�]K�O�*�ք���ݬ�2��ܖC�	��HO�NG�{6�!A�D����N7`�QY�D��������[B"0W��-J��W�)��xQ�M�ٝ���0b�?����E�e�Q�����4�<������vzbMg�-�j����U�*8�"e���_��qD�7��fTm��kg��E�L�=�'X���`��}�gw�8���C�����U��Odʡ�҂�k�	!�oW@�'�颖�PO*�����pP����J��Ó~Ҿ�z��&���Q~vڲ'T���{`��L����3q�0�����ĺQ�3�W�p(}	u�qB)pF7Z(�J��F;��Z�.T1AUN^����"�OGX������-�LM��d���z�Ս<!�� ��Q)���I�,X�t֧:���	�L������҇�\Wp�y3�vT	�Xu��������م�U��%�R=�������*x�YJ�A�qk+��jYMI��:.TWODpސ�Z�8�Rެ+{��zfA�@���pYiT����Q1|�)	�DFD�R���W|���j�F���9��\g��u@�T^��z�i��QL��h���%��}�c�a)�|7T��I�{�z�X�G�k	���m�6��g^�y?�)K�1���yѬ�^,i��:<o�5�$V��#Z�/�Z����e�X�9�3')��L�l��I�YF�m42�5�.����)����[�{PM8�5l�{� ��Vϡ������v��>����x�$nz�b�v�-pnL�����1k���������=(��� r�7!���V��Xc(���Z�	����.@j$W��Yq�c�,6�P���K��Z��?�m�7H>ņ��ǵ�>q�0�`nyt�J��*�a� �C��A�}�M2��`fN��s4F���������s��)vy�������ٚ9�0���q~ϬD9ZՏ�y�־���\l��N.���6���������WF�R�ā�CN2��*y+�͊��etL1��DqLv16�ʖpZ}L�$�?O����Z!dw��Z�/שw%� ����t�K�g]Z�!��},P:�N�4�@>���'!�l'�Yu��-;(nK9K�	W;���=U$���2��\�����W7V�0M�)_���a�B�<}
�e�Ž�5�iY��ƾDm��������0f�,P�b�"#��g{��%�� 7���&:t0�"b��&8�l�T[����X�7��]ʃ���g��	�P�*�/���Ҏɒ	���0���s�8���*{�3Dz�ԫ6�[����.�\ch��B��"��O0�_�r9MM;M�{:�l��N!��\��pi���ݧ�ӦLЗ��pym�����.���7��C��D�D1�&U�9v'<�����j�F%���Nm=��>����?=_�P�[Ko�3rc�ehݵz<���VM�o,�1��?u_eÈ�	��'��·�|��,H���Yj?z� �T��A�@�U���.[e^��������;Y�x֋]Ԕd���{`�br�^?�.��,j�M��\ !��I�^>�z�۵X�xr��(�ـf�rS����^�("�j�7^p\�0Џ�vQ'�LЪ�c�'q]��η���ŷkކ���=��#˄h����Z�hޥ.L,���/j��.5��AU���o	{��[�m�Q}��n��r���b*p�l�#���p�Zn1�]�����H����CrW�7��p_��^ {>�v��ɨ�V|����Ӯf7�'���P�D`�4��W��3"����l���â����A^t�W���o�/��kᦥ���VuO�`5�z����.����.bf��a&���ܘA"� �Q�ea�C�7�QW�V��`��u�3]%q~	ކ��Eٵ ��5�^������';��{s�ʄ�@(�����F�N2�"`���ԩ軕��Gd,r��2�{��\���OԐ���(Tug�諠�V�h�����\��,����S���B�����c������$��[w3p��1�$�*�ī!�%F�4"����Ob���?��E8�j̋L�!s��$
����f����fÒhL���v7S&�ǩ$UT^��f"(����eC��~{Aɯ�H����ֻ��	�?�6����+=�/4��4/18~��G� ���^�6�έ���M�gDu�O���D�]�ŗ�xW�׮LڶTA�E�Ϟ��+aƹ�hÅ
��Y��NUΡ������;�ͻ��P*�u�R���;lU��������{�(X#�����0g�����J#��V�fwx2��:{R�2p Y8���D	��
��*���$	^y'dv���p;u�D��tmV���^ckB[������#�8�2�A<�f��j7�<?j��84��|��r�T�#�)��P�.N~M���[8�3yJ���7� �W�PN�����k|�n~��!RGE����:Z����FI���0R���������*%(eq(��k�MKY��h����qlaT�� �e�fm�Z��I��B�^�T�u�V0%p�1�M}��_ÀF���Dś��ν����N��Z�#?w�.d��ቨ����G�8��nv�ˌE��/]1�N��AF���&��,wu@�\�����W�}}�]��;
����>�	���#���f�I�E0���YWJ�v�.G�AO�Q�r0ý�*�}��n�R��,	)s�<?rϼ��"�Kr&��z�s���	��S��.A}�o�_&�8�G-X×��Lg?�;�UvJ�!���fR�K_�ɰ
ZK�1�����<U���%�KO��X�?��Ѷ���*�A*z��'8P�s�� �G`��b�T���6�l�?�{�aY���W_������'α8���s�X��X��yׂ7 �U�7O���p��o�Dk[�RPWS
"^u{l�P�:kV��nM�dg�50�Չ�����`@4���r�b%�㣲�{���6�>�q�]#8�ݜgtN�R��E�p֙�)�b ���E�`��Hx۾~��͠\W8���p ��EUͩj<�;=�Ե��9���4C�T�ځ��L{��@-zNy�h�*<�ܽ �����b�ǧ��X�ύg�E�`�0	b����2
��R��b��۪���h�~�-IH0eeJ������C����xO{���C~Z��������3VX�5=�Ŝʞ��	�i��Hb�8:?�R󶄪T ~�8e@q�OR��pHn�,�I���b�kn�Ml�Gy����wF�!n2!nR\��oh�Z�%M�yey�`sW=��Q�G�r�%�Z�|��"kA�z���TnU.�2�{AFѠ�^pw+3��.�qO;u��KJ��-��b󃦷+Z�����A��i�Z��	�+d�00����CWю�|X1�++Luǃ-�%OST0��������#i̯|��Jm�&���R������V+6�&�G3��Nߊ5/��p�V��͆Iz[����'=F�'g,�jV���'CV�B�^ק�C��Gk^^@#�[��Tz88�6S�ZtYh�s�=kr՛1����g��+�p]_��i���ɕ��E���/Ky6�PQ ��w�1�o�<w�B]z�����Hİ#F#��c�����)����z��m���s�$F���+Lx\�1���	��	Ȉ9읠�l�LҪ�X��JT��d?�y5HL�
y�v�9�9��&�:����@k��2b�\��o�DF>kR�59�<��9�~�@�C���.��Uʤ7�GE��hЪTwk�]oZF_@OSv�fގ_���[�X[C@�Z�c�����ww��^$�>Ũ�����J�_�W87	7��)"ft�dZ�$��N���GUB���#A'���e=Ȥ���!w/����Dǜ��%�&E�(����?�,�RW�"�#y���|p�]]\Z.y�X�u	d���TU�N&aD�夨3J���Y�f��0���^��m��'�^���W�+�k������$Q2u�?�a�ʫ3ô�\e�k��E'�{��=� wA�5�����w�
���p��S>�?�ȝ�+;ǫuL��|�6f���)��erNU���a��5"�r�~�:�Т�D���HjW@o+x��P����3S�T�^>j�����ODUd%�T��C}�e&QG^��E����e���b��%<���<_�Y�����'�/TH�S���OU(�V�����b�hy�vik`�̙j��lR0&0�~��jXJ4s���A/C��@(�TgCU������u(�L�)�O#��\�N�1�ղ]��)2y�4}�I��,K������~��{�%��(-��qu	�J;J�Xt)�J��ݲ��9�C�Ś+\�}䭽;�bW������̀�`S����q�]MT��X�粲l�Ҡ�h�d�e:���5��4H�4KiH��!T�tY�"kh
5ymx
�����·�'e��>�N�ا�W���]��5q;��-�_s�+����|Q�Q<�*%w��,�Qpj��B�;��V��|gݶ�[P�b�m�M�'�eu����M�������w��с`��`���ҷЕ�q�Wn�~�>JW�n_`Pz��|Bo*���NR6� �����DJ|�BMd��d�@��ImO󨸎N����MIF <p.�m�L'����>�63C�(�
X�r�d�5��a�F�h�ز����&�
��;U3��'��&(��*��ȗ8����!F-��T4���a�h3۔�>��`��v8@Uسؑ<d3>��@ z�����,���Ts���[��۪_��Wޏ�t�5�<�=G,�e�r6
���턩�'��{c
&X,Rw�y�g�;��wI7�o���n8\�a�u\������Zq�����_C�Y��3�Saٌ��58�	j�0pn��A�e�c���%���2�'�!\�Պ�Z�h�xW���S>�r �:F�V*RRm[�f0��	��qe��lw�n�n��hV��~udW�4���6�W��uK1������@[B 5yԃ��A1Ϟ}^h����=��_�K�c� F�]�.Qrp{]�٩�T��<(���M���Hŧp�!�4˟<�c�5n���Q�JTa��}C��.��� V�JԎ����z(�%�o�/aYr7���$�&�X�3���)}����	P9&���}j�Y۾��0 �HT�V��~���J�~��4�	uv����M�����{m9OtJ�!Z!�/�\�U��͗B��͘�����:^p�-F���|gG�P�i�"�_��ż�G����x����ݔ�A�[OM��h;�#�fǨT�C�D�,\/��,O�(bC�1�/�8!w�|S"Km\D1�ŧ8^[G��>>���`*�M=�R�'s�4���m��6b����Π.�C� g���Ix&����o��g�4=0��Ɇ��*�#jn9EY'�@����i<��k�Y9��y�\-uh�P��, �dP\C�0Y�ڿiÂ҅�*)�⺥:�:W����9���[�/��� ��'V��Q�>�O�P�8�ʈ���ٖk���O
n�6 �f!�(D�V2��p�GS]�fW�:�`�1�P#�	�I�nN)��G
IB��b�ݦ|��mF�K6T>��Do��i��S5�%��e��f�������#ϭZU�ɌU}�o�w%�'_
~N6�	O\�u�q���T+I*��p�,^�������G��)��w{�
�)���11�Q^3�z��V?$ �h
rq��%1f�k�D8�Z��A.�&w�J�Q�p҈�Q'`Q���q�O�nt��D��?������V�����g����s�����T����iu��W+�A�*���/c:ɛ�Xn�cĿN��K5
�#���b}�-IN��8^�C����M(,`�,Ŋ���f���������h=??�w�"��dm�=��3\5�vԍ2�R�6��ʅK*�;P B�qc��>]D��5�[�:B����ЬI�q��EXCn�P��O$���}z�1���#ŎW�Eۉ�ٮʵ%�A�J�ik�/���(L�I�BTӆ_,	�z�B�7Dl��^��4S�*��?>���hǢ���ӛ{��ܶK ��pvX/��S!M��m����r����lvv58�����P�� ��{�\�.��5v�qt.�8�",+���F9>iAVNW �[5$�����f4憢)����u2$�?L��>�8I;5��Z'Z�h|�N���w7	M�`��LH!>��^5V�����!'2i��I_n����o�l���>R:,ܐ�վ���8x鶈pR<8�L,J�$�  �<����E�����2�i?�gHo&�r^�.�خ6y`�5r� '�l�+��I�ik�^����R�!A����b���[��"�X� Z��k��l]�s��,��92㜭��M�Ø�1I���JAN��{I�k���#�X��Ѻ��s#"#�&,�`�&1�����6NC�8��r���1,AT������Z�͘M�V� �%ߡn�U��Jw��C�Y�rF>��'��D��P�<8��G���X��"��t�q�y����s�	��X���!����j%v�b���qQ��8��;��XKQ�&C.A*(S��5K,��:�ukJ�6��uA+Bo��<��?�ע�ѯ�$�vk���U��8���;8�p1�.	!�nf���<�$am���5���Z�|rJ�|A�[��Y9J�#]��颶�M�"���1qWG�KÄ�O�R�/��r)�e�W`sE�OD���a|"֑h#�+��@��� �j>M^���ó�xy��V�G��:u�+M4�t<�+J]uЃ9D5^3�<�W�"��T�v�l�d}�Щ3��m��'�~0��;��vs�vjw��lQ�0�uZ���xx�v��L�#?�h��A�i�ǿ��������t�F��z�-�:;S>�M3��z��8�	$.�Sg4�����#�`tu�P����`ժ��ь�"V8�o��S�~�Q��?C�ʦ]m##RGTJQ�7[�x��2҃v�.�v������"�R�
(�����TY�Eݮ��$[��G�A1����ǐ0vӴi��G���!6�v�O��Fr1\!��5R�#�V\n𕼥4�P�o�\�i§��J[�5�� <[�}�	�z>�pbo�Pg����C����Q�9�U��\�r�6�P����Ͱ����ʑ!�̖��w��'�f���HW�w`!�j�9�t������zUs��1�����(EhK��lq��ԬpSD���Y��Ѵ��������jK�Y��2�F=0�t�!J�H�F�Ы�tU��  �d��F��UQ��I"��4���ė.й�e�#Z�DY�Y���?��&a��(�� �;)��m��ǦC����҇{נ;�X��s�i�'�<�z��:�Gee��#XkAm��G~��l\���Y~+�儦��Dw0��g�uz F�����P:2:<ɱD/�V�o���ޒ?��&M�L�RCA�����}Ԣ�Ʒ�oKY~���{�{��Ch��+�o����{�T3L#.�_�qX�L�ϓ2����%��+zS�Cb�f*���Ƈ��(l^PUi
��%�8i�!?v}w�vS��p	ӫ��a%��+{r^z���|q �C>��o�y�-��TL&NvBW��A�*��3T�]D�-.�n���~��8\� �IAd�o��k�j���y��>�IH4�y1`��6��X��2�>���֚_�Do4�%�lZ!u�I������[�U�2�`�mt�lR͹�z=$7`
6�Op�ƻ�k@o��r���p���� J�]��˃@oR����n�v
p�˱HȈyK-�:�*�YW��#��:; @A��>l�%����V���1�X�4��݊�O�ҍ��?����C�J����&�@�(��Bz�Pr�$N�_C7|I&NK���|�p_ �Y�B���.5��j�v�R�+���K4��jI��go��k�93s�+��`��ro��`[�H�G���b�$�ms�`�+�����}����/���ǥ�cϧ�@s��t��!,F�c'�p�j�{�!c`�9��Mb�8�X~�X N������p�`�����`av�a��Ī�M��i�5����p8���1�;{O�S#�N�#j���{�*(͆�ܲ�{ފ,_\^b%*Y>���0	��7�z�X�j�F���e�f����Sa��B�-���a9L��S� �S�9���t��%t�^p�ǿ��P�v@��S��"7Z�Ҫ��u"�L�B�9ŀ�F�׆��u�h}J�[����my�<�ހmpE�v�V�@�����YG��QFHb�9�'��O���B=!�לmu�����4��6�Hn�n��^�"'b:5���,jb�R����;�e��A�B@�R��.P8���>uК)���~n`�(��|�BTV�	�ty�"3�-��6�_3Qms0�!����	�$��Xv��0�)�	��닏�WL���KHW��й�������)���%�r}&z�q�P������V#F��=���]����w�Ą:�Lo��r'����ơ���
��.�+����w�����e ���u^��T�|�֋�>t��"mїq��i1�2��"M��=�:��g��/�b����1B l�F.��P��5�`]A�Q#k�IV�Ȝҟ��BVC�Nb�-��j?/��n\,�9}��P���D��:�iG�@�)���a�B'����,V��D �a�RvC��v�����񰛔>�Đ�5e��uR��ۨK�[�`xqVT��:杙_���h�D�f]t�����˧�:���$�ȣ9d�~	Q�@!���qi���A���ed}�{���Ha����e�7�~��s5�Lcg�*ܨ���j�}���F �6Yh��mƠZ�ç
ٰS�f�ݡk�3�'�+���"�rf�;]!�sǯ�㢒8����Q�mbSw�Y�B�q��kuЖ�{�a���lc4Z����<6wܴ���m�ej۞ԱDcb���
�^T#*;w}p���M�(Xi��;\����Bw��M8�_;~R��}���Vz�� �`��+|E��F<:]D o?�xC����QM��Ȁ�h�#k���-�f��#,�������PB���!3z>�;��SA1%��D�����d�xs���1�X�(���z�Dkw��S*��^�ݾ���[:\��w%bfϓQ�$&N]t����Կ��E&b��1)E#���I�]���z�z�+�{oK�-��O�M�x��F8;&uWo��?�M)͘	��(��gm�lR,�"�Ʈ��u3�1/��A���M�
�г	����/J����!	G�%()��#Y)��Us;�ϙ��W;G���m/� ��"�Dx��$5o՝���J�q������ܫ��P�蛠bi��Cn)-�r�.k��.��r�?�$Բ+f�"��ƛY�t��Nv{TX�X$Z�f?�T��M��=���#D� �r�%Xv�-x�CEX_X�P������kN����<	�W�ԉ�~NZ �4˴����Y��TՐf� wu�aט�LT��-�;�e��b�zj|�6Z�I-M�(m*�?N���lYb 6�Ӕjz����&��U[2�`G�H�"�ie��M�>����;���[��R�:�<���ح��"?��m\T�#.�C�
��EsEv	�_^1���/(�]�D�j��w����F%կ�1
�z�h�����DR<Xa{��1rᴟ��P���7n���]��Z���{��_#�t*>(�g�f*��t���D}$>#v�Q�ߖ8N�t���/�q0\��m��h�<�'w�d��/*��@cJ�h����ߗ��l�AvM?D'e�rE�T��_\��`G��AǕ})_>4Ɓ*:$Z2y��4tВ��Rc�	�]^����}�e&≆�6q�7[�a�[Z*���B�����A��ǿy;\�}��iW���1@��G�^䞋��/��?fk2����5`�w�w_A�KIl��NtP����t����Hu�e����C��h���������G*�1�����>�S�"+�.�� �0�7���ǀ�s�ah�Kt���g"v��*eDFXi�[�y�r��Ǎ�M�a�j�3X���_jiE3�fv7-���1�4 �9��v�+	;ֵ[�Ն���{��"�\[���x`L�P�j�����
W�Q�Y�*rU����ix1/�������g���B9��!���|�q��dV�-o��@��ځ�L �'���b�1p{J9E�/��k�F�C6�T���+=���@TOCW��%)?�>����sQ�?ғZ�	Wy~a�CASw�G�&臆I���]~��ݠ�@ͯ��)0g7�|��B�m�����Y2Ӡ���A�Z::�T�R%�j2��)���*�0u�Rj�ɘ�隥ˌd�WP����/	z�]��OE\�UI4���g�O�u��ǧj��-ds)�H�)7?K�&�$ª��1������l��?�t�+��k[��R��\.���ª\��+�)H�ɹ����,K����H�,��9�. N��eaI7��y���L߲^s(����ڣJ0D�ϣ����g2؊�r['/�d��� eu#d����ߗ��HM���%VC�S��"���&����_��A�$C���p!8QE��mVI���iY[�3���Y��7w��\{�S������sWR��1�#�{��c��,�;CZw5W9M��/��`����A� �&�� ��4[h���?9�}y%T)�����L���4}���65��K����y�`c}��#������c9Ⱦ���嶧#b(�L�?Dfe��'K0!U*S;�o�_F��FC�l�"E��mVC�e)�Θ}H��>*���M�	��Dh���J���ja�hV��N4H�v�y0pe��P�Mx����vlv��4u����.��� 8�sy�I���,�L=7��ޞ�۷i
8Vۍ�KW��ixFL�E�.L�X2�M��kS���1k;�C�v,,"����"N��ИY`���P0�{}ӽD��z=����J~�\l@�}�*�}��0�(����&#���wqW���9�
֞�.{�wo����	$��˾}Gqy=ӕ&Pd�KY����mV�g��^N�ٻ49��+[�w;�7^���21���ҳ1��Ӈw�܅�,�@���8m���l;]�t�iF!��t���&x�R�pZ=d֌oA�����IK�5?*�j%��4��Ь��+b\�k�K�i��ՙy��6�;_	s�m���S7�	���T<%�+�Ew�Bq�'������6!�Mߌ~{A#��9�/șW��Q��	�W:s�����S��7E\��:��aڥ{CsT�v�:�xKy��b�*4e�b
y�)���{�����_}��b�h󘩝���o����`x�����.�f��M&�d#�Q~�w���OVP�F�����J�[1@�)_����Ŝ8ߥaN�o�������(��O�q���0���ܓ `�\��s
��?h�����5U[ǏW �Yz]����XܸI��򜋜];s���n�-?�;C����C��kT���-��7�;#Rg���
ؓ�8@䖢 �/f�
B�"��lw����%:��J�׷OU��?����$[�(�i�1<q#����9lݶ�'�!��ɧ0;4�g�>�q�b�K�[�R���Z�u@(-�գ_�������-��w�2Ġz���~hBݥ�����8��H�w�=,��	����r�Q�N�fV�9�`�or���(T��s�����X����&�Ml�U�^=K�)�J+PC$՛�?<�Yp����eh6�[J�4�p��G��|_��?1�ٿy$�4U����J�� ��ŧ�w$7�KT�]�Y4h�!�y��	W�v��~6-5佀�6�-��Z}m7J	�|�)�ܝ��ge��7�A��cq���]�k1����˨�>%*l������g(�H.@��}��[-���fG@i��L8־(a���d}]�y̩�twK1�c咖��g�i��dH
�����/� ��1₉�8��D���d�M� 4Y�hgt�(xÿ�ki�h�;�t.����,Rʝޥ�ɭ�ŕ����cwT��- �$ʵ��!4
��*Nz���'����g�o��4�M1��N3��/q���}w�ȺD����Iڄ;�����2J�~����ӨKM�`�y��o���-u'e��v��� �>hNP�����L(��0-A�6�]�?@ͤ� ^���MF:un&�S:�eҗ�N<�K�U���X��?ngd���0"���ݰfI�J}�_z�����|S5l@u����1���t#y����r�5��ϴNI��l�a<ئ���ǗV@d��*i�{�@6�Y�)狐A��T��HFO�e�k��MN�XN P�ƃ;vY�s�`=D|�o�ҳ�Zt:ظ��D����ԅ���Q�s���~o�LPS�p�v���'C����U� � ~o�5&��т�e޸SJX(�RZK���=Q���"��ʨ���r�ڑ�'���� 9��N�}69�>ae<{�(�X�4~����,A�$pn�?�[پyn2�n	4��=�T8Ͱ]�T�����hf�m;��Ы�B)BY�N8	�n�G���Dgx���S�N�.j�%b
6V?��/�������Kσg�v
�o%�Y��/��~r�p2�^I�g��a�4M���t��-����=e��c�.Pa����g����PEb�8�����%�q��2�[]ۃ�x����[��*å�f��c�f�������g9�HN�{�����U�s=���;���c����p9��G����4b��].���V�</��9��)� �Hιs�T���P�+�>Jd�,��C�����}9�>(�W�rDo�#�i�*�@Ҟ���
{6���U��e�c��Q���׭���6 �۶˄��S��8�f��&#"�2�s91rh����lI���
��q����IY�\�T8���;���W� ��Js��#�ky���O����AMԗ)��>�$j��?��rl��
9|��H�>� ��'$�x�&	��M���-�p�k.a���k"2A[����"�7��(�gJh�{~i��rB����A?���(گ"��B�g�ګ��t�D�$�yb���d�7\�fߋ!�H��@�ܰT��HB�DM��1kh����U+i
b ��7�i!���$����L�͋g�о3��jrg�U��S�ZG"�l��S�����cI��V���+>�>�YƷc�-Nj�y�����#N������S��"��7�~X��
x��8������,��!sC��\�z}��x���(�� �\ߛ�~����\�	�y:�>%��ɋ�L�`񓉡�Ƞ��z�MZ��8�sW�/�qS�\/Q8@��4� I�0�`��c�p=�r��&,��j�^E4J/���~Q���
vkѬ$b����0)��c_"`���3����� 1�d(���{�@�	���S
�|�'=/� ��_r�P8pw���R�f3���Q��xdg^�%�&�߫�	K��i�����"�O&m��c�|�Ȍ�ӳKN�h���q\[
|M������}Z�����),��zgZ��h4���h�p�J@W��y��/u�I��3`�8�Ԯ�}_��TO�f����hU r��U���!�v��	��� ��SZW� �l�jk �B��:"e5ܤ�o0P���xA��h��D��L"S�M�o	Jl����N+5�'�0R���w^�ˬjW+B�����vV�ϦF�f��=�����@·�����d�gJ_#5�\���T�\uA�;�T��oT���UX�LD\5���b <���F�v���<H.��G��ȼWb����m�I����a�Б;O�ޢn�$d�AH�6	�������|q�S�����Z������e¨S4=d�l�%��E��
����W��o�
D���^*mʎp|D��O�M���B7,j<*�9��@I�5��4MX<C��t���CS{��n$=��񏈢4�Ž2������C޻c*����h��ȷrǗ�*�%}l-��&r*i&�+�s�Rq��[��g�t��S�R,ЅSn�^�"ߊL�i��
YIJ�|�NH$U4�u�V��$C��� �\ň�Ԧ�EǺ��$͏���N�7D�qu���o�v�~o�"��X
�ka��C��nd�w����J�L[Z0#s����R4�/�>����ۻ2%�b�06�;����Z���<+�� ���3Չ�#7-��Q����ȗ� 6��hŀ�;ʪK�W�UXp�|sY\�fl��y�#Ei���͖)B<n+erWd�b�m��)NO�[����ɅzI7b��*$i��7��b�6-0[owF�X�V�l��[i�Iΐ��V����HZ?�� �?t,�b#����(#��Q!-Q� �Pn��]�Z�"�51N�T����	#+ũ+G��b�8����_J�.�Xf�/`�,� >�b��W�v	�>��N#F\'�V��*�[v�$J�w/�7�V����G�Ր�1����oC��BR�n! �g�H�z��ȰҸV	֙�ޠ�\{+@�H4��7�0��-�'��,%�/�"�#2�A�q�u�9W�x�Y��4�0�����kJ3<��R���>�;|��\6�p����L�U�-V�@�W�����:��f
t�u_���x��v����_� �qQ�}��,�H/�.yF�٬��X�$ �g�J����?�o+,hUe+�k��l��3xn�� �:`H�]�A����}��u�T��nvQk�&�I���ȣa	v�=�Q�\�N�p��6p[ܚD!�>|�0���������)b�ö��(g�;�l��r+�g�b꾜-�*!���׿���Tr�& ǭ��j@R���h��L���<Q�����ƞO��<5�'�I�(u�x��v;�E���d���`z}f���d4�S	2�����)�2�o��d�|P��O�~@|�1�!��F�z��0���s46��8�� ���j�;jӑ-��N\��ǹ�?J]�&�d5���Y9\R.{�Bi��k�d�S�����Q[�4zQ�J��zj*!I���m0�W���W&��؛��e����"���\:1��_��Fr�vz�4r�ܸ4n�%i}g5���Z�(����T�IFoJ	����y�-ҹ�]S��>g���D����g�
�T��k�V��?����N�hj��9Q���DU��Z��^���1��F��ą�w��0�� �{�T�>=/��c��WT�#؁y���@UO��+J�5��B����
@N<i w�F(�5ѷ�g��Ԏ�w�$�,�Ry~m�5k�3�_.�f�鲻����9̝�=/U��D��z~��sc���`|i۔R��O��Z0Ww*G�`�Iٝ������X��̬|6I���k�3hh��T{@$��������W���Tk)��Y������Z�b�q��F�{c�L?� �xF��ľ�3�_�Sk�*��G�TzCr�M2�la�.��a�y�v��z˽}�X�E������r�\
N^��{6X���xa�ׇ�C(&���������`�\��$)NRx"(�����h��W��2�
y'�/�vn���X��b~�y�5��02���:c��zK�M��d���D�YH5J��4��6^�e���Q��Ij.��3Q�Ϭ��p/$�L��U ����$⹸��ʛ��S�NI�&�_��C���",��l�Rtu���u�Yzї��A� ]#g�ƹotn�֥���q�w�ܰѪ���@�G�D�C�+���;ą
��{U��s��4/pP��ڦA�
�%��>ݔ&�}mX�W^X&.섯�*^7�lI=���Dҷ>*�=@���74������t��lȓ#���km������yIp335���&$��z������@lh�="[s���P�Dc�k���u�(����#��j������=.-�������}iy+��{,���jm2�wkj���*N��_��6G5���eF��YN����Qb���UbnH��>���}Y��-�S�l�9�0�����ek����u\-��#�F����W�ˀ-��W)N�Z��o%o�FHb;UF�J�k7uq��X���p���q���=E������(�>ж{Cg�j��{i�w�[ЅQ�uςp�� s�P}Q�09��i	E��7e�%epR-�ZJq�6K?�2�@ABɠ8�ŽD
� ecY`O1��7���¼��=QhZϮ����<�.���Zz;:`-�:�c?�a2ZA)J(
�z"���N��ު/;�&<���/�A�qX"�����#�E�?xK ���HJ}㈸��xX���1�<�@iD��4��.1[��*vte�s�,.��ux§�d$|�q�~�D(�O�	�s�4q(�"�����{C��l�/.^4"'xE����p�GC;�w�����r<DH��Q*J!�VVk��Y��`,���X!|���6L��PH��=�,��VQ'����N8Y)w��ks{`���u��!��\¯E�h��@��V��&�΢ݿ�7�;��n�؜1�:&���8����S8g���1�jd�9g�gu���i<&�	n���̲�QsP�%��\%:t(�]ArG�f����=3�a*i;.��I�-�T���1���݂ܧ	h;��_P-��kqi�`;�W\wrѶ�g�o�0l�y�Ԟ�ᯟ���Oj���),!P����6���<�z/`�
/��C!�"�s׶�l��!i���p�|R��Ѯv	�〉���|���8U���LX
Ne�N�)p�-Xľtļ
���J�d�����N���od��+��g������Q��Q���8�x-��H�@�l�M�;(M}K*:	���h�W�2��B<C9��A���P㒻�k��U~+>�`�!��/?�.ҏB!�2� �i�����i�@>�s �S<kU��q~�OE�t}�ݭ[�Yqbh��[����.a�l�gQ�X^D��������;�l��d_�1T�KԂ�v�0&��}��������k���>7�3LD����M�G�.��!�����5��F���J�ko�Ry�e�K�I�W�L��ĵ�<����wp�� g.jkj�pW�LK]�xDg�v��CG��qviә>��8ѱǚ&�9P���)~X�I��!���k,�1h��=_&�%R�v�. �\�.(zC4��ܙA����0}�@p�!���wvv�Q�j2�����T-
ɆP���C)V*@��xλ2��D<7e�IO���Iq~V�A=��`���T�kg	#���K����j����� m�y�n���*D�Y��l��$�M�[W�UމhZ�Q�m�xe{ne�K?�a`����;\D%O�0��#\dμ1�zW�Ə�b��0�8���Vj4b"i����Y��U���n�Py�À��.T�X+,�����\I��9Lc.�������i�X������i�\�a�M['��hM]W͡�գכ��l�����=
��B�P��mA�Р�p��Ҷ�}�+¸Q����D��&,òTv&���'LBJ1��b��I]?�����!(8�d�}�.t���C5�ɣia_R���	�����SZf���E4N/ D�:�N�.0�͟�p��Eo�@��K��v����h�q�;{���Ų� �V��kV��,�hR3X���S<Ǽ���ö<��wQ&�">3S�H���CY�C���Ao���Ro���e�ͨ��,�f��W�9�=�<>"L���Z�'i�,���N�ڧȋ\4y���_��-��G�^%��vf�I��۴���HBik`+֑]ŦE�>���ÒE��G��櫫6uk�w1`+�J���%]�\~~-��a�r�D�j1�Z���)M��@�u�yW#H���\!���n酟:{f#�j/d�dL�`	��*�V w��:�N�F��ݰ����TzȰD!�d�-���5��?6��J�s����/&ol��8�
�sse�Q=��&[�����P�[�=܁��/�=��U�a7�?���ևO�yΊ�3iȈ.d�S�N��`�3ٷ��b���-���X}MwPBR=L�Mo��Y	 7b��x��*(Y2>��a����Ss/	YJ�������b�2��?@��he���!���>�>>�	���٪Y��3=�ͤ�]�P'0���Ig8�DAu���O�򏑨�!p���}"�����@�;=��X0�&.��k�Hw���M?�T��u�\ҙ	aȡ?~��xdN�Rx���+��%\�,، �-̪�q�tL�7�6F0}�3?�Q0��� f3�^$o��ބ����7�����4�2�g�ʆ�C/Q y������f(zʂ�60T�d�GٝF���>�ӛ4<��T�I�n/�K4�z���lx�
M��~���D%���O�FҦ��sɍCD��6�<��q����{m�0��»���x�Of_4�~��p��=6�R��)�ZߓAm�o<M��K\��{�i5��/
C���(�^��/>C�nCz1_�r��c0}�w�DB��C|�5�=h0D�Q�C��`���=��p��2�!I���+�*�����v�����z���;&x��y�	\�y3�<S\,��$Q�V�	�5{{�){����Y�R��z�шo�1�|=Y����T]�H���������-���z�En۟U�Ν���:F��S�V��i0�9��м�XRN�.:��˖KN��bXFHw����_�]�%���9 �Y��C6��@���Fc��@\�� �Q*\d�jh���I�_��xΩ�����ˁ/��`8��x�s�0ֵ҄��4��I��t��kK}B���ڼ�y{sPw��UH6��oh�C�n;�v$*����>=�YE42m�a�C�j��[�b'V�d5����;�2֟��@,����<���-�Q�_�4�7�ǵ��2���A��k��w �{�S8ū8�*�hF�򗬸��B4
�B�4B�,�b�;�H�Eɴ���[� �V���$�%{~148�$bM��X�')�����܆(VIH���Y��h�ٜև)��{�����������is����z2�[�2��P���m!d����f�I��D�5��u'�U>��r �E��g��u����NF��S���%=��ִk�a0 ��\��)K�]pѮ�W}����8�؉����8��+�w�2R�S��9�����fw�V@�c.�ց���+C���"��ަ^�&���l���J���~�t����PSp3B��.��a��U∗�H�_��w��W���퀘|b�?�n�?V�
\9`(�������P�ǻ_�CA�����"�g?�U���15�t��b���&�����YG��c"�W̧]\�w��m��Bpze��ˆ �� g���W�b��i@h�������ZLn�]Ϛ�j�+	��5�c�o�E5U"�c�C���_���F QB�{�#e��	Y���%ܐ���oތ۝�dɀ<r��y�*��R����xd|�r�����=���I��?&#����)�X)�b�5]�ᦏGw��wq��\렴v5)��	����=�+"O;]2a���5O)/��-�p����?Wy�D��_{cڷ�xf9ܲ��=gY�c� ��/Q���*��-��~c��/��vf���+��L�܃X��F�s��2 ���!�v�C�t��LDtXDa���U�
P�R�^k]�}zBB����r�&�b�.z��Ȇo�M�`�$+�<t��c�.Wi���F��W�ן���<�^�7X�t!��r[_�ڬ�s��$�G�z脔U&���ϔ~�4�)�K}���c�����q��S�����n�$�g�A�|]��-����yt�<�T����܃��޺�(�x&�ո�8h)�ѯ�B��X�@&�(�Vm7�vѝ�}D����LS�æ�\�w.^�������g�.Y'V���ḁx���v&���w����"f5F�:�@]��('���	�����%[���M���Sl�`	��y�*�%�|_G2պsxM�M�1��D�T�zR�R��<x}��f�~&�ӝ�_2��-���\�rC~Bt�ƘPxG�m�����G�32�d�h�w�)ߠ��&����I�=\��1����B�Ot�%5tn��2~���mdHn�ie�H M�i!�ѯmד��^���Pܝ���6���C���78�N������1X9k~�3�1�~(2_�j�\jM
M��a�2*���;���s��q��"gf�GcBz��`��F,�y� ;
�+�bqyC{�o�����޽p*��/J��j �	�׋ =�Wd�H�R�EmK�s���q

`�Aru���r&�������M<E�V�8E��4��V������0���#��V�ז�����:u���f��H9�]jK汞6
�p��Ti�Q]pd���>&B�ݻW���&�l�����L��L3��D=�1;����T��<�_[>5�Oy�V��k��I1^��ۭ�UIl�(7̎��{P���vt��^�f{*��v!b�>�ݓ;�)� �� {m7�Ts��Z>�wf(x�h`����d�/n�A��h����Y=�FT݄��������m��G�8.����;Я�B����3p�A4��R��'�U{�b�8�_�;I�*z>d�F{/u)k�/�`��c]�y
Qec��ݗ���Gp��[������#�Z�[��A,�!�B��.d}�����?c���W��.�zvD��Rʍ���jyL�s#C�l�{���f�r�d�E(1���T�ا]տs�Q�
n�a$���Kt$!W۟��Y��taT�Ea獈�>:J��,�.,��g��M��#11*{O�"xW�A\R��V/���V<eƽ�&T�L�0p���S�Vu���z²�H7���7�Rn���A�����&7�,/�'��!�%Y���e4yJ�=�(�p�K��}m�����5XG:�H�_[L�Ә���?�q.�p�
̖E̴���؆,V�.CΞ9�P�!�\X����"���]¢祈�ݍA@����exR���Ow�3��Ny���C
������ǼZ���2���(lZ�|5S�W�R08�\���E����9�Y���p7���Wyϩ�a1�ͅ��iJ����/��N�]򃺻%{u���}�Z��S��e�I��l�A��� ���҉m���k1���L&
7��齑��C郼k�VK\�]~E��j�sÑ�i�Ӗ�Ei��( P}}�7�E��c� W��v�E/��hE='e�~e�_�UX�s1�r;�أ,��7�ɧZ%���^#����_ӑs۳�(m ���B�x���|h��f�iFr��[h?�l�a<��V'I-ocVǉ��3ΝSG�Z�k����樬��M������#�O��.8 #�C��Q�V��=凜"���x:c��]bq�Z}��I���,_�V��Y�tz�����ߜՑٹji���r�Z;ǆm��dS����z�VB��pJ,4g~���X��]U�#~-��.m� \��c��Ԃ5�pR�K�r	��*��_�ÔBq{��pIu�(�[��':�>o]����=�d�/�֑��a�������Õe��|x���r�A?F0�[��F��ӃC�|��!�,'�����������n��F���z)���7ƔC�Ӝ��Ǫ`õztH�,�����Б�[�15j�"���E�z�zU��dв;3F�� Z���?�Js�=��e�R��;$���$ZM3yM�+���TF=�t���x�������s�@����Z�5�8�AF��u���C�Y�i�C%'>Ad�t�Ժ'L�c-�ϝ���iT��j�N�c�iy/��&Ҹ<?�Z�r�
2��C~� 	���/^�pM��~3*o����^1��5`)0�J�L/�j�2}QEO�=2 |�'�T�J�d���8�HȚ	�Ɏ(�6\	u���j~o[�6�a��o?@ ��f�/�9��>�>h2�`}z��>G3g�}p�˳FY,p����1�����W�b��q-��ZoF�� nx�G�0�x3RO&�騀�t�^[���,��X��y<Z��
u�:��T�����$���$�z~�:-�j�չB��ؑ��6��P��E��f��	4���u�}�)T} �c�yf�B>0\�OδO��ܝ�R���fw�P����CB�3�N˅l8�x���.�~�|)���D�H=$[%,�W=��L>x�z� �ͻڣ�ϳ�4��s
�A�%����m�Dkm����@�Nb�")�#���.���0�+�3Y�
9pG�X�#�22�wl��	cM��L��=g���)8VRK�����mEv�E�7���d�_�uc�s@���/�s�j$&l�S�CE%�ف�$�pE�'�l����~�TS�s��Pak�� ����� ��� ��%�.|8��!�[t7�C��C쭆�U����A�}r�LɅ��8�ToS��4���fL��1��z��p��,�m�ط�[��^�+�ͯ	�A���ۺ��n*�T�y����J5�~���Ӵ9��g��_��yh���Q�p�̪��ʔ���{�W��֨'+n	��K�p�Y��]��� �];�ϲߢ����ߺv��i�Zf�>�ק���YAf����4��-���(�
��3W�.�FFҺ2�6�ƚ���\/�a�PR�����T�V�	�(�q�W5p���I`rs9�)`|=N����p���Vw���ʵ�ck�\q3w���1AH�_��ځ��ڿT��m�[���ͣ�6�|;�~n��a~����#4 �"�^`���~�ޜ�8$ې��߱�rC�Ь	�^I�6Ȫ?�������b�z���V��tn9rϻ��R�u*e⓿�a�bL�O����C�(Ot��m���ʅ=7tuSVo��\5e��~����k�w���]|>�c��u\N���2���Or�կ�:A���y�{�VwU$�ǵ�mnM�����k4: 8Q��c��Wg�!���B����{R��S�}J��s�]@��0%�1f���{?@X��UY:MK�ŋ��,|�gX�]\|�c��j]���<�ۘ�4�ߥ�E��dݗ,�3��E�Υ' ��.w��Å�c�5���<!z����i�`.x��=|> w�tvy����&Tp����Q�d�r4d)��w�
�{�*!�'��RvY`�*���aNa�oA�����2�-��i����[s �X�l)�!�M�5]�l�>}z	��r� ��@�_��9BČ�mE��M�+�g)#)�\�l&�5�@]/M�<���	tLSѴ�����\�т�/���M�(̖@�����,�0eY"&�ƅqA���-��s���_R�V-���E��$������3�/q!�R�u�`0r���������v��䭼�g�J�'<lS��U�
��Z���(y�8\�] [��k�\ē=fƿ��u���'��]lv�t�vE�煍q�A���ä2�13%�7����-Ԃ�- )�M�&�9}���:����7�d���K��j<bZh8�'����`��Ǭ� �&D��U�1
J�0f6c���O��1b��ǿN�7�8�¡�d�.��T!<�p9QEx��i��,���^��u�:����󔳲�Dj*���Cө��
�@p�1�UO��M*Ҏ������1�c�����0mguV�s����2��w�b�W��7	�ns�g��l����D/�_�&��w`��2|[��0Z��͏�[�Ai��38����+}mms�-r��
�m܁fl�I�R�y���\=.��W^��FC��e=�z��7��	rDy����~���1�(>��Vr2Ta��-�op7���c��^��T�Я1m�J������=T�,�������~��Ś��Z��i�.G�<���c#�AewD� �|�����_�k��Y���7���L��'/�D��b3������Ņ���\򑜓w�mҶ6��8�4��y￀� �K��@�_�*rr�\}wY[��"�Ng�Ig���p�k�s�7$<�1&�/���t�E��趈��v|��ۜJ3�ۧG�v��+�h!{mv>����ŀ�m��M��a;���j��2��2T$�Υ�
�6t5�\#��k�s��J��=�U�Z�7�՘�z֧`��=�*����{������������ݭ@p�)����!C�b�&��7mt5�ۘd���2K�z,��e�]��X�:P�U���?KTXRq|����x��%j�mq?t�1K�A���w����eG�����'��V��ϵ71�o��>;��я9H��F���� �ڠV�7Ε`={M��ӫ���8���{������j���\�/��t8s	�-�64�Rh�l�ew}���@d]���-������L[qSX A�]�K�t�cǎ�0lk�,ŇMrW����&���1�g�\/+�� ��w/��/�AI��)m����,�:Ⱦߜ�ǧ����IK�qJ�Ǿv��S�������.W��^�MO�ld�H9X}O��f��ė���H�F����ݐ\�O�p�fˑ��� &�7�=F��ӷI��'?����|L�>�-�t�JH<���)S��s��b5����=���g���@b�̳0��Ȼ|2����/im��;~�����C�C";J�c���o�f���A���2�b��ɶd��$��8ɞ�-�	�qNO�k]���_�tAϧݕ���849fl^E��rD���m��CkK�>q�f(��\A���CPM!T��$�%��b:��+8�F�7��O�㙹��NU�)�g^$���̓1��y�O�F9�{�}�qڔK�hw<��F����ޢ_ �O��^e%)���E>��{aJ^�'�}=S3�&Q�K��t����`u���J���x�� �È�0C��e�E7�Y���ۣz�6�SHs��Gm��]�{ǐQ&,?���`rǰ��4�}��R�oAܭh�X}�,����.���B�r���wx��������:��]c.-�+Tk�����>c��3�3+�䉃���S\f���� SSZOT�%G���e?�����d-�'\�e�m��1�y3�	��;��4��|I�/�0�o)_���e7e���OLk��5�s9�{�8+6�Ld�7��#̺�K���5����x}��Z����tƁ���H*�uļ��:��ec��+#�� �-���k�.�3���3��d�.Y���%u��r��P���x�U�� ��
S-؝��V�5�80��Z���滛4���g��e%�>5 ��k^��^��'3Ғ[h�ZQf0�Z�������p��j� |J�i��ss
��0.�9���[ћ-�oeއL����u��)q�n�ҵ�/x��k~�L��-� ����޴9(f��E�0�Nek�A�[O�ww�����hR�TPY�:�$�`Hu܂,�����5����D���UO����n1�P)�j���^KZH:��fk
Pe?������%�����p �'<��"���94��#�$�;ݡ$�3�m��x -�/��T}y����*��OC���TĦU�b�d��R*-��T��
�f<��&��%��� ҽ��Q�ci�1�r����ϡ}�ې+�Qv�~��6{�]���	q5�Q���=��n�c��/m�='!�E�(�����Ƒ��9�w]x0EX@A���'�s�JI��ɳ!��'��n�+(����w��G�"�'�P]�z��l�d9�~h?��!W��~D�I��a�R��o2��S�`H$1W%~1~���O���3���� 䱐�]k6�SAW_�y��=u���q�pN+�d�Ղ�I;l�DAY��ҙ���xLڠ�~��nt�:U�ˊ�������	VG~i֔|�+r=b ���Ů�y)��&Q��2��{�)���d7ݲ'�Ea�E�x��C
<��x'44������V��q�(څ���G����pa�$̭ Oν�[��������g!�wuG�4)�D���)j7,X�H��*�y�I@N6 <�0ϛ�-b?*IR�W�tN��%�v������N4�޲���ߒ�����ޡ��m\JI7�e_&_|k�;q��):3�6���j�o
F#Kt\tAp��6m�Hb�;�7��Bv ��YB��:	 �_I�%)�;''ȥ�!�*6���hத|�A�%�"�p�+;�<��9����9�XݔůDrpv,b![e�)G���A��7y����+M�FAą�
eSO� ��E�?mhg����}g��>gl������W"�e��L�Jee~k�y�n�g��Î�ڈ��E�$
�4��o�0��J�sG��t��8g�59����ms����H��0�{�
��ȉ��bq��(sM�Tv��w����6�=f�؜�����ɨ���no�7�~�?|�Wg}���$�an7p��Y��n�N������F�3�o����j��C���қ��D���g���x��_���Xx���W���{���S��3V�@�����<-z�q�n������Mi��0�4Y.]��0EV2�B�G��� ��w��J��\����]���X�uۨ-b���G��	'����ŉ������T�r�t����j6��������a���y�g��rB~U
�����y\X-�k7Z5.��JR��`H�df��X�P4��Ĥ���JF?�� ��D	����;G�, ��?gDj>�M��hk�#t��p+ޙFZ9أ#:���E��$��C}��I7놪��:��xA�nL��o��9]ښ4��VIwiuf��R >ɘ`@ȿ��*U�|�'�ws,�i��q*��ٜ�~���g:�Ay���]ƴ孿�����.��j����p��m���`�
%��3Pp�S�7Fv)\�JSxV�Mν���gs�+3��������t�0����cm�0vbrxT�6ì.�!ֱ�����N�bn�xe�0Y4�؄, 0�C~@hc*���	Z�,ykeg M��>��qd�Y�Z��<N�#�!�~���Qb�L�.	��fU��Y�I���j^�p=�7�䲠�b�JV�:B�2X�F��)�D^���׫̀�6���l��sZ����o���^o��'�T�)�(����#���eR�?�P�(��r
���/�H_hEՆpg7@�X�O��ZV]����}E+��`N��X"9/�j�b8�S��S�]Na���~_���� �Zz��c$%|dt���o;$�3�5���R�&�T����:Z��v뚊��V��	T���h�}�ۂ���ѣ��H��؝���~�`u1����L�}�q=��|�5@k�c4��۷�Ӂ<}��ӯF�GR��6�\�(P�GlZ#2�� P��4�6�����P�n�`��!e�e��
t~`�(���9�#^�W�!�K��)�K$@�,��*�$U�c����eb!��-���� 2�F'KK5sE9v�-,����A�F����=V���Z���~/B���2?��}��e�����Ӷ𮎟A�����Qژ�8I�':�Ry��'���G$��})��x��0����\��t�V��J���rJ��H4<�u(Z���:��5O�\�g�8G����^I��Ŀ��	)~�/�Fi���ڵR$6�m��Z���0�C^�`�0���ьĨ-k�'�D�������$����Z��9�/;>�V��DAlB��H��qUì܏�H_���?��=����;� �A��ʳ�g���|5@Rvj|&:�nr'8�{-
���b��Bn�F��KT-U�[�����,eX���ݪ��|k]1E����c�s�[-�a�c^��G�F���#��_R�݆Ҿ��V~$���ہ�'@ /|y���G<��@��]��B�¤�H�([�/�L)Z	�h�G1��/b�Գ�;\���6�R�6�?�ք��V�)#�"��}�8 �B���o�c��p�5���~�˾��<y��+��j��4� /�
UzcL9��2JwL�1qgSfq{�Or��r�dcB�	L��U�++�fP�O;gq�����������{�{�����L'd6��&�p̨���y�ώH S��!�qT������Z���{���������R���7 &*3DA�C�<�|�.�H0) �V��Y�e�Oh���b�~:��c��~��w%59H���Lݪ����#����U�s�S �[1)�.��~���	-���+v��#Om͵�k�~`�H���I����\����;pr�w�k�嗪0U�
�Hd�`�l$C�A|yJ���q
e���,Jf�~����G�y�c<����3i�)�!#��d�A�OI��:r>u�<���l�Ws���X�kd�/`vj�G_p#x�M�����8��f�p�0�;E�D8#�:���Or\Fu��HGC}�íg9�/�̯�ރ�t�e_�}�����B|�_H�����	ݜj�@/_�f�$��>�itl��\/Ţ�$U1t����gIb���D&r�q7S��?ɷЧa���>�ǥ�f~Ҿu��Á\؀�ޏ���E�,iq$���k<�m�}���QDCu�.�`�KX8����1F�Y���I(;~�������/��ܧ≂����@�9�j� ��讑r�8h�B(K�a\۽q���[0��kֈ*by/Opߡ�\�}؝�YO/G�7�s渎��1�#���Y�b>S�ӓg��A�T��)O��&(I��VlS���{�ʃ<���b��$Ʒ�+�Ln�/d
���% � I6�A1�q;����2����@:�,�����kɯ���~^Q��8U>`y�:��� u>?=՚:]4JjI��a�����WS��W���J�3��G�ŋ*N�W����h�v������Od~7q�ҽJ��c�+�"{�Ч��'���/�)��aD���qhqqͻi����~���?u��fk[��t�o��r
)VRru�Y��l�;�HH���i�p�ȇcs]�����Ƨ�+�V(��	"6����*�JW��=Tm�b�.��7 hS�~��ʆL�ү��є��{�R.V��s���fU ^�`�����~w�S�1���,Y��/f��5�S�����8�zZ~Ӎ�	�x�?�Ut<� ��^A�q�rg��������K��J��+���[���iK��%�4Fa�T����u��S�������@6�W=-S��q3}� ��]��KA[|�v�cц'���Ovr�!Ⱦs�љ�1{M�P3U׼�Y,�෿wԺ��Wz���h�����;����h|5GvRL��j�LM�}����-;!�pkg2@��>&���v��^���=��l�6�M&Q��ِ��5|m�J@"7�����zv�|p��D�[�q��Np:��Z_���$�6��K�F���9���ܷ�@r���K��gJ쫸w[~�����cwK�$��Յ�R����w�Q�יb�U�/U���y�s�f��=������fC�XS?㘫�{�䗬�Yp�'�4�1�IFh��0=<{���PmAt6C�^��9������OĚN;���1�"ː�eV�Q���=���;�	}d�=7"�*a�@c�
�������� 	j�>5�6��QfT!�r�̆ ��ڂ1�i��D4^���c37b��8�K�.��t:�����r���e-��<�x��`�z�H?����K����G��q=�1��Q�����rMm�����4]ke�	���8�ގ���BmQs#)�	�a;�AΥ�d� *�N#���k#��u���2T�Z��ZGy1��I����)qʣ��@�7՗s#3���ݴ̣�И�bIz�ݍ��� *k�^xv�}2�N���E�{'TE�rQHci��֜�C�5a%�i�9�u���ɖ�(�8/&E���հ��e�c��G����6!�(�t�k�u��eHֽ�����.4��+���ImnķA��o9�u^ш�,��F{D�"eO�$V0�$�����l{=�5��.�єx,��~-� 0�/��-�C�!)�5�,����A5~��͕�y�E���61-�5�����`4���G����>bV�.C�ī���]j ;l	�k*����t:�`	�P׆�&wPU��:iց�&�6
�#IT,1�zf���.{��/�
!§�J4j��C�رW7���#�[��֓��#��y�v���ݖ�O:���UA {}��wǹw�� �XGŀx���P{�-��$�����8;��Qa�6����_���3�ԜN�;*B�WO`��y:&���pX<jS7>�ʺ��u���%�x�p���P��ع��#E�Ϣ��y�����I~�=�����*����W<B�x��݌�=��g�-|+������Sl�ӈ5�P�� Y=V���H�M�Dc����k5D-��ʊ���@��&������Y3,I�R@� �m�@��y��B�S����O��8?hńυ���+֒�V����<u!�Z������Kh�e���`m"�#���Q�>���_�>S�vz�~Rx���U(j#lБvh=�(�t_i���B]���{�S���L�+����Փ�SB���!C�)W��Q��3�1�Qn�ޕ1߯�9i#��g?$��"J��±_�������W�kFN-
6��kO��B;�-H['Ɍy��q�05��ƭB���j�:��"�=��?�ţ�$>~?T0K� Y=16�w�D�� ���#�5	
_i�o�QqBb�8%o�G�S
捞(xv,��ݛ���UQ�b-��w�zu�70_KU��=�#�W斫;�}��9�k7��4�SI��E(����}��V���P9
�e���3�f�g�]�[��q<n���3�v/�Mk#^Y#7Sc}ߙ'�ϗ|a�QE޷��D�E��7@�[�Y�V|�mW��l	���*��<���8uO�����QĦ�����ӉyЏ����R��j�r�������ݥ��{]����7f����~�01�Fk<�TԔ��TR�3�'��a�q���0tL腽��O�WLcU*Ż��$�5#�:|[�8�q�?YfB)�\,0Cc[	��fu2��b=;[@YQ23���)H���ڮ�ʭ����F\�A��q�C�8y����� -��Yv>�x�]t��US�R:��Ie�;CD���\;Û>����EM� �O�rlD"J����^�gX�m�*4�.��h���?Ճ��FI�"�s��4��Ezs�cn���h|IHB�dm�[�)�p�h��,U��&��A�Ja�q�^�X�=&eH�^����}�+�[���joV��g�D�|@���L^�ƀ̠U�pi-o���p�:,B������̠��5'F\k��l휽���_��Ǹ�������<���&ק׷�9�y��XA�~.�b�[��n+�?lÂ��Nm��O8��Ar��JJVS�|�M郓�
 c+�I�<v��h��'Q�Mbls�֊AL��:���m���_��S��u�Ί~��' �#�'*���#"�.�aBኁ�B�w��!O��WXH�wBS�=-�9c6k��(4Nu#���[�(o�$g�mNw��Hhq������ ����!^m�Y���)���vɣ�白f�������}�η��5�ړ�O���k*�E�)�tf���V86�sp�k����Pɣu���]����&��;�&��Nձ��a�l�;i��R0�>�?Ȧ�x0�GS�����؂��B�x��[��|1x�XhAaN'��f`�Mb �e6����ъ$�`&&H3+m��g��ՠ5�)�(��i�o�)��@���֏?��}�t�pz��k��S�˛������I���Ծ���}���<�o?��&�t��3g��'�!E�]A���	��ЋQ�l��9�,��L� ��q[X@{�H"L�&��<y���c�GE���~3���_j���j �m2������并H�*�1�p堪�����o��,��NӴP]z;P���zS�X�9���O�}�+H��Ҳ8��ɕ�!LO�������̄�΄d��̯R��@�r��f�C*K _JW�5��b��Cמx�7�\w%���3C�A��@H��`O��ĽAGr~�Y�;":U'B;0K��3�Qʄ�D�at�x�2y`�y�kVbB��ǡ���He��Y������g�����}�{cM~%��� 3�h9"�i��bɛ���S"⸮i�4a���;�V�yJ�	΋&����R��.�e���Y h��D��(����m���Jw��_h��_Y�벛ɾ����.#�ȂS����|[Bx� ~6Xɧ��E���y��̖�����Υ幻�����aSQ���x+��_<�y��Ľ�)����G������P�d������Wԇs�z<�8Qº�@�1��%�;e�=~,(�J�D�O{};@�kl���>�s
�Z9F:ŕԲ���!�x�&���='�Sp�qÄ�Eڱ��F�C`9����3��6����;���ɧ�zu~�W_�'+p����~E

:*�]�²�2���C�jEQ�ĸ�%?��;,_�^m�m�W��K��+~�UD#�y�l9w�C��bo�wEA'|�m�Z!�in�������s��91.:|�[��b%�ܜɼ��ubt��Ϩ�E��"��~/M8=
Djr���	;�v�C,�z}`L�4�~�������#b������[ÆU��>��h�}5�fM�[�a��F{�g4
���@�W�����]����sNKBe17T�]���4<tz���^�׷��w�4�O�:��ğ��=��?|-����C�@j��s͹ oa$S�ER.�b���q�Ѹ-��;�%�d�	p�BV~ZDƦ`��7Z���K�E^	J��bx{[��_6a�ƺ�8�_ٽ	BEDw�vG�L��o��3���ul�,{2��#���Z��i�����#�;���;�O0M]#��H�SF(�88�f����j�r��5I�W0�lM"��+L��q�׍��h�ÖZ㢕jHm���eF�ܾz�%��ÀH�3@��Y�2?F�:�h_y�X�BʵAr]nĉl.t��V� �f��E��D��1Õ���tr��^{�UD��=*K�J ���N:����H9'~�-���{���лT���-1S����w�J��,�/n:�$��L�4�>g�H��=��}���
�탠��"����L
U��tw;4WUڴɮ,F3��+�1�zJB����'�-<7R�N����+�_jt�Zk���%6 ^p;]r���j\��;�_u^f`C�L������T�j�R
�.Y�5(���5���?C��\\�8��o��;�a���ߡ�=�m�",��}��V5�N�e|P�':��sZ_�P��*�(���^�;�-DT��L�}�N5�Je�\m����������⣷i�'c!h�$'���b�pGN��܍Ngzk|�ױ����F�I`VŖ?S�Hӌ�Πz���e0������H���tp���Pn.^����q3��z=J �Z�� p�\�]�e��}I����?`|�"%^)��UW�}'��E�+o6%�>S\�tR�ٗ[����~�ަ���Ț7HNv%�TĢNΜ։z�i��@��_�1����{ؒ�AD˻�_�\>xTCL%7x�SԔ�d6$�o�����*���P��\b��b�M�:L�Az.�7��ң�3�o�m!z��v8�-<�q���7�}n)Eg^�s;g�{8����J�h��o\�9a��"����1�.�9����7�y_��=���*y[����k���f��(ܝ�ځE��f�_l��J���LYY�d8��A��\_�ƁK��$�*�j��dEi$��.]�2ǔz��Zj�b�i�@����fM�6r�@<{� ¿[�;�j�x~*�`�NV�y�li�L��/��#ǰ7=㜔��8�{�ڝ-1���`���u�v�%Q"x��D��5��Gf�4^E�G�~�^�}c;ut��I�F?;w��LKv�c�o�K�h����Un���Q����?��kl�Ǩ���$~m~Z^� 
��3���X��г_�$")xr���fAx	��/��L�O6\ʻ�ޫ�����R��+����J �Y�\8Y�WN8����cp����d����:�������Ǿ�o̹������+��8�,n��+�ۓ��V��J���,�7����`�6!L&W�!u�}x�W���Y���1vM�	�K�N�ūз6�uv�����#b�-PE���|�HчJPş�c�=�Z�x�0%��c{)�͖'HΓ<T4V�F�He��Ae<	"�-�R�1�0�.PL#���Aֺ��`�6��g�F@�pW�Sb�0��4Za����L$w���h��|��g��`��1�������? �{�Nan���!:�F_�;��¤��r�Fت����G0��T�v)^q�¼1 i�vg��XV6��#��9��)R��Y?ܻ}���ߠ����R���/,��v�E�r��cQg��s��j�Q*:�z��L�n��,Ӽ}��B�/T�V�8��#U�V�ȷ${*��ے�?DOu���m�@_z�S.l�ʝ��2>ݐ�,)!����E#��Vn�l�@��Ĝ�jN֗��nH9��(�հt}!�B;���Ƃ�_&a|9l�]��*��S�QcH�'|4��h���I6!̿H�hC���up�中E���h�^���yw�͡p��q�9�&��2�C?��Vf�� b�}�A�}Q��:�& M�1���|�}l�SJM+��y�@"�l�U�`l)�\R4�u�>����T��5�� =�lA��Jq�l�!�av��B�����mj&��9�Y�e ���"�tXͤ�5���N�>��{�Qn*�&hI����ۺ^[�q�-?��H��7�4Z`,����V_��}e8�>���������+�n��)�D^��|$�`d������M�����Q[�$EV#�ʇ������"�[SDg���{n���h�gf���>��%$SK��q@�L����0������
�D�2��CZhg�^a�Q`6�i�ρ�o^(��vH���C��6�"l���7�����D�*ƫ��u��D��5_����껇̪�3\��H���b*���A~܃� ���/)��gǽ���:L�ܢ?M�л�|������T�r��ǔa4��J�V�)]9j{o��=6�?Z'��!�y�Eʕ܈O}���}���i�9���7T��	D>6�7��/![u�����^v/ߤ I� !c���#r�I�!i2���▾�O��M���i��<�cx�� ��W-�x���4�<� ���0Pnص�4YU�m��q��th|K�y��H��\U���W;�g�`�@��.j�>#If1cS����|�Z�e��KD�dt�nJ�{�b�g�}�o}0ja� �T(p��zXJx���z0y꾲�:�6m�W������c�Lu�%;��Te%\7p�����s�7����A���I��	l����ˠ7�a��op��Ps��d�S�<�t��T
���#��t�|0�$�ܷ<q��#:���+��g���[8�A[|��[P~�����g���tdB�^��`���b��G�s��sq��� ��|�!\Pdo�Br�9\�E�����������e��*��?UT���Pq �j��[��Z�ME�MM�ɤ��3p���j��x���u��Y��0G�nI$���p�5�h���?nuQڏe��m}��ב,@JQ�8usG-K `|X�~��������h~��Nt�%s�3|�bޥ���
�;���`T���	�l����.�(|F�PЛ���d9S��n�N:eݫ�t����*{�`~-`���1�U�gd����������I�*(�S��ﴆ��wLg�[�n�jH��e�4��m�w�`�M�*�,J�������_�wP�)�.�M�8V+x��+��UM�p��2�Y�!��a�z�]�����L�:��g�7�����Th�y��z�9�(�RS/oQ�끽UcA�p������H�+�s%�%�C�{�\� D���44]��Q�'䕋��#��F������F	�II!b�������D4Gj�2���a,6%U�f�wuI�M�[[�cbm�Y����~��s�qU�I��y"|%�6�̭��\�����w��b��G�*������,a}h�Ca�{v!��yg'b��I��*QM��jx�&t�P��N;p|�"�	g�:���k�ࣇX3�*3/�;�3���@`9�Lu�{�U>G:"7u�k�<�慿�\a�K��_�Q��C��5>���8s����1x0�E�s]g�ő���b��ftC�J���k�4���q��l��2�̰��#_��A�et��6��ed�{�J]_t_�,�/ԌDd� ` 4���"2t����*��8�̑�ny��d4ڧW���U8��3�>�S��X�ݴ�F�'�w��-��Ov��2���vqK$��C��z�B�a.�{�M[t�As.m� �� ��*d��"�ٿ����|���:-�x�a��bAu�d�@s��p�EPr���lB�y�%4ٵa�ϡ�}L(��jBR#�`���1���B(5q"�ҝH�V	��6��QT\1��ｙ7�&�"+C��8���mb��� ��V��끺��P�LD����й�IΰU�ٴ=��j�қ�|�/B���Vٔ5>��L�r�}w��9�Jn�i���a��n-�A�Ԥ�%0 O.�3�$^�Y`����p��������z�q����Q�+�@��@j���(�2~�Ħ��x�$����=������t�'��E��/y��"fe2j�l��2�w�1���! �y���?�3[R�a_�"�ˑ��?�9�۾=����	�H=00)�!�c�Vi{��~t)�B�W$���`��c�ze��5J6 �~lO���i�֦�Kv�H��@�>/^�'
4d�_�P�;?�ͷ ���A���1� Tbѹ��,���Ӥ�+���{1��z�Xf0Y���	����Jԇ��IuL�@�&n972�P�/��>�|C��!%�GXЄ61G����2BǺg[�
�-Xn�M��z>8����l�]~s]>葾�P�_���c�`k��:����}w�����/��͜N��\�K�lPh��7�X5l�~d>��'�gy��\�C/z�y���c��WcW��er�w�W�{,��7n[g�fʨ���U:�,hA�0}A�O�EžO�v��'�0�I�-`�$�d�'� J��V��mU�q�U.�?�:�.I �y���M�$i�m�B/jo'��MY�{K���)t�-�K��=�6�XI��~j4'�U5����/�J����5��0����_'=V�j(�`�6�����ȱ`#�B����A h�ddk0+YV��z2o��Ǭ��$� ΀������[NA'�0���Jh-|2l��Ú�M����z�@E/QC)�e�2�S�nd�Z�mA~�AG��'���U���\I��� ���������!�H8Q�����z��4R�g�����^�SU�/����`oE+)��j���`�Xl�l��b�u�n֏�>�����u�s���1�x+��3Cp�pw�%]���R�e¿^��H;�
�>���i��{V�QUHGG2��7t�%3��7��tSI��ңڄ���ė%�� P����7/} �������I��p�j'd�V8
���}�jv�C>��u6"�����[g�b5]K �*`���(,l)DH�}8'�_':��3�+�@HJE����L��Dѷ� |K�K f%ٳ�j�|�u����z�L��.D�<Ӊ���]q��M���2�-��?]u8�+��5!�rӞ.b�*F(4��>���$L�*�r/R����$�3O{��٭�3��^_���(�T�<Kb�[6�ap�'&?*:}�P�l' '��8?Wf\���(���\b��[lE��)���.�8���B\����68a��o��k���0TC�6g�9N91e� 0�U�f]���'��H8�6yD"���K8/�i��e@j$��5�M:��5R�㧔5	ځ�E�Hx�]�y�R����+�濖b-����1��n��*�a���R���g�rz��N+17B�1˦�>j�pht8���S�p�C�x���U��&�L[޷1�W�L����j��;!���-}@��p���+��u&��>i����/���'L;5l��c1r�~.����~^�s3�*aL�@)�Z՗6����Y��7N�Z��Hr�gQ?�7�2k>y�[�r�J�.��!<U�P��o{O'ww�+�m��#'�`o��'
���Kwk|�`]�p�qz
Ğ�Y�3�Cl n$'�YY�?H�_]Z��3�)<4����YxHx�4�Pl%ZYVN��T�H	�р��ߛ_
�����MB#} ��k���R���q��y�?�h��G݇~���vl���V�&������d%>	�$؜�fZR+�j*w��9�OzT�q���vy, �j��͠�%R/�k-n!�aX�M�G[��O��12j�d�8��~&�qN� �>ywnx������g �(�e�m��*�L�Ut;���N����XJd��;���f���j��	���%t>/I4����)nq���Z��sl�k��(��l� �o{�ȉ�-�=��B�;�%��O�kW��:�Y�W.���ym����Bov�[��c5`��BD�Dx2����N�H�����ݿ�e����2��q�ǧ[ݾ��g*��BW�2@H�o��Z��4A���0�>N9cx���\$�X"���	'o�!���4���T����U��c%�&�,m,+��qE�O2�_RC�h-[kdW��U�&�Ϯ����в��bRW��҄��Y�d4\�SQD#�T�o���@E��%�i ��y��#�x�A�[��@���Q��_
s�����O��B��812�Vԡm+D�׭���a�>�i ����}��תsG���Ou�PB�Lh,j'p}�$�31פ��<�Zprz.��4��-s$�?�Uf�S�7+�����.���jO�����B*z�\���6Z�H�r)�e`rZ50�^]a�'�u<ć��'���F� <�dM�����*eÍ.q�ot�UdI�O�V�]��D�R[9d�t�t�v�Z��d���{��n��V��>��Q��qMqr<�o�9��zo��,�
�Ι�����=��H����bC>��w4�q�H�z���h_s�.ڏQQ@"��h;
�n��i�
�����˂Rw�H������o�v��l�g|NY?dA3a���������F��`��o}��}�@iO�3�e-iM8����l`��S����y=��i�G��k�dJ�X� ������n��4��dV�����:U�q(t���f���?�a���|��R�$>`�Up7�)P�o�#+-�a�o��2�v�H1K��I�6GGi V�Gf��h�<+�(V-P) ll(%�i�G��BҷP��{���Vi5a'�oI̜���]�/�wJ�/���v��h,�8��Dt�@�7�^f���
\cb��|���H<�������� �sy<]-�0Q`�O;%�%w$,�T�JF��0hS&4�%R8���l��>v���h9~9D ����S����� �
��Dq'��$o���1����"&��z$	\V� �)~�P������ ٶ�+5��5[�Y������Ǩ�ފ,�:h�H�9��i�x�J8����i���x#e��{uN�|�gu����P�Kl�����С�Z�[�7�Y�'�V��vZ@b�� ᳽�g�W0�o�`B���F	�l�!*�a�$T^�߮�Xé�h?RH�ǋ���̛�U�I]����k{�6�=���+X~6|	>�C�&DψF�rq#˫����o�1R���O ���S����"����X��x5#y�g9z�0fci�	CH�Un�[r^2�pN��lVEd�M=}5g�I��!V}��xg��ȤU05v\�f3<J�b�F=����'���)[�{������-jyi�'���`W�u�
�q���1fN�EL���uBvF�?;!p��حy�oh�v�^H�)�@�8�ݴ	�����-^Q�p�s��n	�_&}���<]N��jm�g@TO���A�]�[5�{)���g����(��n�����B��Ж�p/vX�vg({�6�3�,8��V sz���q�R��fE��qg�U<��~���Gn#��m<m�5\�Ι5��+�i:�"�`�����4�p��}�D���5��t��*T�L_���2+�A�z�\�oe�_
��nZ�	�fw����f�6QA�u#b�*��1�`���� �wƏ��q՜�HH'�W"0�:ߤ�T����<�:kHUN��5�����~�!r��< �=*�B�$Y{Ԓd!}Ŏ�:�ljɼ�;�U?�ߢ�.�?����K=!��g�y ���O\���/:S��A�\S�����yZ��U��J��X~����)a��v�]6x��1�7��a�:��3<�`^5�Z���Mʷ,�{�k�Z+��W�������ߊ�	�ԙ�x��Xt�.��D��N��s(񎁤����_�Lb>.���l$���� 1���9�D�8:�zd#g�QR}g�q�H=���m���T��M��D!����λ0�&����VԲ?O�xgz|�����-!#eC��~Ц�d�����$��&�n��?�@M�A��~#L���߆���y]��õs�Jo���Ǜ��2'F�H��Y�k@���?���u�H¼�(ATSR|�}-	zb�4I�¡X(h�����ˉ�ۭ���0�G�:������?�r��TM>j�C��c^��᷹�����]Q����[x� a��؃��-���=2%j���O������g-=��N����H�E�?. �y�<�+*��~+�Q��#k�Aq�WxwG��BF_�]���=ml��Pe&�y�6ǕEk� T72kZ4Kj��P�}N����fJ��ڦ�R��wb�r���K]��1��1�u�}D��}C��1��î4v�'v����zF�3�.�^����p��Xr���Y�Pd�Y�*Y���L TJ����QE�EX�B 8��3'��#��j��v�#��L���gz��h|Sd�T� ���"�=?�С`��T�+�U��킲��Oo������nW C]:}V��g�IF�f��sa�^wR�:�)sq%Ѓ)���q��$�ذۥ���.L���_gj<!��/9!a��\�7��;v�{X�_u���+O����*#��G4��9��حS��'���c�֎��.�V��΢�3����2��F�z0�y.��Ct�
���g
&R�@�����p�|��~��&n�Ņ�d�z9/�`�tc�+�:.��R I���|��	�t]k@�^�B!��[=�A����<>�gVۙz4u}vT@.3N������j�'�֭\�2���f �Qb�(�C�w��Q�E��1�hhQ���?����*�������<�5�֡	,�>5�Y�+B��_-�yj�ц�?���^���b��4s8ώ\�)_5$3}�̫�@��4��6��\��3��;�|]��&[��$�ـ~K/'�&�p1�K��*�=��hi��m�Y�(�~G����[���b��U2Ҥ�� MQE7�������Q˼�u]ȼ�3Ri6J����R�VLi5�<c>�	V.��[����٪Ϗ��bnk�=zI��6�
v�.��O��Y���_G;v3"_���?/��.�)��F;�{e���$=��K�I)TUo���|p�H`*aH�� �j��$$R�K�����~������F��̙��h��'*�4��CQoY@1虩���i�h�WaZha�{� ���Ǩ̇�MH�j��Wé�@?���L<U���zx]��F�)�q6���| ���z�]�;�ag�֥=j�r~=�ڳ)P�%�Dc�*� W�5�F���������*b��b7���C�E!���)�O�S��}��Ҥn�7Fa>����t�3P]胣�oc?�>׭A�e��k3�^����R�����Up�-?�7~��
�N1��o��xs���h����09�;)�����e��ÖFzW���k����Aޓ�s8����<�i6��)�M#�S�<�F�+��sy�,}��D�m��d������d�6%�� ���W�.�=�h42��]�6���}�WG&WX�]]c��0.3�b~KB�B|ΑH�>2#���n]w$�b�H�5�܌>��ن���	�I��MT~̓�Y�l2��p�~]U�I��'#j���"��n:���W��	�p�f"�Z=������`�:��jA�0S�!	�&�Y�C�����\i�+_`BU$@U	����)���7�hY�pďE���ȟ6�Q����ռj�	��7U5����DZ�,�?)��λ�\G�j������m��� �`ٯ�*�����H<���q-�#}��G|�w������&�G�L��"���|���yNO����I��� {-O�m<uZ���Lb���NIߠ|�Q��`n�q�,@�AU"�N�H	�xN��w������f08����	p��3�o�7�*׻��"�?�;�ˎo�M�����H[(�m�=�Z��N�x^Ұ��h�����.��m�5��U�f�� S"4x=�D�m�C���]�B�u5���Y�Y-�c}[���s,gI�ƛ�E��v�g|���ʢ �r�B��&O�J��փ�@�v�.!��!�q�̟�6�ʪ����o����'[]��!ڛn%�R�.&�S��x���qa��#,���B��ϙ2.9�j�`D�=���Z�x��jm|�R��L��M��
ķ�+�i��b�X�u��x7#�/��oa:���b~"W5ҿ��z�/)�a�P쯵�����p�*�ad??���?w�b{���}���%�N5��`g0� 4�Ǩ�[9ő�INHm�X�g�Ԙ�f���1��]ש�ūi��h8�|q�z�e]�k�*�����lv���Y]�M�E�����
&�'NM`�ya�g�m�_{��?*/b�^&�)�I|$�/��}0(����e���+��y�>D�}M��S�_G�@��]4�Ǽ���;ȂRS��'�H&e٭���]qϋ�#��$�TR	~�ry�g��<�}� 	�[$�mG���a�������4�[ceK:���x��T{ `��\kV�;ؓN�n�+��:ewf\�L�'��(�wE���9��/nry$;�3h:f��o�Y��.��o����]k��󕌈䐑����XbWm�A��,�[�QVS.���cx���dO�'�Hg��w��kW=~x��9��"y��䜿t���8�piF��!0B�pwq4N��,l̶�lK/�е�S�=i��B���4O*-Mˎr4����,�C-���ߣ�0��]z3�b�,Ŋ��[
8su�粁�����p,|f������]pճ�%òekfH$���"�M��i��uGd���v,.�5<��%L~YR�
�f0��9��v[�]�6��ߟ�uݺ�{�"��[����V]�0E�����w��F=%��ro�n�;���8-Q�
�0:!SW&k�G[4�����2D���Bޏ@g*͑-���B����i@ḙ�����,�5�T��7N�T�
~��fa%Iv�m#�0��ٿ�[ <K�'~5�*�Ɔ-�
���Q�9��HM[p��ȺI��k·:�p�K�[z锹�J��a+3B�2�+����m�}!�c�E�ip<����>�@᷂�Q�\b���R7)e�;珸�I�X��9>5�2�fxmq9b�t,S�`��ۚs(�S�����K�\��,�`"#zvs6k6��1��u�`e��bD�y-��k��ݽ0vJ�֍�T��TrB=i�`?��.� ��F��($�*Uc`4ڛ�%�$QM_�`KM�E}�a1�^��|rM�hw�l�<j�r����=k"&�ӆ����'�~yh�/+���PB��.��E0z�=��)��1�n(�^ё����E��v� ��I�k��F����x�槄��"�a�>L�ǘ2ʥ���hlj�%`�po[h��B>c�R"\(�_�c��#�i�Z�� 1����<� ��Ƣ�3��i3��2��i���r��OLu�1%8��0������*jNӘe�Ś�~/Eȁ6�{�*$נo��h^����'��⢦Fr,ŏw��@S����|	�,�_}A�7�˲w�h`�?�ݓAK^�G�U��S�Qp	�羽��¡��x��nj>`*015�����ރl��1��t�`Z�����]0\3{����a���1ULA�V�\4�&Ʈ�{�B�L���4YNl��ymP/a�ZD�n�{���o�R-�,�?�F�o��<~�.Q���)?�Ҍ|C?������>�.�}IuKδ��B
��5��/���2�>�ij�$�ǻ���T6TLjj�����  �V����۶@uo������25G��7~����R�?�>Z���IRoF(�J� ���S�ML\Gd�?)��|�ǹ������7��i@�������xW�l,6�kaQ4�a!��`+&���(6�D��gU� H��S�*��%T��S�z����2�^|�ꑀk���b��z���������B���@��w�&�������K|a�������(��_O<�d���`Y^ܶ�&}���V�KY����5H��QJ�^�ۭ�IMȝ8���쿺y�j^+�G���Q��*��bN0ltۄ��E�#E�)5�җXp>=b�')_F2�{!����+2�D�(�Y�L;��ᖎ�z1ih����"Þ/��pd�O��~�����A!���ey�J�z]�6�zRH{���f��1�1[�KY���`8M�Kvm�� ��8J�+�b�T����fǹ��v��2���7-Bv��C_/�&x�鱬�2�a�#E}�h����&���u��ݮ��b`�FSP��e���Y��ZKPR�k�Κ�9
��T��r�cbkZߗV�h�G�0'O#7�Z�8�f؈�Y.�?�h�B�ܝ2�t�#H�aOrB���y*-? �^�a�G)e�E�V�P�C�T�L�y{[K50y��vs΢Xkt;���6�N�lˎ�Nî������>�R�?}��1uc:�D�<v=��Yey����;4g�C��οt^u��j:!�a>Ρ�@*Н)�ƊҏsyiV�49�{1�p�;�0��)WA�u|�b����
$�'u�!:]��-xT~�X���%nF��T֎o,����U�wA�G�Sޠ���ٙ�"�v���Ye|g��)�1������y@�������Ss޸r�#*)����>�|q�/�&,�_3�멵O���r񺶧R���`��X���^O�C���}�^O�Ɛ��3=�}�Ej��W7�c��f�
�ߧ��J�ʠ�^�7�Z�tN*D����ˬ�pMM�D�8x�eeT���h���2��\��/o��%���i��"D�����%r�
��`�� ��b�>�uyy0�P�-�`J�c�tW�/k�5G�̤�9�UNUC���W��%c�Dؔ`����*�N�مl�E$n�(�l��عI��٥<�t��0+�-��WZk��Z����l��`T��+ضf)���y��K��q�;��3��]�5�_�����Q&[͂��>�Ut��>@�/��ĭ͗~
����g��n�w�^����9<��F䤢X�nב`���X_����d�����#̉���:R��s��P�,5�-��s����"(@�&?�9���W_,��-���U8��5.��5M�֟��a�"��jQ�9�#��CW���]N�j8�Ʊ>%�
U�,�4�M��P��-�g^�{0I=,B�_ֺE$}��SG+���t#��G�Rx�܄�~�ރqO7�	d����mk��~�5l��+��ن[L�x�Ϸ�P�0� **�E- J!��Uj�gnA� ��.��6�^��@��~U!�\K�����8y��0�vߒQ_��yv�P�ŏ���ǥ�ga2��k�9�Ǝ���.��!.͑��{`#Ov��Va���!Z@��+��y���6�Tٛ�7J�Y@�\�*;��;�䢌v7
�a���6{:�^��Y��;���IE���_����W����λNW7�Ĭ˴�L��K'+�_��;i���*�3��B�P��8��
�����@�z���&�� vZl�x�`N�rj�Gׅ4�:�����tl��e��'���
I�}h��6����O/�u�0�U`Q?�iF�Y�*(�Ʌ��j�GV�L]'�gL�Qή����֊�#2W�x�	�No�܉����8�g�"���z���%mw¨��U�����Q�({�X\������X�a�	 M�=���@I�~�+%Z����06��l��M �L$F�ɀ%�p@�aBS�!1�v�����Z���&�R��KV�QQ�v6��h�&�J���T�d��㐯��C6��oB�7'����F3W�aq��~�O�	)l�	�n-�O>�M�@4N����Q��7Q����"��{@5=t�_k��1�XCq��L*Q�9O-Ѣ�8%^rM"O/zxȝJV�;%Gj�n?�+�I�&fhA�N���Cݬ�V�����n����P���IJ��@iR�I�@:1�ފ��K�S*���P"I>��ݘrO�nN�fGR��!}ЩY�2�i5�D����/�b1�OVn��S�U=U3�g��z�x��m`C���M��Q�1�X6��V5���7�*]f�7����㹙�k�_�D�N�Q0Po���e�=UrȠ�
���I©�w2�j� O �?)f1d��z��b��q�dg%�/�"U��`��űL��4�m'�\/�$� p��E�XU6���y4��C,�N�����b��8�j�X�/G6Bev"-�K�U��|������R��ԛ���v��U@Jk����}`E�����P���1���!Ho�z`.��i��c�-5�x�tzD��
/��&�/Qm��`k�ܞ(BKw��G�<��|�+��FN�A;(���2�	���t��A�6��,N��ԧ�O���	�/�#��3��	l��ń�+:�އ,��=�8�;�@2�j��T�/o{�rQ~ b ����<�d2��ҏ;�bމ:B	>Z*X�7*��|�����W�kġᐛ������!ݕ�[Lk�9'�zb�x 4�������dV����/#�5����_��zNZ�[n�81g]fit/���c�ꕻ/˞b�����o�R�OM|n��M�I<������E��"�վy�	�lvZ�~��Jx�����v�c��2�+��6�/�{��,9�
P�<��CpPDA��D6�M+}7���1�A�8�����5����EC�c��aK�!$ѳݢ 	���(�G�|�@"�<�D�꽢�����qգ�Ƴ�a)���h(U��. n��g��m ��� 
͆PbK)��6�M)�b%�g������7�D�A�)��S���������)�CyIfvf>��X%�ҳ�(����dYz�M�S��?���y�UA��"G{>P+@n��}�^'��(ΖP+O�[���������荽�D����/��M�H�#���3�w���n��n��2���LV���+i寂�(��3mA���Ә<���$>��3�a���x�ү�_�ї}�-}0aB�I!�gK�
�caE���yX:�H�����x�4/�-6������i�yg�=����MDs�e�b$��K��OW2�ژ�X��h����U��)�W4d8ق�7txY��SK��qղ+D� �{Z,}OZ�!Pq=V����������u%iת�m�heLA�F�A3���ώ?���6dM����R__��T�����w�.\140�SP����d���0��Rf��m[T����\�䤝ߡ55U������������w.�o�]�B� �X��U].U�J�~:�����Z`f
1�S�7�B���బ�\C�hn,D6���0?�4;��z����f��ia^���m�6�E��뱄��,	-q	3�æ�����jW��i�)^ͥ�9b�C��_���dpVs�)��ܥ�W��j���!to��=�B4bM�B�p�aG<��u����T-��c��?yל
W�6%jr��g�� ڭp�sO�L���>e��ʖ|v� +�r*��I	#(K���H��j����3��������c`�/��lŸ2,
�WBF����L�"�p{UF��a0#�e<B�:!e1�����5l��MI=��~��Pr:���O���#��7�xw���Ǹ���`��~-k.�j��.4T�QiP�H�u�o'��	K[2���-�
��yw���U�jG���8Gu�5W��;�d�t�k3{*ڍ�9��KO�4���"��U[����IJ����l�(	A�Gj+��MV�咘pa&������$h�*=[D`�`G����0 .S)�i�T����1�]�E�a(��q�=����oz�ɺ\��^Sr�A��r���9�t`�&��k�I�T���E�g�;U\�$��sS��_M	]eM�������*�l��MF<�y-8�j�6��2m4��)|�̔�T�0�'�Е%�ʒ���vӜn��1D닢_[yؾ��)�Xu�gA�Vd��X�����W���I�ɉw �8��?�w����&��|�Eua �%1֤�HRm&_���>��� :���v'G3��F�QOn�_iܱ:b�:�K& `'ٕ)��T�t�G��u���A�?�;��Pk��9�� ��V�?Ⴜ�䬇 J'y�,O����O�)L�!�Y�m�T�j�<�Q��bWo� �˫��et�
Y�^����$z
��b~U�{.�XZ�L��&/���zyzW���|7���S��
�e��G��n���V�y��3��qk{�U+�2D�G������Ob/�EYwS��"<}��!ό����1���\<8��t�}.�(��T4Z*�*�J򎉳f����$9���,!w�H�X8���Q�K1�<��ͼ��Il�zu�]�����^/%朏i�G��
Q���㖵���3w޴���L�;��Ŗ���!��;��"�8�s�ZK�k���r�c��)�W�[V��VO7�u��6���<���:�����/�����бpak�#� X��ۦ���F}��N��"Y	�`��6�]�\��x���N���(�[�)������C����Ŝ�����0��i[�&Y�Q Po��_){�>|�quBȐ��r@dT���J����J��83�/�Ẽ$ޑK��p��v�$�Z�!������iQ����!)bm��me����-C+���y0[jL�����Q:��`%o��`0^�z�Y��u,�F3m;���Ku=��	���^+���l�	�%�S�WþT8n����i��l�jo
���#љ�0`E�{��|��rdAz����@(-sYy������@�8X<Ak1Z,RS}P�NЅݣ��$�Y޼�`�1��r�x*��BD��C2$?bhv��8eu�ְ����.g���hO7M�߸+�
N	����_�	|���v��*P �Ivh�����
1� W"�o�y_�SV��D
��JT�t�����Q�PY��j��.��e+��{�.�7S�>�G�Imtzd�9ũ&����T��J��u�L�\(�gNZ��z '��h�$��%Z��HIYYQ�՘�>�,����M�:��q�����iI����a�/+d���3����b�y�b�|�2$ĸġ����j�S�����݆=���)7��M��5�t�BD�U��x�V��槄��}CA.i��O���L�������q/^�c�+W��SL	�R�Z�N˝ɓ�}��{�����o���0���%>zP�EDd��K�>4��G�<|���������{`���:m���"�iFI��	� v�"@w�Gxa�wEJ�3K��ָ�H����zq����#��Mo*ܓ��̍@Ft�o�఍rDq /3����o���>w���������
����o�q�a���CfȆ�� ������	�
����ki��5��q��������e�h� �&�5��f�9�h)���p�p��}�� ]ꀂ5I���6�L�1�����͂�H����ޙ��`[^˷��%�/eZ���,��!���zbdŗOz��W��1:�m�o�lI�I�9
�y�1�U��u�sfPJV�ރJ3�)�n�⓲�1�:�m,��9⫗��ҷ��*<�Z��u<_n/�wU�-�/#ɱ�R$�
屐�Ƒ��_~sK%{ ����<i��:a�X��Y���9k`�BZ���o���MV%fC'ސ
f���D������s&����gp&���8�F�BcP�4��wp�����R�Ў�]J	ί��A��+|ܡ��G�����5��u�b\���6���W�V@0��!U���R������ǖ/��	j��7|VW��8�ٚh(u�q(l�)2�י
3a���#�y����:J�Q��o�j�o�]W�y���Z�c)'��zj��/�9�1>�f�����W8
�y���m� j�BG�G��9BtZ�C
\�)c[ ��)��Tfx�K�%e�I7�����Ϟ[�
��K�M�Ka�%(��
F��k��iE�e�~��<�vd�����H6�꧜*����^œ�HШ�� �_6q��'���2���\��~�/�h��%$�������/��4�n�y�>���MHv1t�ȌP��vw�xn��P�+PF�r�j��5a#��T3�����h���d�e�Mʎ���-�^��05�`8��f}�@rC%�"�U>�$�&�\
c����v,Ȗ���BG@`]��{�<(tsQ8~%;�"�Q.#1XyIYx1�{ ���D�b<ۿ_mИ�c�d�p^R�D7�T�W<Es.E�alA6�13����5�o��6M�$���o,x�G�C,^Ͳ�G�`I��(��M�b޴���Lj�-���6d�;�_�kkL�Oͦ�b1�<�O����O��Z�x��6�h<���_�;��u353���_��>�Xh�2��������c!�b�����i��8־Ӱ/Fv&
�;ٹߨ�_ŠJ�JZd���1�	��+-��7�s�pu(�!�F�7��|��F��띛�{�	b�Va���0 N*�Y<�D��"��'�����N'��)e�s��|s!:y2^&��Fϩ&cZ׭!�n���KP�sI�z*{Ka�/���V[Hx����'�D��*������	��M��G��#�L�@nŃr�.�<�Y�����&���7��#��#V�f��8����i��a��k4�
�z*m�����C(�Ϸa�!;E3�{灊=s&�45ν�% '�_V�[K�D��ؚ$a�,5�F�%��K��!�|���jwU3�i#I""�G��da	$�Y臓�h��Q����(z|<��Ԉ!J�Q��u�H(���0��%a���)4�Ё���mMʳ~�U��o��G_�������q�!H)5��Y�/@T"]kF�O���
�����D�ާ���*ڨC���uT�����m�4c��j�_c�k�Ea�=���%�?(�tP3�gl2r�`|h;���	����7rT(i�2@j[�k�e���d
'�&h�e�a;�j\V��N�pH�q���H���21��.��2�h��Z��$ϼ�7_m������:�'�[�[��c��L�X�*�1i�6^P�	���R�_���l�l��Ϭ��f6�s�����o�ǛC�I���So�KjCvi-εG�V� ��dU )��NM��ڑ;`��H�3#�.=��.�e���NX��p)C��;��79����P�g�~qסrz�s|��a����*d�8Aj����a��f��@\b���B�~ぉҨ��_ʹ�6��e!,zQ�YO�ܥ���JaQ���-���R�����h�з�����~E2�m� �̓�8M
�ND��,����n�B�Sn�M��1��cYޞ�v�?�r4�97�^�"��	����si��S�@���-ì�$�����m�.rR?m���b,��=�8��������
�(�[5c�Jbׄ��R�8to�gkN�F�/�_�KfٙC��,����M���&>"<��-"�2+���}�,�O'����k]k�f�-���qer����@�%b��j�xۈ�z��i����6O#k-I���	�rD���Q��Ho$R�<f�H������}���"3
�F�@�*4
�;u�b3����v���bg�[��/́'Y~J@@׷$"-�)�n�8=��0-��N@bY����y����J��^�n�|s�Pn�H�3 }�<�q�v�L�3�@����G��^Niփ�;mV	�2�rdu��ꈁ��h�] �8 }w������^�5I�ꓞ{|�3����s�bmƐ�P~h斵�S؇�K�=2�C��&v>:oM(�{� ���_�&�s�9<���M&��QE�ϩ�",#��j��`�9�-&�8�C+_`eW�
rH��[�&�Y����?��� 0���瑮�ى���V��b4��\��c�✢D��DQ�� 9�FHڍ�e�}H��Ӌ��lŵֲ�$�l[T�x���U`V��_{^q����W��N\Y�YP8��E޷�h/j����6�o/"���^�UB	�b>��#ha�05��[p�mV�Ⱥ����i~r��lI״�J\�䘩oa�I��'QX���'0UL�TJ���@a)��ك����b���V(f~+ەx47ϑ7��
��7*rl#�*c��.�����eVG�-g���yhk������.B�#T7�ې͂U��dZu ��/�(�԰:�'�C���(���z�x����[l,������U)<:�60��q-ːc�ݿ9��k͓8B[�������O8���8��%u?Yy��G�c#_����֚��c�t��s��K�Rg#k�-)�O�*�C����ȹ�1���6������5�}z�Y�� �>ϰ��R )eKj���K\��<�v"��7�KJqI���g���v,Ϸ�����/G{��Q���F�B�����碉�	$ �pϯEx��n=��P���>��b#տ�ĥų��,��0ڑx/���㱙�u3ɐ�3�XXs|U@'th�?�~�}U3`��.>��_m*��`I���*�Ҧn��<H����N�93���d�]}���t�R��<;0D�k�����ѐ��$��b��6R�f��"'(Q�gN�����C�P��R�[�M�䱸\V#Ki�H��!fT�i�u,�r�6����0��
O���2�ϻ~V������F���1\{v��nh�Dе��$_�ZI<Aq3g�;���J�Å������:�!�� ò$R�Y��c՚���(��8�LCn0����Ql����l�ů��V��dؖ�?�����Y+l�Z�~�E��m��y����2���Z�:�˟0�l�ޏ���$=~����@�j�fJ��Ds�8�EYc��	�9te���v�f����0�b�2�>��9�MC��rb,׾K/ZJ�%_�}l	�\����!ZJV���߾�ߦ��4}�
r$b��֛bi�o�5�G$��%J�k7C���Dўʧ����-�ES�>~Gw�n�ڸ�����������Zґ�<W�d����ѱ�x{�l4=��W����9�,�����X��*ex��mP�=e�m[Ai�L�I?{ˍ��t��n0q.�>�Q�r�]a�&��s^�)���i33"Q�O�s�����a�`1���,|E�uC�l��~v`�+q`�ru�h����v����bHJ�uA� �Rk���L���ģ&Q�n�<��x��׃�oj���)�����6����5m�#Ϣ{x�."F�Rׂl�S�a��(���&��t�O�]n,�s[Z|Xp�b�`�O-CH��x���hS 3 ����e���D�5��/�:l���Q p�~�,Zu�d-W��|G@�1B���S��I:�$H��$C��V�(��ȅ�$�q�q�#�}`�r�6��B���w���@��I�V���FB�m�ʺW�}r"4�1�[��(��O"���
��W���j�f$Tya�4��JlK�TN�o4��Fr����:�����s�L�4w����I!;yϘ)a�X$����Ih�?�v���a|�vp?#σeN/��6]_ů�{���9WZڤ����U>�����;g���-&�%0M��I'4����48�`=7O��	��΢׼1"q,u4X!-c6~x��P�z[�a��ig_�A��Ƴ�,5-�h��!Ԯ�^Z�#�;"��W��'N�k4��x:��u�j�������5�VP4���O��㤮@�P�#!�_�Lr4|/ڬ��W<����b���U���������U)h��M�ى\�> &>R�����O�Y���>ק�/��lT� �y�`)e��7�c{�Jě�mp�3u
�B��{��`�3�J!��ȳ��C����&P�֪O�"2�RI�a;�N*+�<�F]Z���r���|`D<�.'��k��\�:Ro�$���t�i�(7�T�5�å|� &�\��o���a�zv�7=�Yg_*���k��I�c�����)�7w�p1t�bL��!��^�}ч8�l��Ր���&�`�tG��Ю�k��BV��q����A�Tp�cx0��`A	����(pHȏ%��b���o9��%��<�c+|�b�8ް��R��E���o9�p^�j�ٱ#��Ut�,��,���r�a<f�����S����]�O�]m����ֈ�!����2�^%|i�QF`�<r���{�f/�$u��z����/��H�,Z@}H��{n�5��U�h�7��������tY�����L���d�2�,F^K|��BujM��&g���y0���O٩>�=�_Bn;�;�` XA+���DP&۪�?>�����H�E�I"�(O��0�@���iN�(p\��A3�Qv/��
a�S��~���$�Y��Gh�E[
�	�n���_2;%�3�f1����y�b	wb\3�o/�!E^\����Q̴e�R��{NQ�x�������"��nAcR5�#���&����u/r�eI:�>���� ��E=?����L�/��c�?SI�U �c���9�1���&�7��:�( �b'�$�oz�Qa��k� j����C��*[��G��q{���A�0S����c�R�;&E�rv�<�\\J���/S����<rx�(�HEM+&\��0�d��_�O����Q��G�7�B�"��*i�x�̢�-��>����g��%fg���"�H�z��A�5�m�Ľ5+�"<��J�66c7��8׫,?B\5��J��!���?��D5��:'�!���]�Z/�N�Fh�U�4#��H>�8&*�˱��g��'���A�pP��}�����Z�����HU�1S��F��	����_����϶���s��$�N.	�o��:C
m��9xj���|>|��������L�U�q|�2(�]�����k/Iﵝ�&- I8^P��^�l���s�H!Z�{<�rs�L-w�o5JE�����!��-�a�39�4� aP㆖扠�n �f�]�]x� ���y�L!�}x����r>X���;�Ҵ'<Ql@!q�Ō��fG�t<��?x-W��a�5��W���'�M�ƽ-l2�Rw��J����-�����-2]i�\�� ��g�cm�v p�����p��у��z!�����z6Љ2w=w���/^d.�g��|�r�j�@�i�]�.����z���� ���F��cd�,��k�fr��A)�x��.�Hӣ��%Uc�x�g��QN�MK4��!]�-l�i��!(!b��3�Z.4������o�}~�xѬ#>�Q�>H��C�
]�۹�Ɣ ��|W�C"N�Rb5�� LAW,�oB��T��$�-�L�W3~�05uMJWΙ9W����Z�(3��%�����4��TVT
]���	�)�ꚄK���f�u�R��N��p(�.^vcL�8�{�(�JD�yQHh^�C�����At3j��Ll6���|Ŭ#�ْ�![��I6zk�6�n3G0�'�rE�K�V�ݢ���A1ت�p�Il�wA��<������%�]�eSz�sċ�������}�a����S� �J·1z���yy�u�&m�C�����E��%SKK�/v���~B%�aɛ�3��G�>	�M�N�ۆ�`���Ą��n�ȉ}�q�<2��\Y'�?�%U�hF^�S�`�=WQ9��XR�ߣ�B�o@J�"<���瑣��=Z~�:&b�.��W�u�_�z��IY��Q�X-�\c�z%������Z�Z��z�����5mà��eol�9�ªo�q׿����B���8���Ƌ����R��f ���}�A�QT*]�Yۂ.������|��j�Pz&h/�A�J�ZXWgi��^�eް�6G��l�唚ۙ3H�y��%CY��"D�͋��>)�_s�UF@�mH�;'�p>O_�l����NF�������;{����č��&g
��S��w���� W�*��ҷ���Iqq�Я�r�o����Q�]DT�G귑�K�P�F&@�1b����W��~�2��$�
�U��?e�4��HS<���%�B\F�M{��s�>*>��=m���U\��L8(T��>�`Y�/=��Gt�sN��V�v��[�]�P1���n�{ғf����|�ѥ	��-�?�5#��7�S�{?x� �w9��zJ��-��B�*�QG��)�疩Y���Z��Vm��;�vYȏXG���7���R��L?g[�zv���}�e����h�+�����*�_�U��S�T�� ggD�i��xx�r�ŕsEnW���J��$U�5����Tx����[��>Tk���wۜ���]�UC�!�90�^�� ���?� Kq��;�e��+Q_E����&���d���� �G���P� ��d7:�VY���X�E<�z�H�1�&@o~�|��f[R���B�@���H
i}��h!��_G������ɖ[�S"����`[z��-�@�O�M�4�rn�TU��V7��v���G(2�%� s��7mg#���?�y�'�5:F��w�~P��I���er��Ł�t!��q]�K��b˕�i���Lj'�`oc���L)��,����e�2F���8N��FbY�TMޔM�;��꿻���Ntz�i�6\6"r7=�V�Ҏ��$�́큮'3v�ɳ��f���.sX!��_\yp�V[R��Y��f��#�n�Z^��,�c�Ͳԉ��N�������?
JIMݠ<�xn���xa]JO,��Ҷ���]����H�!v5/&D���=��=qm�Ĝ��ޢ"�_�YN'��cr@B�h%�n+TL��� u�U�}&O~YD֩h�5)�ŕ�b�ػ� ��q�-��֨������8@x)Y��Ē ]��&�
�+Ĕ�<�0��\=�>�`b<4G��9H��f#	���@���95��!I���V�,�y��@q��踳��^*RG�D���j�[U?���2T,*b�L2��Y3�_`Ms�!�)X	�[���i��RtA�D�@ax]�Bmj�D�������Pf���ٽ���N�:�e0�M�%W�ֽ'"Y�����qh0����0����e�P��C�@_���#�0�)%��z��mԚ��v��OCAC���	V��:k�蕀
8;��4F 4Ka�ra'���;o���3TO��pj"�8�]���A���%��u'ݜT�ϧ��]~F�[9+�p�`�8���?"�{�A����V}�4����*���āp�l�М����I���r�ˁR��s4�NBa�����z�����W����t���O�+a �9&$}t��?,�QE����H6�T9�y��>�*u`^���=��?������e�t�.��$2�!�KK7`�6|Qهm��g�(�_{ϸ`����)��uc��3-��6&��k	�{sH��|�<��8�y���������bvٚ߂��F5��RA�NT����xq^du)Zv����@�E�f[ bx�~"���<�Ŭ,395Q��V�f�L��q�<�y��@�Ӌ2.X�AC�jaE�H���R(���Ez�0��RG\JH�����+��Y�u��-�[��,O�,s��Mw��!���7
8UMd��M!�&�s�m�ܶ�i�O����/�5r�O�M�D/�~����{�#���b���N�/u�I"!�Zv.���ݎ�&U��#�`a�*�L�,��٤d�7�[�=c�͑��js�{�L�mr��a%q��T���'��3�mk�;K�? �Y\��Sc@Y=��|���11�8�<TWߢ���5𠠢�,zC?�A�;@?F=�C�Ĭ���ÃB�-X�8j�'8�-�GV�G�Z��T��	jY������������>mP��!\\�x�;0������yO�`2��;l�^��a�+���#���w��_+^Ѥ��*�\+�1�X%.���G�,:n�;����˪~�����R��6�y9a/����t醊�YZR|�$�����(&�9�=Ã��1���QL�ϋw���D����d�(���U�O@�r#��g/�dϾO���cI�qB��hY2��Bah�������=��;�I���^��Kh��<"Z���a8h��v1-��Y��9i�z�tgDː���B�a{瀙�R�S-a�z��%4��ѓ��'��0f��Yw1c�����&�2�c#
���P�}IO{Ʊ��A�R���\���[U�ߒ�)f:0ҳ��2��'K�!nǭ#� N�J�f�X.�O�*aR�>�<A�D��TZ�^uP�?r5kEJ}%�~��1ې�]V{~&l���u�D��SD���7���m�P� �PfL��Pռ^�DLL�\z�Xu���Q^��Q��:������r)m��3�.�����E���&C���ͶP�l�7snU��"_`(��y��i����!�k�WҤ�9�RZ�˵V K��e!�I��o���S�̵f�"#)���\x�6f7$fy�g����*j���Z�����e��L�Z�|��?�K��``�y�M��{gd��iɟ�1��
��#b���sNYج�O���Ej��Tz�0{ꄥ��!�Y|�!�q�w�u��{���EX�ԗ��|r}�\	�~7�����$�dcjm�A"���ݭ����E'P�� !��P_N�O���{g<G�P9#ؾ��-�:�����\dT!�zOF�OF����;�	c¦4��<,�p�G�F���y�1��'�D����Q����K��Cѝ�6�p�.�����ǎ�bn_�I ��X�k��f�}��a�]�R3�	�H;�'K�V)����+�:�ɑ왚��3�'�a�G2\��j�mlQ�~���7�U	$��c[��	�ٳ_�J� m��_���S3��U�������X/-'�\{hlHJDš~ף(�(A��-���SS��δ�fkxz���0`"?���{���>�wp��p�hmlǫ:&���a��/��
n��;)Zr�Oԝj_,��8�R4�`EI�_hl��W�*Ԕ�y��բw�R��L�4; ��A�ՐMڢFUΞ(|�<�>�i�j+�2���A��N�IniT��d�`�8���q��Lr$�ʖ�~o��WG:�E-�,�ڲ����0�Ο��˚j��f5��aD-�Z4��S�0[��}'5v$�ߴ�ۖ@�M�\��D�s"���
���|��ywt��3ۧ;��ő������#���aD:{��b�<�^pʔ�$Q(k��޵'���F] `��D�Õ]��Z*�ħI�0�HO?�uY/(<:�oG��u�ߐ�sġ���%K&���f�*]Rv�նW^��f�Ո��1#�#���M��(��x��f$�D՘H[�!�G/���k�K�O,A�M<���J�lL/�i�]�|j�x�I�n�%Qg�F�wh�p�/l������s��a��ɛ�="0�!�#���]!Z�B�����:�}[:��
�[?㳤��JZ�.*r�|�y=JH,������N����KR�o��.�a)u8�hdKo���8Z��~�)����^�m�J�߲9r�+�A�0��MK�4-ە[O�HCzdkՉ�|�s���������[o�`���9ֻ3y��d��+���f�+��׃/��D�P������'D3.�f�G~�����N��е��Uޫ��)�/IL[���)��'�GrF��4[�,���-�ʝ`��p�G�W�UB��*���ga5��U��v��5�2��c����X��8�+A��3M�wҸ��t9�W�}"{��,d��Y-훢n0�%�"C��cd~00b�f�}g��u�vq�Q�CZ�����?-E�[R��W�+�fr�-D0�3}M֏�$�(�>���Ay��j����%J	�M�膂���ܭ��������>��u9c\<Q�u^��-����3-$��Q_�)_y��Rހ�&�/ᄀ��n�`	1���Xr�y���@%�5�n����ߐ�n������l��L�K�в�@"��}�ڐH�NK��[�AJ�����6K
�?�2P3��X�t���5C�uq��Ԍ|����pF46�A�R�O�Mq�^�x�;~ V����w�AfЩ>�B����#����b��/���(�:T�V^�+���ĕ�N+�,��n�*Fx��)���{���.��C��Zm� ��r�s@�D���i�0�"6V9v9�Z��h�nY\��ȑ����U������Auxg�]-w�iǔ���1I	�=��B(>�\�����1����ډ&11i��# �[��������Mh���,FR�U���:��Dc�&��D�&�Y���ĩXJ�J�rtYb5t�υ蛻 ��C�e�X�h#� �"�{H�����]y�$�f��[�ɻ�ĤlU���(�/g��?(8$�5��+��~�(��3���/�U�Bs���Z"�����?�nY���'�o�LF�\T���`J5���lWM �*:}c	J�+��C�s�"�p�dP[Ƥ�3��WbM�oV�GvB.*%&96A5��t[��a%h�C>#ȇ�[o��Ø([��1;E�p�����vQ�/�x�_#�LYݶ�+�!��?fJL����\�|R�mR5H8,n)�l�uc�Xd���'OjW^��cc1��1�-P�'[{*3��{�����~`VpD͆�I0���T�~�������c��H5�gbYt�3�%H��oX�4�󯸅��CZꬑ���@�[�=e����-�-�P[���6��4�t����j�x	���	'�zs�	,���_�GƎ��&�S<�&�o� 
?*�ـ��F���Wv3n��O�I!j�b=��d[\���=���4�K��H��/ԔjC�+�U��z�⬈�tH8�qa�#p�
նpapv�� J`��g:dA��(#EY�H�ǂB��=M��4:��Qޅ�L,'�ֻd��X�V/nk��X�;q�W�Q1��>�Ү��F�a1��oC�>��a30$������1��a��&I���1�"V�7�7���>�QJ06�!@���vv�!��R����5��?�o:Ď.��a�s�'��+76�E��*�n�yؚ��E�P�f�DS�̦ �Y$qc�h�S�����r�fofqa $�n�{���ɝ���Z�)�*�6����x&������^q�@���^OKr�QxiD�*�#�XJ6 �d#�]ik&�g^�0�P�`���x����մ�\�aEEk���Z!���)oty�d@�9���~�q춑tf�D�J+��;�H���mGY,�%6Β ����������G�#��Bo��8؊I!4�d��룋Fy���:��Ku���V4��M����w{!
J� z=KP�b-a�J�%�i_ ��c8��ۤ�>�� �~�,�b)��N�*g���va���aGIB�<f������d���:vZ�ٝ�B�.O�1��g&��93ڎ��֬��U�?2pO�?ˌUH���i���:��!�����P4$(�p�x�Y�P�:K���a���#� ��n2��Mg�xw���(��c�x�<24�2o�o����b�G2y����-���%j-5ƴh;�Da�	|?]�T�}��s�d�m�r\>H�O��e��n�݋7�i/
F�h��m�Uh 2K�y0KÇ�ƪ�x�gxF�ß۶��M[ ۘ�DΣC�;���9�|pq�^1�2���6�LKI�����y¬Ia7.��V�_�!��Y����&���氀re,(��<�'�IE��07U�C?q�f$�G�uǬ4�gDD�1e���GL��╒�:|��(�X���_ȁ�,�
(�Mv�c��yY�	���ʹӵuH�u?��/{hX�I%�/����(�$H��b!��&�O$��j����Qr��Rw[�q�A5푍
TV6�_ƙa�n5)�h-�ˤ�*c�H�_W���T(���<"G��YsyM�v=��G�U|u��yX�vC^RA�?�	�T���eP^�Eο!�,���^�M��}�h��~LfӃpq/���9�=Q�1�],�,Ԇ_�o��T�> �u�4���̠9��&Ӹ�ˈ��c�9�6.]p�K�0�"?�oq=�bĈFd���+�^�'��j�r!��D�Kĳ����Z`���a�S�R�"U������@�?b��g��E��hS3h�<��Bba{�&Cj�>дWu��0����Zw��{�<�M�YD+�{�Q��1��r5�i�O�%��wAd��Rŀ9_IiK[s|����5��M�ѶzӓmF��ɮ,"M^��i�{
��@v��R��lL�{�hu���S���ۇ�1��^}�r�;⣭ޖ���f&�`wN�~��Ib�9˒!x�"�, 48��?�M�TL�$�����=}��|��AM��
�;�����P(m�zb���)��м%�Lߙ|��n�x��xA`I/Уs�c<�0q�S��m��&~*�`u7�̀����e�|��E����cqs�P��|�veJ�~?É�rxzj����+W1�ptm���1�\q���{$V�< �����dS�TA�8���If ���5j�����'�;�LBa�d]��
2�X��B*���V��WC>����9'B�����kR�����h����ş����p���x�\t h��q(px
��<���Da�b��|�z�B�����Q���^����OHY�m�h���F��3Է�z;��?�VX�7�=8͒���宵��nxG��7!�6kҗ������Ʋ�6�Q=0ko מ�Y:�%J��^&NC���^� �t��G�x��W`$�q���������!r{�]�ڭf�H��B~�K��w�3t�&uhu~'��$����A��wo{3k���Nz������r���������ԗCzN�y�U���p�EB_<K侯P���|LP�Y�iv6�<mp��0�d����~���|�떶[�՚�gU�*w+u�RY�\�������N�y�rr������������	�*�-}P��v�* �6"io��r�P����o���+A'}雀�ߟ6}��5���Oi÷��uѸ�V��LW}P}�y��׫��{��}��JG��`Y�l:�7�S���$���Ď+.�L�?��P�ȑT����ľ&�>�G���2	P� �2>3� 8A��͠.j�.	���l����j@�� T�s�F�F^ L�y�.��';�9re�� �R�^lɧ����{����:�؆k�̖����A��X�;Q�I�����^�\^��ǿ�'TA*�8�ٺ�y�cS%UxR���V�0��&7UQ]�fE>�4R��/�V.ri�?��m��� �1$F-[v$ ���Aam<O(�~�܂h��~<@�����F��F�F�j΢/G5��@����/�k�D���㉈Y�C ,vho�9�50��?��y�P$����ֈ~5���;$홽���=��ߑ�Þ�Z8W*}��WPU�?�e���P2���w�X8\C)�/4Q�1�Ƨ��bK�wW�-Ƞ�<a_rm:��B*�~��H�'Z)d*�#���0P��T�~�R�dd�r"Y�hE�`Lkd;��(�U�h�R��g��w�^��v�p�]�����vm�Yٹ�^�;���xUpX�7KW���M�N�>�-.�<��kWq�� vX��� ���8G������'��i
��+�x;:���1��#8
�ez�����`��3Kr�-M68�=���FMVw�Պ��Ge&�v�Ϣ�ʆz�Vo�8�4w��HTj|�*K��ŭ������M�Jx��1$��5�g�2C�xc��OZ���|�Q�9FrMzF(�Z|�"��g�(��gjw����8�ђ���c�v� �Vɤ����\a���aV���u�4�@[^�2� m�Je캤�Y�\a]��w>q&����,(���ڿ��3,���e�jV��#��VB�L���`�au�����c�Lחy�5���TlU'xc�>��F�rΘ��1�,�@��{	� +EtV��m��}E.}~�<o���u���g����c�}mp�(��+��#l8� �Ѫ��)��Hz8r.��yhdz��VXt�Pp^$ N2�]�UDT�o<�K�6+�j��[9ޒ���p�����L�k��L�#����[ꑦ�����$��)V�;΢��e��������vײ�zvK5�/�����-t \��GP~�?M��S=�Vڄi��ٻ�9�+��/z�\~�p2�u��)�F�&�#��Nz��L|J�sRپ�?}y�%�"�����$�?��O�
o��FA���ۈK��Υ~2��:TSnS��>�Sp> <��1~$sR�/	+[�@��(t΢�v�+�ה$�jk�x�[��m�N]��~�DL�����ITɩU�#&�`G�w9��8����(�MR�Ң�`<F���vM�Ѓ��j�?ѫj�VN�9�:5��~$a
�7�C��)b˪Ǝ�D��O��� '�)U������.a��#�x�O�pOV�$���Wж��Jp����>�� �3r�:�Mޛ��E���&����(B%V_M@�3� `+Ϸ���~�>��N��)��n<A.�#H��L�>�H��Г�"cK����%@��0�b?j�6�Fa�<u��X=5��Wh¬�<s��.��%�Ȑ���%�U��Y,��g�	���Ȩ�D_�������@9q�M����C�8p�S6=ϧ!(�f������#���o��-�`����Iiӯ�e�;�f(���n�����W܄�F��r\���Oy���"Wf��������]���:�D>\5h�9-������g�l,Y��|� c��la%�p����o1j��`����i�J�q��������JUG�ȸvF)U߷[�	�������:�u�e5\^���d��*�h�3,��T�����x�*���|��˟+������Pe��Ƌ���wݠ:��M��H׻�h��Lm�t��5}~�[`B<:�y���Ļ������\'A@t�a�_U޵�L�'B'�(_/�V�V�/\�(6L�$��>Ɖޠk���,����~�t�r���E�45u�*(tZw��l�� E<x#��!���a����a���F�m����Ӄ���X}*�	�/p�Q+�����D~���0�����Кȫ�a���N���*����S亥�H{��h�?����ܖV�`(�_�<d��Dh��wvSTd��*�$�[�LU(HpTMF�'٥b��|u�qգ���Xĵ3\yc_��'��pk��E+LPA�����d`x�7m��{�^��s'q3~�ϻ�Ǻ��$C�,*sذ�o�7+�讠�M�|�)b�0��#�ڬh��؀���&�ɀ��f���rIAy:v�2�y#�^�dD��lI�)Jv_�z#�v�j=S�|���S��NS&b�_�U�>-���4^�?0��(L��I>H�a�C�u�"�b}��H����4�u,C
B�Y�A���!6n#{Ô]�́�����h'�/z��=l��l�A�*��6 �M�Lp3m���.���n��L/�>;��=rO\�8  YÑ�[�
��w+�Ϛ~�B�?�� c>ު��Ps[:��r�xS��O�ptd���X�0L�"c��~��o=��M���{ۘ�]��bq���J@4#bQ��w�W0B� �C����w��BH�cΗ~��A�R������B�H�����ֿ���<&L�O$�� b$*nE@�9�W�P�6����QX98�|�l������}�k��h�K�����,V���A���<+�7^�O� 9�@��j�;�i�G�T��!WU�&�(teɁ%s��oG[Y��"�s�����F���8��\
A�[P��Y6�u>�m�R�N.���`�5��tU��|N��L=�k6����4v�P�e�wռ����|��è�͖N��q!u��4�"rQ�!�ȼ:���C��-Q�.s���� bY���U��!����)iGQ�&](t��Ȩ��� 7���PM�0پEyݳ߯{5+Ú8�w�xa��`�U�M�u�b/m�s����p�<�]st�1v�-��	5��5�8Ӣڈ�uA톋&j�h,�пQQvq�u�"@�>����5^�8*���z��Ꮆ 4�P;1 ���
"��y��G���}�ۦ�����ܺ>������� �"� ������������V���>�v��ַ(�9Bo��M�P!`���(1h�R�n#����47��
���l5�d���m�*�p�7	E���F�L/��M(S/�K5B�W��Wl/�1��f��ʣ��� &�胨u"�������-H�4�8F���U+2�r�-7�WDq 
�'�9�[#�6����t���;�~��g�z� C���S?I=R�R`e���IA>�������=$�6YZ��#B��
��edoOY�X��H�\�̝�d�ПJU=�bPF���܃MX��G��i�kHYX�>cY�ޟH�(���_�㸴_�C�ùm��;:g�WN:���Z�f�$�틴�b�+*~a���US���k����q�s��\�{<�Q+9��T��k/�J�C �-خ�Lަ�����9�<��_EA7GЕ��4a�n�7�;Y��O�� � ��'F��Y&=ǒ�'�l�X#�����1O��u��p��7kf�椡Y��d�������z6���}�1�qC�rގ䟑��X'��f�xA"���5�xmJc��[l-׃�|T2�8{�u06�'�F�g(9Ʒj��������_�߻n{'�}�#XJ��'��f%\�.7�H��D"��>�&L�Lyڹ�3��!wr�y#�h��]��'�Nw}>dr���\� ��rռT�K/����Q����O#CŠ=6#�{�����M���1�8E9:��L#�2�$�#!�����8�C����c�p�3@p�H?��XA�n�m��c�>�8�0��X��C�V���V�2m^֦�\�K�lM�|�4>� Xq��f*��c]�)�Ù�'#�0����|4AL�Ƕ3:��	֋._"�.6I��	�A�W!r�7�k;ם�R�,�;Y�
h�G�k*ּ@R����kw�Y�V�����c#��������C3A8(��7]�4��vWr�-Tml}B<����5o��6<]������Z�t����t��$4�?�d4�C2��@����ǭ렍.�M�\�#a晄�se@g��Q��{�����[����*�Ɲ���4ҵ����;����{��m;\>�6
�q�j���7|������$��Ew�����\�di��L���|�$�
��@ԭ�/��Oi/[��u����C�n�m��g��֡���]^�"$����l�n�ŃEaZ� ���Sv�����ӛ��~t'=.��!��6v��Ë�jT�B��	;Ԗ���.�ȳ!�;I/wF$��(����7�5p�^�Wa(�|�P-J�@���:z�+��ߌ�L���dʺL�\���\
D=�ܜ�'�ҚG���'UU�B\�P?zB�'DK:���ex7xA���(��s���Y��B-={��M\.@p뭻���\¬�C��ϔC3J�䊦�a_Y��&^M�T�y�z�3�#��!,�Z�Gߙ�Ī��Bڡ �9V�ă�ҳ�I;ƬDOQ닖��n� U�l��
_�!T����^�Tp˿~�͌��_��/� @�8�}~�x}���6�3G�?.����C=a�mJ{��Ρ���o��	
79P ؗ���4��J$���;��p	�O���Z�/�(@e��wY&������븾�^�����]Z{�0�γ���Z���6N���۵ 8�-o�+	8��	�1�k�f0���*.^��+�6I�ݰ�6�*!��� �]�+�v%=�gO�5�=o(~O���U�(�Nߣy�I� b�sR�ZO�bjq�� �uq���D)��D��,���)��|s+�0q�xt�%h�y���,Z�{���1ܪ# Q<��s~���2�)9
��#��N�S!���^��L1v�K��<@���%�e�=P@�&��ȭԤ��6Xқ�ҩ�L'ڕuq��	_�,�,Wua
�i���Q6��*�0}g�j�v���}2]͓8sFL�*۩S���md` ��&�i��coV�i��Q�y2��8L�:�k�Kn�ɺ��i��5��qw�2�!�nzt�J��Da��L��|�C�-_�T��tRY�C�!t$2�ӈ�\��:����y�z��g:p���i�������0p���6=�����#�Y
 S�����1TA�d�_k.i�\]CY�R�|��A�Կ���
|��t��Ncp�]���bרlE�i���������3�[Б|�<�;��ҕw����cJ�z��U�x����?-���^5%w¢�鎪sm���v98O�Y�����_ �{<��T���
�x���E
�S����\C,Z
|m�%��d6چk�P���W��I��bA߇~v����W���j��Mv�)�_"N��:ઊ���ce�L�����ʋ�Vn�KMnEOO�-���djOx�k)>�X{sW�!|��\���^5p��V��>�0�^�sX?���t�5��ra9�?Gy�m�)W�����]叄f�]�qnS�q��.�U��Y"�e��*��5�1:�gW;�;�iNA籺���Ƣ�$�O�(��-_���
9p�PQ��G��-�L-&�M��E��#���Q�bV��-���M���S�W������{H�J̒~�e��.��V��`�?u��J�6�
��©�\;� f�+��s�h?2Z�M$E�g�9��/�)I�q�䊀}z�䃏3�<�j6c���@�� �$���k!V��n��殑��`��E��}8`1�5~,��� /x�W�繐��N9Þ���f���2/f��5���cM�?�ĢQ:2tf�GO�{X�6C�s\�s��岗ۢ�yl&7��0~�@�k�V������َ-/{x��JQ����%����|��,@���G3 *h�~��/�w���� .C�}��/���Gᦹ��}�����@�����4߁d�S�*M�ȫ�i�,Īw�by�Vl��Ѳq�0�q�V�NEao�u�%s�t�G��oT�^U���O�.=�R��%H�'��1�g�{ۉ$���[�t�۶�����;���Dn�F����ȏ��mZ�8WT��XlJ୺��b�5�^j������N�z�{�����Т�9��(G1[P �z?��nwD���S����:$�6�rC~R�Ad]��C��ݜYH���WX�[Y���BQ�1���N����>���ć1P7��N�d&�=��H���*���ak�Z:��x0矧d��X>����3V�1�e�(n���K��aT��9z�Gp�
Er��
��;���k�6*I���p�������f�PQ�$�d�B�r��c��.���s��-=w�'�߼�iV��L��A2�m(�Ү4+�J��6i7���2���t�����YȬ(��d(�[�1�RU+M�!U�5nҘϦ�q�H,��ʑ[ja��r��̂%M�&H��Q�$D���k�	rD}��D�
c.˸T�U-�ýa��y'7^.:�%� /�v�SL) ������������&QJ���w*6�Dt�uuw)�Xdc>�Dd��xT�4C=��pw��w,8�L����x��'>��U>�_/�_k،��c��fP�-F@��[#�%��zUOo�� lhpX�{�?�2]�*'�rf|Lr(n�ӚM�Fxb��7�����l�nT�)6k����wQd�pS�`Pl�&|��/���vѸ
��M���).װ<:k�j#��y��Z���m�����y)�/'۠�Ո
 �"}B0����!������;�SS[o�:����/�BBu0�R�bfu{w_�}�̦m6C��*B�P��G��w�n_���	ja��T����*�8W�� r�"�#C|�Xa^�*�e��/������X����q�V%vUg�E����nO-L�@�ߡqYn���T����?�>_9`Un�,ń%��ц���D�� �5&�f:�K��X��%@���ˋ�u�_F͌��/���hx*�QZx�R:������3�@�mwϰ��D?��$��I�ˉmí�S���;q��}(�}�.Qm�|���鿦�p�#}b֓0����hSX-sY�y��xH�mT�	��^�����^5� ��d�n�n�:��䌀�#��q�O*u�r��Fd�\M}Sj�j���X1�d3RoH6Y'=[&tԢ����I.	<k�����;+���t�f���$�g��C�{��̰�+>EŮ��Ӣ�-�59kX�,��a*"�;��<:�����9r�n��¦iy��X�Lv�4��oZ�����]c�3�*����~B���d;�ަxl���Km���P��������n����|Zs#J?�����~2J\׊�dؔ/��NY����,��?1g�&yq��S�0�`j}OĐ�.��s�����M��!(�vfg���8�9 E:��O�T!&{lk�P�ĐI��q4Z2�8�ًJ�cY��m��s��r"{H��{޳��ٵk�!�"n���g�E}�!� �`��$,�y�"�#�������G�O,��{�TwQ�#-u�������T ��vEV?�-N�;�JfLgI�ns��~�g���>����YiHB��a���Q�5�wB�*���[d)���D�c�N�k|��7��8��$�riR"�P�Xh��`m1�%/����
�}�}-C z~��Yl������]�ܖ<�9��K>R� TC���-�f�RZ:�D��eM��3|b#`v{��D���7��FM�?�C�Nf�L�,T��Dbz��kc���4f����<���BZ��a�C�=�0(�յFk��¡/�P�e��g��d�8���x�����ql�XRմnJ�a���7�`��P �56��)ut�Xg{u���<��_&���x9�Ѕڑ�E����zg�?�9��~$p��
E��,r��O�o�N��4CL��crׂ6�;�o�'\���h��@}H.0*9��&��Ȑ�q;�C�M��������YDj�ʣSݤ�$8[:�%�����Vx�5�``�`�e'��;���{���M��+�o�ڴ[����l����\��*�/UI&���"q�M7^H��N7���a��2��T���=_zx�U�'5>'�0�姪��;v?>I�EWk�%�6~(k����J�hV	 �F��
�}�d]���]��h�H0E]��g�/;�<� {6 ��zT�tT��t�`T߭t�8|[N�ĞH�ڟM@�mR�+fWh�ڠ��nA�`ڲ"�q���;%��
--��0�z�}��p�P[��5Cg�|1ء�2�E6��2�)�id�A�d�9u���[h��	,��7��^��X�"�U��~�d�	�;/ҷ�ՙz�`���ݳ<zC�Y��*7~�^9��ňY���s����"�p���
y�Wʴ�i���Tf����|B�t��U.쿬Ç�&�2FH]�Cd*��h�i7._!�
��yg,�X�y5�����Rܩ����x4l#h4h3y��Gx!?�@m�������V[�bB��ݦ\{}2�� 7"\���1�S������#,ߑ3��-��@�x�Y���ڑk�?f�.C�NXt9-�&�֔Ŧ]K�ò	�I���$F��nE�b���XВ�F$�����!GJ�Oǁkyw�Ń^O��!��Y��a:�A�|�����sR�}�R��rk�ۄ,dA���_5��m,A����uW�d{����iJfX�E��f����yۯd�/�~�`|}��q/8Ř~Ҏݠ��L��ؓJte�a\M�����3.�	�py��(�|?:_\d�$��cn)���" n�RxL�c�+�C�J-�rk������p�'���bJ(#5&�]QI��DoO��o:�ؠ��f=tii[��Wc�_qK�,��= !��*D�O#�.Q�8_���/�oخjN�utf�J�"ۭK�����lU��C ��3���z��x�tA?a��f�gt��ZK�X�%�����%w(�bk��w�&�x����k���}PP��X�x?�R�����_N]�tR2,��\�*��(K�Q
Rh�MEj�b]Ϝ aV�ѝ����@��!W!p����Q��q�Z��Y�HP�(	�ۆ�P׎��E���~�%0�@����=���#���_�~�=����>�h���>3vT3A�Ct�p��<�M�>����&!s�f���:eN�Xdn7A�jq׳�[�:�
�#q����~�:��K��y���e�������N�!�� ����Q�(X��fjil��RI:����y��V�ˈ{���>��9a\~X��q�|@ܼ��� �I��D�@.<�a:�+���2��� Ehw�LV!Q�'�<��O ﯠ`��6� b�S�����L�Y�P�5
�oV��V��z�cR���ZsK����=]�}C�jL�]��q�+��(G�������ҍ�\�J�se!���^.�$t8.��gq3�y]DALDC��8��&p3z�&���S�`8���Px,��R"�t`�d��!�}L�z�sD6�t���_������$?saY�嶚<�qȲ5u��\V>�j⩅��>H�s�*�.T�J3\��Y�H�/i�`?��۠�Je���3���tv~F�K�f%e��T�vݨ���xO��$	C�t�wl�}�66�Œ���>��#
�?�Mܢ�¡�0���xp�a$���n�/��|����\�N��gBj�&��.��=���Z�a)���)�X�t�U~��O����ݨ_�+����<DI�_�%B��x�]7@O�ƈ��	�¼y�E1i}���(�oM�o#�4
���-$m,MI��WJG�Jp�p�J%�x��n�YV��Ƃ�����~��]#�cǞ��9��S �D�'�+�4',&js8�41��ՉUhL{j������k���w9Jyx��Z"�MR+��\���l��gKԸ/Y6�%86�ԧk����Qaލ�bZ:�1�ش�ρ�h}\�z�p���P[{�ֆ�Z�k��s�~R�R@�Kr�� tb�=��$z� ��B�'��'������L:�O��j��w�����i�'���j�:y�)�@fe@��k�rRJ���� j`J2u,�!lM0���1!9ʮ��,�\_b�Yz�.+X��c�/��g���<}��&?�Q۷�y�`�	P�H+"m�<G{��hȳ�����cH:վI�� U�JiJ�
EǺ��s*��יǡO�H~���ʎLH����I�A;U�Bvƙ�ҕ��*,b@�%4�+Q�!�.uq����UeJF�:�gw�;\��p�MZ+�O�Ѫ�
���2B�ވTsa���6��/��x�~/��C�Z���˻��gz�%��a���#���7�]+�RU)����&�Ƀ�}��%#�+,5<w�{I�3j[A�OBs��<�Dh�����9	�y�>�x��P����t�+����t���
��!G���G���l����ly�������,�H��-��6�ޫ:I�E[�D�'�K����o�B�M��� �;8�ښ�2/�W� ��+���|7�o�ۡ�%p�?�@0 �z�6D�+�x���j��>��:��[�E��F$gk�؄�$���mUU��kb� GF�|���B��T�E��4\��+��<A���_o{��k�
���1��e�ɠ���<������+���7��� �p<.��+��T�fqMX�nL~[��7C�=���1�ߕ�XRb�Wi*�.C��}I���UH��`��@3n�Z�Ɩ@��ͧ�Aptf|�(��0�����|�+�H��f'�C��Zu���H��o���f����ꊩJ�/��a��,�H�9���p�;��KD�Q��Ol��fy�E�sPa3ۘr�栎�>r�&:�s��a��e"w7��G$h����s����e�[���'��ܱ)ʇK� �a~�9�G� M�߬FVW�R/h����[Fz"����(nan���ή�^�WYd�. )�Uh Ҹu����x�w����T����f}��+��p�%G�c��dd�I��h���8aEq��kZ�8A��5 ��3�&�e��|�k�JYR��-�nA�U�<���* �����|�6�?�\X�wa�-#��Ӭ�%��[��_G��j@����L5�pB�wg�xȉ��	�xӖ�B����dy��v��P\x�ġ�d�{T�_��l2c�P�.{y�Q̒�&Ē:�g)t�=p-��~ɭ�J�&6��D�n���������͘ǿ�2*�3.)e������e򺜩��E�X	F�(��H(+�,6�����G!h�?}���41+
l�T%�U0�Ȗ������L>j��ܬ�n���Oڒu���Vެ�)��٭%��3b����$�\���Y��d�p+�?������v{N��i-_)��;��l ���rdL�+҅��3r4��գ�7��}�y�G��|����~����L�j���z!��7A����7[(aN9մ���˭���+����ɫaBj��!�^�u�ZOI_|� ���(����P Q���,�JDr��� �=�����ϝ�HG+J�����/�h�ూ(Zf���cX��g�!z�2���iK���w�G�%�Z8hA��)!��}��������L lя�� +�9����N�aZ��n�P��4���픇��_�	59<��P����� �����kjݏ�-�+�(T�G�7��XKDd�C*Z�bꩿf
��Ec(D��.ӱ��0���^�ͪ/O���l9�1�%�Q���]'x�s��m
�_i}ua-K��o ql�͠o\����^��9�g�K���:^3�>\'N� ��YT�=QvQr!ZP���-�:��Qy�C~��Y�:����L�6�i��C�{}�:�j̽`�S�Ǩ����g��� 8��2�Ǵ���q�<!��Y������Lm.����}� �o���N�ڸ{.9��F��Ą�it%�}{�b�i�D�,�}�読Q�=ʶ(���8���K��|L'~��ps�=�k�%L�i(�# s�@M�m��䝮8�Z�cl���n${��i������L��A1���׾k� AJ�x�6�b�(%�x�L��B\v~�l��yz�ʤ�s>�c��G⍬��'�Zk9"�<�<����)���=�Ɓ�ni��l*�v�@`m��Ɨ��G�Z��M�%��%�Qʃ�hEsv�ƽ�R�[hCR�Z��6�	����Ӱ=ߔ�ŉ���0���{Z�q(�m80ґ5d�9�2M��)2��X�5��<�n�pM5s���]�h�c+��l��# B��=5��>��jiT�̄�'N#���4�xu��StM�ϛ��~�B��;s��5�n�؎
̄zμ��Z,���ӮJt_R�o��'|Z�_��
��d�`�Uh/U�|ȮT�A_��i��ױȤ .��y<Bw�,�}�"���VF�"lU{�x�GB��)�1��l���4f$GS�~r��Υ��-��� �<dfX����E�7�4L�O�"AV�U>U~�rC2j�F-t���ߑ��'iQ�7��X����=����'����"�#���w�'��M����y����KcwF��A���� =��㞺'��\(�+$�_E�#U�,D?�#�-�zu^�ڰ8��%����P_v��-����7�l�ϲ[������Vx��L��xk�vm�5ظ�IO$��e�f���agz0{�6��\�HKG:�H��uM�F 
�'ܘ�i�n�AH��ˢ��>�(d��4���?ׄ����̇X��>Đ�?�Q���{Jl�:=�sɧ�^g�D���?�2j֥w_�l�*�F<�� S��~���0lx��bmH�K ';�'x�^
Z�8��p��M!l�+��bE>S����� �o6�,XF+ӥ
m�kqb1� ^3��-C�<���k�#�#f\�����|I������J\�����bZG�A������wv���F�Lr>0�)��?q���T���,�A��>����=��^��	:�c;��0�ԡB�G�6�X�#��@��Gۋ#��Vj���K�����P������0����h{�,z��1�LL���j|/K���73~�T��Iޫ��~>9��a&!Oɣ��ur���&�RP^��IL;�7-v��BD�=n��Ԑ�	�q�o����
O7�V���[���c�I��ĬɃ�~Th�+�Ϧ�0kC�.+
�g㮳	�7~�Y��}֎��S��GMq3]�dTs��pHM�De��Mn��L�n�����$��7�H�w���[�B�I/q7P������@/�u��0�4�Ԏؙ.� �������B�];����Ё��6�㗑�=�x1��F.UN���M*�1���%Θ�2r̪/h-v�;�wT��i�=?����@��^a��	={�ב���=�49N-nW)Jg�6Y�+����|w�/�?����2��O������6	ܨ�g�B�����V���N�&�!N��γ��t]CA�J�a�gcF�Z�yی�WA�`���m_��b����뿈P�ܓ�ҪO��:

u��
�t���������D]�����@�J�}����'0�S��&���҆�V�;J֞=���g��$��Vd�7�`�V}��6��a1����z��������rh�Eө'��ցi��o�-M�i�:��3�5[�{����SB�{���.ڊv��_�.��	�yq����~�
v��Io�R��U��������w�b�K0@t�T�x<;����fv����'�� �/��/��ĭj4�K���Q��Z��:���V}Vx&��1�تb�	F������8��U�C�3��t!Оa�L�K-�������
M��շ�R�g�I|��s���M���ג	�ߣ�Y�W9���� �ݜ�.�ݕ[�iB�����k����QFZ��Zqw|�Y-��Wl�}c�%��w�j��q�-vl��D�T�+��B�<��C<,��� ���
��KZx�)�����f2��fQ�F[�Ӫ��{�o��� �[�!�`��k� )�c��y�唣�:,��k��-�g���L��Yo?�Fp�)f&_ߒ�W��Ơ�V��41np�p�@��Qe���Ez@<�#F[�[��_���r�����0�?XM����"xc����<��H��%U �:XFU��)����S�z�]���}����=:����,���g�TB����:(3�˶ݰ)���(*o������L�UYfp7�ͧ�!���,O�l��r�-�o2	r��h%mn��;�?�?�۵9J�����JI1�՚Ֆ+��]�F�n�C�M�ʚsQ4��p;� ���ý:�:և�;�%#�[�FhRӺ>��ȣ���Ʉ��q��h*9�g��]��%|˪��EG�ʟ�װ+w���h�.�Pj0�N�K��E�o�ϴ	T���L¦xj�5�ch��X���"��o<�x��}��t ,�	��'ZЖ'�i�=�-��&���vŷE�K�LW�����vd층�3-� ]�?%b�<݌�H�B����٣�J�4�����]�H+�~A�z�Fl���xM�BN���i$���=R�ҒϏc�-�nY��)����j[�1��#[�֕��v GΩ��(s�>�W(wʂx1[��{��Q}�8�V�1�x��n��m~ӐP�ʮZ���j��'*�ZI���jrOqB`���?~�|�ݲO9t�Ωǆ]�
��\�RT&/����݀�����n@�jg����*U�!�h�E�>�0�2`o����'�|�0���A3 ,�C�ѱ��gm������W+("���G,�b}��
P�P� r�����c�b�2C�u_��M�^g�sj
�L��<���x)VV��Sd��X�����&�wc+�86�M�(��%�cyL�^F�Ng̞�x6/<E��H�3���y��WqD�;���a�$`�Tx��v!@�;j^JN��&'2U�Do�,��� �"6V���-�:K�#���/r�������m �"P����Y`Yu���9���-�=��l'�t�N���
�^,��W3�H����ߧ�]�BW��;�v:[4G���
�L^i'I0�`�yH��?�4�p�����]>���:�h�\�����J���;����M�dv;��K��/�\,���2�e<���q��q�W���#��3�XY�9���A�?�ħ�Y�.����5��}w��Kխ��_�UkUg�d�p��d&40#6�"�:�mM�6���L!�UF+<RY$�y�f(��7�[f�(䈟�����D`X�~䠎��()����B�X���|ID'�l�,�B���\hm~�ϐ :�FN��y%F�M�z5�۽nY�g��w�h0/�x�s�Eׅ��) 6ę�Y��'tO��
3��B~i!㹥�RYВ�]�G�0vJ{_r��S�P��)��JRs#�̹$R8��,�D�lG�( =��]c�����5�x���[ɊvǮ��t��s��˹(o����%$�|
�0epn�W=\�zb�\�?U�]Q�{e.VJM�"2��h��~خ\x�M�T����7�!��.$7���$�boF�ԬKau1<(10@W��@ ښsn+]�N��{��5�t=Iw�c1��th�~�U`�߱�~�^���Y�姃��y����אGb���N�ĜI�=@P���Σ5��ZIR,��hQBۏ����Ok��k�!mYw �7N+{7J������?�?sg��)�n�r���y�N6o��|��pGy�N@��� �ю ������*��$��!������H�LI��P���C�[ڰ�U��}frؼ�j=g�)����]ֿ�Ђ���~Ģ��0G����a�A}#tѭ 8�b��?��6��;R�[6���|Qʆni�  4� "� XTIM�Ǜ���|?�N�Tۜ~VJ�P��^� |�y�S�jc߀k��oD���g�9oH�xy@�?4�t{|�*�������dF�'�O]{�By�A�� L�4���"���ƒ@�%� 6���F�?�����G^9�PQ>N9��01<'A�dy�dT*u�������> �� ����emӢR.��g<lD�����H��$�2��L.��P0o���0V��d����BZ��f�1���G��y�D��*�rF*b��?l�y&�s#�E���t�l�E�ˎm��ך�}\�� ��H��������h�ɮH�<�@ɗ+�������ʼ����+
n|��l6�G�OjbJ�zΔR���F+#y#�%��9}<���D,�薠ݔ���K	�W5o��?�B�:��<����q���S����S�je��.v"��R���Hy�u�0�˻λD�t��+tX!5���\N<����p�շא�����D���z�6#H�I�zH	�w� y�w�ڝ�]Y����:%r)��8}�=:����4�r�
;��|�'���9q��f?����;�\>x��5�䞕�0Tuv���*^7�/��۰�h���{����M'�LH�	<�G��XPE�}!�F��x;�EtG���&-��E�P��tT%F����3鏩u( �y.q>Ǒz
o�M~��i`�m� �����㟺*�*��,B�IpX��o];7�(�z�>�=�Y_*�������������nv7��!�����D��_^1U�'d�/��XVE���3i���1�dt~����}�������%��c�1�8�7�}�y�&�������5w�Vp�H���Rp�+��]!ZL�Vi��L�7[�4��(�V�����(3ژ�r�~4� ��!j�q?�KT�ܴ��t�5�y�ӽ�rkލ�q5�?�ӗ~�n�ы��+�N(*������?��4�	���9��q�G:G���QJd�����gmɢ��Fc�RG�nm܏�Xi�Q⭣;=��ܩ\ί8��<�O;ar����61^����]�K�<�l;��K��?��J�������a�v�x��!�t���Z��WM�R/8x�ǃ���(X�8r'�;>�6�TY2 ]y�.��	���E =��GN\��Oư)���D:�B����1���Cα��t Яk��J��Q��%�P�V/o�EV�l\��z_�S�m���L'GW���ذ`�� ���U{�l��.�9;�=&1� �)\��3JM����mUҺ���e�j%`�1����n��ǿ��_�,���y<���ۼ>Q��(�GyER��H�,�Oer��c�@�b���hi�.�A�w��m�7�靡R��sTX�xhi\zF^�m�� �����)(�ħ�U�6�����N�|�4�b!�&x��}e�[!���0ZP��~E�7�Gܖ+��V��%2)M�)�nm#�YGz��GS��'9
t jŞ�k�x���%�aL��5|���aH�<1�Ɂ�~x��^ѻ�-w����8b��U���&Vi��㫴�¦���c��9�W�(Aߺ�!�zf�U ��6���R;��9�؁�����DMP�q�]��~	r����;�am��SE���\���*�ąr�?��:>�B�,��i�	`)uנ�����ࡪ�{��9E���^I|l%\��7��{�\KE��	��_T}�S�޹�X������m�EU�7�ϪK��2��';$sR�k���D~n���0�amQQ>��HgkBֵK�=ӱ|�U�zy�/Z?P/��P�Η�0����f���G�����f�,��(wY�O9 w�{����9�q�ݞ�VU�q�K_�\p*ՋxRg$�x�\?��x�@����ÿ��V��\K��0`.H7��w�g���bN��&�`f{�Q�R� �=�ូ�hXq�%�C��(y-�_�س�࠙<.��0�n���&� ��
r�>�k�G(�-\�Fn���W`�j���rHc'�"#CI��f�;A��*��J~�cAdu���O�L�,�u�F�$$(���!i�)/�P�V��>�/����1�ܑLڝ����<�������~�*$d7