��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������-��
1����yr1FUb��q�ej�IϢE^U�nA��a��"��� �AMF'�k-���޷n;m�o�}Z?��$Ĕ��L�h������g�Y]�)�}�"��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�?2zֺ�i�UCv�~��t_.> �KX�d��@�����O�2H�%��
����)�j�6�Q�؇0��E��:��r�;xՐ�>��~U�Љ��ӎ/s{p�|2}���/�&u��y�4�蕵���b��\�������Յ(Xî���A���
��&����h4�J	�k���F[��{����G�l��ّ ��t���3��7�=���	g�%�B�������4��/*�,1U[���_���	�J��pq'��4;0��^��ȑ�G�^k֞�٤oJ�\;ED��*��Pl�F"��}!��^��	Jة{����j^����%D'�H�s�/S��t��%��~pN>���Kǉ�{�������+��}.Q����|��Q��a��P��3��/����j���n&�F���{���b�'�Ji��!�h|h�Y|n~Ω7!&�}bd� ��g�kT&�"'�$�Ƀ;o>0R(��^> d��l��m�C#9cZ	�y��Gl�����eK��k5دI��������u�B�2�d8�F�G�{���5շt|yj��E���Y� k�
�Q�ȭ��7�B���f���f>r��7'Ѷg|�G[�,��Z\�C�Fc��iWss'\E��!9�LB�̍o�����S�lj��K����^]��~{�1��������3�&W��A�r�IM|a8.��(���'=Z�}���(���ԋ�3X��UI�N:�W���6�gѪ��ai�i��чL{�U����J�L��"���i���@�S⥔�K���S�8K\��ݫ��0�9��	L���DK��������<>�h��\l�l՝+��1��t!�v��_eS?hz����������0��hf��@�:�&h<��;���?��)-X����]�n.�����Le:[�|�{d�`4��9W5�k�\Ēs�we���f/^��.��ܛ��G@JY]��T�!��Φ�#���b��*�i�5�om�=�P9r�K���Ȅ��4�5���U��}�n�c����CZ��ɇ�T��B̕���84�<�vq�GC?=x�_X�Q�\9v�L2/��t��öCN�Q�Aw#����J��E��������{�[>���<�j��5�(Be�4�0��+(0��{��lz��z°���bh�U�	���L��z�+��9������]���)?��!����������l����rx�8��T�
kT�z�ȺK�M�e��t�����V���#����!���h3t�Ҙ�]��J����Se&��~6�>�~���W�	!`g�i/͈"�췐n�t�ǀ��_�j�D��Uw+����H�?N�Q驹�0ؚ���=^�cwȱxy��K(yvM�j���?1��)�x�_'����������J)v�b��17TiJ�*Ҟw�_���b�3n͖��;�v�<E�z0K94(v�*n��r2_��3I�d{��H�L�9kU �����a�o��h����!���Ør v��9Ks��E�uˑ����!{R�xj�K�Ӏ0���:�x+��./��Y�`ĩ%��ALR��S�D�\���� ��"�f�ػ�8��Yh&�"�&f��Y3�L��ɥ3��<�+�'w`���/:úu�t��G�~���(ʌ)�,T�Z��?�ޘj�Ƶ!���T�)�	?�|Z�x����.�_�	nʊ�iW�諟�?"��=wG%�Y���=Ǐw׼�����7�@ݠ�<Z+6׮T|���S&OӧX1XP�h�T"?x�����rx�lɲէC��a�肤�ND6�`�$�4J��0D2��7�4�����	ƘV⤙D0vW�Ǿ��ݿT�Y9@[�c�EH�U+ɫї�m3�]�ذd��+Ձ���Az0N�$[��p�9�zrrww�K�3�4vb��Z+-�]yj^���^p�d4�
ǈp�Y�kjp����]W��9k\K��ͨ� Q����d�}M��P��d��v��{v��H��5~�">���wCy��җ6QP��|U��]*�޷ �o��p��ĸKd*����m� �UࢲX�^���	s�3*��d`�t�^�~��'����>�& �
i���\�+E6�Al�rR���nBZO�X��_`�3��u�}��B�F\����PF���dP��4}��o&x��G�ߖ�x����ZC��I�+;Br�Ō�I�L ͝������$��<��#N/�y���ޒ��YN��W�(�����Yq� �C��Hy�з���tW��?�Tw���T�7R�'���%�*Żھ�񏅶.˝�O��p`�����u�@m�I�fr�<G]&�~�]x����ōF%��j�ϖ$���=ô�G�k��/W�`h&����f�Kz�.�9����F�8��n��}2��wb��+���b�q�[�Q�����!�ֻ�W��;������N�5����hCyE>U���{~3�.��tH��1����.sj���\�Q������׫	�LI�XK��b`����4ڪ ��H���0����,ەMu"2f4ś�RS���!7�/�`2��Z-g9�R�_���i�Dvdcщ���+�\%�{O�"��r�ܰ�h��n&�*x��*��? �0]5<�[W��g�t���,��y}�.��w�[S�� }>l�e�zQ�F�+8]Bۇǵ��`uP���a���T�N=ޢ�<���AQQ~4��P�j��c��f�e��@!-K���,�Q��1����<��fΘ~�����艈F�-Kl��K(�-l.�°t���t	tp�cz�ݗK�2�G>q+��D'n1�eS۰[IP�i@ �����j��@Z��0��	]<�$�!�(��N��k}�9���]�@u�W,8�7i���5���(��vCOwEo�����\&O4��S2�/h؎.��r���nc���˜�&&�nU�
]��^��B�4^[�	������ι��ɛ����� ��M�%����a�o��T���B�~*{u�Hr[�K8Z��\&8�&�ܚ�Nފ�]FCP��t}!퀝XC�^�:����:L����l� �Z�'�Ƙ��n�U{yjW�y�_#ћ]��B2��m��L���	���m����o�Nm�\~��O�x��x��_�1�s0�� �"L���#WA)S�o�Bz�m�S&�:ٿx ���i�_���%>�Ә܍R����.y�9园ԩ�k�/���YU��	4�<Y�;?*4�=��$�DԬ�I���O�W t�C̐IѢ�!��k$��d��[ |j��+d�3$��f�C���Z��:x��}�*H�VH("�iD�wQe�Ƣ���˂�hh���D��f{�_����̸� iU`�'��n%�(p0�����S�n���S oT�u�Tt��n��id$�+.�{�jT��b�7i�S���Q8y����$l��;�=ѱ�_&��m��ו��nS�1X�9KƆ�-�ׄ���e"~���C��A<��,�8��X��SmA��"�`vxC'�NZfآ\b���u�蠐]a�4^�S*Ι��vy�t�k�3�W�A� u��ɂX!4��J�Ms�6`Lr[u��V�F���]Ǖ\P��س�d$����uc�,�ϝ�E8?�l�mk��rc$1�{��>8���� �X{?�ʧ*��ڸF����� ����&J�I�E����k�eZzQ�-UI�1Έ����f��E��ѻ<EUM@��KqB�;�9Z���7�7K|����\$R>_��s)��[�7r{�K�ό�* UQI1�uA��X����NU�^'�p�X��?�(c��A� �y��i��r|�ܷ82����
Eؿ�pl3d�Ð_��D�W2�������;����_�X�߲'���� 9a�{�Ez"�'c*�\6x��B&'1H3���KZO�`ԗ�9���K���[�������]�kd- �ux���I~\l�k��l�Ʈ˘C��1�	�M���x��4�wA��g�|��ذB,ݹ���!�7�4:,��sii��%�	y��"U���>~>M=2��n��t��ᱧ�E*Z'%����c���7�WQ��am�,�au�>G�-(�V"F��X����4���׋e�i��[�]Ht��b�.�.�`�q8g�Ndv��{"��_�h�V����$s�b���稁��]�����`!���<YzpG�OC}ܵׯ�@� &β����^WE���S��̎��3y�δ]G�8����֙������f�A2�n��UN�ۼ�Y���)����9`�Re'�D����E��s Z����u�mH���+��_C1�&��� �V����d �R��҅��0'z0��y�#��q�G������y\ҿ��4e�7ȹx�0U!f��>�!��;�}��k�f���(�/�r�yg������Op��Z��}�/OkV.Q���hF:��2�N��X�S���#��S��"��K˥P�YL=�Z}��A	>�R=Gݸ7M��I�=ഓ��{g�5`�x,�������v�������x��g7�UK��i�.N�eyfY�=
�u��� MC�!i��_��hXy@���C�������]��V���C�q=#)����O&[2�&���~�:��I[|
�p����7�ȹ� �H�m���,�2�x~��68��bkFE�Ϸ0ʯ�=��!>�1�@\���>X9� F��G���Cw��՞l�e�x��^���!��\��[H�3w#�4��;u���bёD0��K�Mk��޷}���*7j��t�AZ,"���R_�!g^�
���B���)E�#�G��$�1?|��HO>s<b�S򋩢$UP0�B��A�4����]h�u