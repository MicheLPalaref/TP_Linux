��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�x}��j��S�b_�)F�1�(d'Â,L.��ꙺ��e�˭'�{���)�Ilf\�@,�y��Z�n�X�D�P��c�����=���]Od�w��yD.΃��o�N�o?ղ���	5��P]���t|�՟X)�3�׈��U��1Z� ��~
y�k�-�@pSy>8�Xy�T���2$�\K��ޢ( v� �r�s?W� ��YpH~��-=�R7Zc��Z*
�}Ӱ���]y�U����ʇML�D�Yt�a��!z ��r�w$)ߊ��h��M�W˖T!�ID�.���Ta��\kna��ͩ������
34yƸ�UdK0p�֨���.[ �8o����[�[����mڄ�j��� ��B��.���)N��x;�~�Y�R�%Tz�	[���Hz"�iƠ��9��vT#�e4;E��C�t���Nt����1o�w�	�3ا�����Y�S�l-_�!�3�8�	7�g���<2Á����"@�KR�M�I$Tu9��-���a�(��Qzɦ�{sb �k���-�Bڹ��� ��T��I����7�q_v#� Vi�)�Z�D�Ӓ�J�!�꽢P��3���Py=t4s�`\��%.��J$쾝�{cC.�P��@��{�����X�Zۉ��|6&���W�չO/)4��+v�IrǑ�'��5�T�p��f��v�'Q�2[�F9�`㺘v*Zڏs�D�#�<��l���o����	�M�S��$ &<V����jFW�R�1�H�ˉY+�j�d괫w���<Y��щ�lѣ��16�����xx����S)�⎲a���{�TJ��f��N�����2	b�Z��@.mI� ��ѻ>D�F�.�󧊶�*΃��͑߮8����j�[T;C��S��W�������H��Lɺ������Ѹ��ۿ��P����S�G]�z�%�UyؾT����lb8��1ݜز�3L����
eb�N�[�s�_Z���2xV4���[�%��ux�gt���h˒Wq�yL�	OE�Q5E�(/cܻ��z��r�fu�r�	�N�i9s���\yFE$NҒ�L0b9��~	YQ���E�6¦�c�}$41��'_��O�kn���%rXf�E�@�Kh�.4���2��G��.X�E���Q��W�n1(V^�V_�47���yv�]�v�c�!�)���D�	�%@�=��ܯ�|P�b0��,�{*J�~Ȁ���g�\���g�
a�y6�ā�K�G�A��:πx�(/�Y���ț���3�nD�{���2���V۫���`P�@�������h';�7}�v�=�$닷������c��+�����k�)i8��;�1{gS�|>\g��bUy�H�Q��6��n��R�mG]Ǿ�6&�k�ޗ���ܧ����x�9>7�K���AhܯA�}�sP��_����E{�_�;N��{(�J�roE��>�Tt�|��@+/&�N�%G�q8���KN��Ю�tч���"�X��+}���c��P�Gw{_r,�[�4	 ��vI�i���@^����5��(d�;k��8�5�1M���kP��Ї$|ML<����Gypf��&{H:�BLRE<�{Q��SA�G~���_�D��&�R��%�\#�l?���C s���p��+#��l0J�� _:]��f���(�I�=�.X�3Щ2mJ|O�r������a�C����k�u��Kr�/h���8A?�.�DE���>�&�>%	��?D���I�e=2=%��?��˿=vOs�gy��	Blͱ��dn���r��Un�|蜯��N%y�۹�dˍ�o�W@�A��E���ʩ��-�h�?B��f����7pL��=���-,���K�̓�z9�P��١�����S��ڷ�951��!�w}c��A���3y�q��\���).�Q�l]���٢`�Z�����O��*����a�Y��'�25�p����.���D�
�*�Z�e��0y>�:���ۅ.+�6{��_(}ݠ�v<ˤ�MP�
_Jǘ K-e��S$4(��)SR=�<-��S$<(��k�\`���'?1X,��B�]��`/����(;:��waR��m%h�}�I�5'�oR��N _������Efgb�rH��M�d�Zܝ���fVa0�^�=�lA�h4��xpU�S�_3s�b��>�e���m��B�b��z�	lm��P�g�a�@l{��2�����X6y��p��Hx�m�&�al:i\�'B�Ah$h��r
K}�:&^ ��U摞��1H��`� �Y�,���)�)���ٷP�,�mn<P�y;��H�ȕ{�`y�9���Q��A�x%v�6��e f�p�&�;*�t��ZB��B?����$)�V;L�A���1f��f���:���oFD���}��� {s}��V���C�]y���rl�A��%WLړėEu7����^�oԭДѼ]��tQX�|=*6�8(�D�j�ыF|&�6�u��)~>*��_�/洌��	5v�tP���
e�3�F��3���Rzu�d|���E���W6���5��lM9�sy����f�~F#s���g����r�#�嬙�6�I򘤩�����y��awޫ�Im;����h��Y�ǟƄ]زnt2'�M����Ur_�Ʉs�H9W�?�_F�%��0� R���b�g�b��v�h&!^+d����o�*��vDf��5���DE�~���Oe�F��cH|E�ܦ�� )w�����*l��>��h@��)��c�0R�T�x���җ�� �3�(�F�4Ȼju6]��U�rU�����ԋQ%c֣����Q1;P�vsn�5�gQ�-��������&
�~�l��7E՜�������f��a�H��>G �gr��1*"J������M+E�j�`�lI�lxW�.|%���m)��K��Wx��)��NwQ��PBC�~t��[�@��^����Õ���p"A#޿��Q]��i��"��f����4	�pgxjF�Z��;>�pN������E�����l��x�L��U����G�����+�oC�Ż�A�K���EeMIT��T3P�4w�ܑc�]c�i���F��O�n���0y]
چO��确CZvy�t�s���{�%h��8�������M?�	kAS~��Õ�Nս����~
�ά@(t�!,�KV3�Ru����id��L���:)$@��-Ȼ@Mw���:��,:����`]�vo�G���Sw�݂�ʨ ��ǳTQ)P�ꌕ�&Ԟ[�@0��;Ϧ��P��ӪO�?���Ҋ�J,@���S�$g��N�tF�3�]6n\��ɗ0�9m�ݓ|>/�$+@���+>��-+\���}�����g4ľ�) �@������ev�b����P)�}�N������#|���l{ĺO�S�Z?���J�`����w�E������߇��K���B�A�v6��W��&X몦���I��2�����'^���"}��;����ߗ5���AD�ܦ�1ΖۚP���[��2�����/�M�\Gx�F��h/4Uh�T�:É��t 1���J�U����m�g��Wz��7����%�!�ej:��Z�
շ��;���~T�Cv�c.�����>p���^�0V%���%� F����H�zl2�YĖ�7���!o�u�R�k�-����<�����B�*"�F��g�Y�4p�>`����_!Y=����Uǧ��d�&�����Ǩ�P����
0y�����}�����(U1��Ka%̔�q��#eX�TL�Oĩ��`��������M��m
#���R���X(����<�N�9�
&g������M���Ҥ`}�{U��#����"�}�}6S8�I�����\�A�t��լ�RyB�&?�.J�9R�,hc2��T����e8��ݟ�0T&���e�&�:5��8D�,����Cɏ��b��wd�2�4��P�������`�a�("�&#��"2�����Z�g�M2�c#�ٖhɰy�䛹���<��ʌ�PN
NXx\�C����ƾG(�t�2&�b��B��uJ�� hҹ,�\"�Ɍ����+��^��@�/ȟ?�Wo�~"{����h7{�n7p��0(��-Nb��i�����(B�K;��QD�����/��|��Z�g}�>�}���K+O񽜞�f�_��|�.��X���4�C[$Q�����?�9o��E��CH�� �jkc���<�t������N�� �a�/-�S�;ܹ��Ű
$.DC-����\5�_�fX?�7	��B>~����{�qj�z�� ÿ����X;w������T�G�u/aWy׬��
�,j���._;��:��q.�@�`��u��5��B��0��׈^t�Ze����7�t�CZ���:��r�[P(��z�����M�[�����߶Nɧ\@�����(�4�/�B<����'ʭskTH�0� D�1ং����c
�l�+�D|��ni�����WWI�Y/�?je�%���)\��@$��cۓ59��A�#����da�O�L�ī��b�ԧ��"�	�y��+b{����EG�5ү�����$3��kb1s����&1�BF��Z���|`TM��}ԣ�t]wڰ	I�ژ߬�b^���F)�rUHᓜ�}��Y�:$�u(���QO��� P�]�X#�7c�]8�آH?y�WA��b������_s��=%cMd}C����4]�p#z
R�i�礄�o�&� +�v��j�|�������M��fb׾v2�#��R������w
�Q�>���Q���-X�)�?�^'>�WP�w��W/��ڽ�A�a$t�u)�X���~�d���T��˖�OZ�VLKL\`�ō�/F.u�?A���G'G2�?��	�ᙨ��s��Qhu�F�H �Q I�QM�8I3D�&BP#q�:�����.�VBৌs�<湁� �xH�OX.I�]���|m�5V�/p��V$�l�PA6���m������ix��хe�cܯ3CF��3�]5ط߿p���Y�g%t�����kX������-V���q�79�P��F}��z�lPIH��.|{����8�(�m�գ1�¿��<{�SX�њ�X��?ˏvn�+M�G�$�t��W�B�Y�Q��0���qØ�n���4��d�dL?��}���Y���иcV��Ɛ��������πX�
��F.�D\3Q�$�y�j�S1����L`�Z��}F�����<�>/n8�w�	�py����Kĸ���- X�O�0������ɍQ���<�2�Ļ\w3��O+;'"R��x�i=�<��灀^�,
�\z���:�y[p�m�JGl,Q��D�hnӭ�/}h����H�
O7�	�-��0��v�_ ��Z�E�����q���Oc�&�p�B�6�r�����iG��3q�H�@؂��Vs�K�a��|��_��k���؎ʡl<[�J7t�Q������rj�;�|@F�n�����FG؊���Y��^[������K��~]g�ų��F?r�
.�;�ֈ�����BE�����y��?���������s$�
ӿ@��&��$���R�����9�a���YU;�l��=>&�
%�R3�#N�o�7εwhd�:�n^�7=�?�q�wv�%���r�dT��-7�L��٦��>��CWy3��t N�@0ר�gr�_��s��jW��m��Wk%�9@�DL�����8��5<����֦��u�h��(u$��s�4w͆
��43~�vjnA��>�,u��ɭ�J�� T2�Ī|�ıFG��G�g�AK�_ 	�pR��D��'�EX�.�S=�S�!0wZ%$�=R��2?�8�X�:��v|�5�@A�DG���T�Ă9դ*��'�E\���Y���Ϯ�H5����*k�8��atȶL�e��(C����5l���,�H�
Ρ�ۜ'o5���KF7#�8��ޤ�ؤ-Q��cZ�k;(�9�k�L��kʮ�T�+��+I����ER�G_�G>zq �*�H�L��l+����T6�UƄ�@\��`I�f��a�/DW�%�]��v�"-��_�hz]���H�$��{� {)���
�h�	L8~5��X����0w��bB,E���}�6US�mKk�=|0ݻa�?��_	��/�=�Ƙ��>2�=����q�P��^Z�����k3�	�ĳ'���҇���ϧ4Am�P�w�W��G�o�T#���Ou{�mq{���X�j�Dy�ޑh���?�H��
i,p_�G�[�j��z��8x�U���溤_���oP]�-��_s�a	3����x�:�<��ڡA�/\K�E5�{���h�/?��[�Т5�`�R��@��1���&�k��H
�#��ݞ���Y�xX����q�����w���~%Q��}�����8��)�0[�]D�����T���c�����ˣ��K����ٗ?�D-jʹ�����SϠt���U4���]�q�N8m��`�p�0�Cu�3����~�y����K��d�Sg1s������Q֥���&8�,x� d��Σ���I{�ו�Ϩ�8=Ŝ���q�.MM����P8 ��8G�ju�d�p��Dy�`C���KX��	�{�P�y��u�D�ț_M�2,��5���	[���tX7b�+� �;�r�c�,������Y
�H>D���+�!�۰o��Ih"�v��q�v��+k�����>�E�f���GH�!���� lu;�5i|&`�c������ϝ|���L��#���%�l���B:������I���e6�V>YY���Ɲ� ݆k�J!��;	�Ne�}�i����w�t�a��T,t"��\v9 ҢO�p�"��(��mg�m�_5�W��M��4�{	��;�,s*��L�OgLJ ��8��M�~�nX�2�.��t+2ҥ- 8� <ܽ�5���
|��@�7���@<t'�n��`׎%/�ѫ�`����ǽ���@�����/Y�@�-��G�WmP��=URd���.
�v���9�a�0���ѣ��ֵ��f�sD2$�yoO�/Un0��Ё�lH`۫<P���
Yt�	{�Sp´i�٪�D	�!q��q�LE��Ln��&��U�O��~�Дu��ј*S�D�r%�4Ө���z:z��uJ5��*��D\X����ɹ�&mL WpXD�'_q�,X� �y���%���a�k*���5�c;'�MS�<^��1�6}�fT�\����`V�}�x��V�Ձ�[k2�C�W���E�Gs���[�d��C�e��RkI��h�4��M�mS���Yg�ʷnP-_2���W��S��=�oD���Y$���ѣ���R�M���#����;���-�\�x]Ў��iO� ���b�R�%���F��#�TF*�wdz�c�:�6s7��Fh�G|ac�$�V����9$�m*Y;�d�MN�������{�'pxT����k�l?��Kn�[N`��A�S�3�r�M*�Ȳ�;�M�{</�f������d���a��lw��wƲ7�0��{�fܥP�Z3ǚtF��(�9��$��t(�Yo�)	�Q&�o�ż	v9Ş�3�����O���p��y7%��c��Ӫ.��ޤ�z��1��M��U��L{M�^��Q�B���i�c:�.�
l��qx2Į����RA.�^�&�m�yJ�S�!�U#��W�K8�$6�jU"��#	 ��DK�f� �����q�CK�)\h�t׽�#>�M������O\�ݲ��t��l�y)��u�tu0/�$�����X}��*�4�V�	}�� ����
@_E~�X����W]ofƈ��jkc�k|>�=�_ 8��OU�Uk�����ЌFϋ��#s�<xȧ�i�#u�SN�Sq6�8�
5���1�wwVYL�+��>Y.Dx��'��@��׆w@A $�%x�	�������ǒ �|Ё�Qn�4㚲F�ݤN�X p�����5%��'��e��W�^���*%7�BL��li�n@^s4�k��X��N`�?��v�8�s�w:B_���r����c�P�0,le��c镥�$0SBg�O�.�7.�)�]!����y�d@�������hc�p���m6�ac�k\���З⺣
'�X�ABk�;�Lkѥ���+������
u߷v1W34[s&���ff����_ڢҼ˸w딯v #�D����O���gby�u�?=)2wg�W0V|Y���JFn)%G���p�vP�������s.������Ia*ӎ|Y�N#Z�V��]�5J8�+� S��Q�����߻��L]�>���i 8\�3��_�
NcDQ��C��Fu�A�gU�ʭ0��ZG'����X�"R�O�2^ΗV�GJ�c���X������<#�sI3pe�� ��}ò�?>ݟ�E��zo2�;��|��c�
sN��@�C��Gȁ����E�U��z1�-۟-�ݨ �*�1�����Y�w�:�m�H�7U�@�|%�/k:�^��9�R����GIQ,GU|3t ����X�M�U�x=���k��X��h��s5�6��� ��.��@p�&�ub�ݧ��%� ��N�c��j����>y`�v��2�X���5����3�L��������������˭� Wq���L�z[�;�m����KVr��-Z�=�a�1�펕4<�:)B5!쪺Qs���{w7���x�#s�R7	� �`�Uk5�8d6p�*�F	b�C�ZeIT�z�%;,�y7�.���[�(�\��k�I��Kj�E;f���f��8;W��A���(2a��uׄ��
�u��	F0ufE��t��}��o|"\=И�KMp�-/�~���v�q�#Wc``�Oj�B���{C����ℷ�/�9`�TC��2�GMb����G�ជ�����ۨ��u��_�p����5��t 1�'7��	<�f�
7��j���˛�p��g��W�ͼ)+S�/�Z��~,���r������Q# �C��U���z9������\r�ڎ@w4z��V3����c&�h�6@�HB��S#f]���tU�̑|�>�I9h=u�o�j�b�J؝�bƕ7�B[Q*5�������6��k�:XC]zp2��r�ڡ "����`~hO�v6��������W�?S�7}���t	-9%N�\��%D�'6{�ߺ2IU�9g>D/^6T����nb	g�ˁ���'����-��1��B��Ċ ��,8�c	��n�V�@��.%����5|�`�X�bS�����M�H�k)-�߁�#G�r@åʢ� 
�b�.z'���Q3,��Ej����	��>ذ[f)R���Gn��\�{e��T�15���2EV7Cȉu�F�W�0A����٩��_n��EZQ
_�E!V]��}(��50x<A,�z:՟�Ss��/�s0Q�Ѽ�WjkZ��7P�A��$����4U�Y�EA!HH�7�0�$a�b��'Q��&w�٥�4V�v�Lb�`��*�ʫy��P�.hZc� �UJ�ےE�ZE�J�6y@�N_�ś_���y���O���B7#�$�V&i�S���`�e0C�2��F� �{�JBF�~!�$M��4)�)�zT���
< fDC�<�>XsE"ʯ\��[xZ�*@����zq�ur �rˌ�?g��~s�@(�()��!ӽ�7�J��<@���M}���%�5�8��N!O�?�����]<�N x��m��`X��]3��X����r�=�o���HC�����;��~X�T�o�7������%S�u[1Ұ�\�:����xM�oGFl����(��'u�3e|9_@M��И�`���Y����̤0�ڮ�hR����e������y�<� ����_�̌t�ٔ �߿MKD��I����>�$$O^�A��*�X�^���^�ֻ9Հd�l��e�~����|n��Ԭ�E�P����T/���e뿗<ϑ�U9�"�֗���z�'��┭U�E�\v��o?4|n�0p�|&���k������M\g�^�L�ؤ�'�y��Ez���tZ���9h�V�䖏��r�����5��v�=&������f4��2�^p�ٱm���</h�����f/�G�l�X'^+x��t���}� �1�sg�Y����?�
y����V35Μ�a�In�RS�l�h�v��lh�� \al���UO��'xy�_9�Cx�ʨNj�5Ƙ��d�����\�̭7���H��(qC�m&�=p ����l鎱��6�)N�q�V����?*s�����}�OɽF�X`Gv\JO����# ��E�[��o���9od ��S� }wre�cJLM3�P�����n����E�����?���
����#^����z�=����U��Sи⾟����Q̮���/���,�&	��k�M�hM���DŠ�1�WA��}1 5�x�!�J���M�<����R��6-vJ�fqW+<�
�U8S'1�&�̐(Trg�ɏ�fCK������A{(G�y!����|=J���x��H�����-�kM����~���i�Ϯ�HݛZo�����]�c�w�m��6��'��j<i�<��0�u=��&�L���V`v�n��2�L��63�d�'���JE�pY˶��lbF
���|"�Ε�cg�7K�B�mN�0B�Wy|.o����w"��I�EJ��.iRs�Ή���-����2�_L�Y��b�#�!��e�R	�яJ��|H�����#�e��;1��7S�փjˣF�&���(_A�?�4ÿB�쑽���%T�kUR63��0'��E��Β�h-Kpo`����J�<��#��b�=�K�!�	�n�D�����cZ'�"�r�I��L{0��E��3�Ѯ�(�8�W�-��gC
5�O��ח�:��[��߮��9�7��$v��C�*f��mXVԏ��G�1K�8��Vu�foM�-Dd��ѴF��5	K��	��9x�g���90�K��6E��C�)j�W��a_�:P8�sufN���g\�5�NA�}v��T�O�}`�)7���O݊����cL`�ֈîr$���2R���@ �d���4<�'�e���.d�R���"K��J�p��gFzybF��9=�pINC�ZR��$��n�!�t��%��ģI�T8eWL9b{��y�6��7�=��4���l1;7�ӵ�h��?�'g�O��Y�c�A��/ex-��F�q��|���yÇ�o5���h����
�2�}R�@,��@��������~�B��c�v��5k	
���v�����%+���!�ԭ��Ϭ��W{PΗ_K�v2��#En�v�j���鴗�G	�$��|�9$"g�n�;���Ⱦ�@g��Ÿ�QN�����'Zt����r!���ql�F��Y����T*&:��|R�Aʓ��n�m�^R�]j�-�Df����nmc��Z��S�⓷����sB}2ʌ�`�/���jU����ǌ����0%	�F���y�K�������:H�tL�Z@���Na��u��$:����	@���g�y�/��4p�����u't�/Ub �(u�
�v���׋9�)ݥ�#ɲ��}$�4���@F7S}�|:J�~h>���
Ct�{ȅ�����������s
�	AJs�'H8��9s��<q��IYe�4T�0���o}�1y�t��	��f|	Vo逧b� ��0dfŢC����@���n�sNo@ss50eeJu?�h�S�y��Me����ҽw}KQD�[J�o���͡�n*���hD0s��.�]į$���>�l!�O1�yN}*��̚2Z"`Ni�]~c�~*)%%o.�$�B_���W�����N�U�4i� +d��z�;s��]qBTl��H��X��y�8p{��#�;���_zx4,�C�I��v;��1�1NW�K�?��b�^y�����F�p����!^�1/�[�V��b�!��D����x#�3�C%(��������'�Ɩg�?�֌_��vT(?i_���S6��Pf��yh#a�R�{�j�����ۅF.m'h�zߑ��N��F�=:��	�$s9�\��̌"dL
O�n`�D.ؤГ���z;E?���3�ʳ0Ġ��B��B9ݝ��*����Bk�;:t�U�H�j�د��u�b1�c�N��<1񰩭�۩����6EQ�"�;c�����Ӓ�8�.�G%��. ��:�g�Cl����:6��x��f�#�o��R���g�8�Fc�~'�w�|8�^"�.���vǫ�r�4먫�"�qF�]1)�R��K���e��! =��lڇ�um:J�v���n�]��g䖞�W�	�Q'��Q����{s:��8�u�Q���h��������`g!�Z�B��W
RK����Q6��5p�G�?K1������+��+���+`iw��}�$��	��ۈ5��c����wC,M����{�6���P���K:A��"�!߼��ߡژ��x��c@�ۀ��	솞��:�s�U��]Vݵ�sG5���t�bG�����U�	�\�`�@��%mh�C���Ax�#�iW9E�X떜ce��L@�em�flQ�ߡ�T}%���

T��Q���*����}��y���C�/(�y�y��%M���K��kB���,��sR�u�B��=u����(%��я����	�o�e��,���~�m�z��z��!~���q
�f�;Oq3aȱ�g��{U�Xf?��|�Ǟ��y� X�G���1�>�a�>^'a�-g�<��6]ݭ�᤼+��ҸL�OF��?s��g�3�Qu���k����4�����M8?���>A�V�~4����W$���l�t-��J�E�
c���r�f��
>.��f�	�i��	}�0Ӽ�=h�e���Z���
��ø�I�$��A�G&��u0�9�wXۤC��@C���=����Y��X8״o;`
Q%�1���>� `@&9�k=������:^{;џ~��j�$5Tic��ށ	RpIa�f��AC�@t�����C����3��S�̇�1�>��9bŔ������,�S�喾����JN��`���PRc_3by�U��y���Ec�,d���J��@Y�@����ΫP2�b�����LG��A>�D��P�#~�E�ɔ��>0<_�LJ��=J9���)��q$�WԊ�AsY��	�W���||�2�M�O�s�E>� ��%�O୓��{��1����g�����[�9��8����UHš�|�M��wnEΡ*�����C+_n��1��8 C:î	r����d��["����z�?6�s�������,��`�؏������\����
xBy--���cH���s�7�3�pG������17����v.�6�8�GD��P�d��Q<�}{)��"��H�K�,�H�S�C�
1���qe)�\��
u�1&DY�xd�=4�$p^W�R"Ūa<��O��!�,ƙK&�&6�P�~�w��㻾�ԩ�CFiAE+�F�vQ-}1�t���4,�Gf.!\�����jTd��S`�hK�l� ,�4�� ��o1�O]��`�
�:�u�^o�l��I����2R�m`>�T�Y��t���Q'{b������H��rN�0��c����M��w����)r:��,)�V�(���BG�{[�C���^o�wB!/QZ����T:�Č5p@K6W�٫��Ğ��ު���1�� �#L��e���Դd�	��ߛ0~�E��,AɡD&�9�j~O���(+]�8@�Z`h#){%�)�9_�#�v��y��fZ;1��x�?����Q�[�k\2@�ভ���w�%_a�����P4�x/���kN�j�.5���[�F�T=�uLp�^������R�e�?�U��&-4�E�4����b���<ҐaV���\@]�A}����+��_!X�q�b��Tu�yht�K�y)nI�5�%]V8$����q6*�[��Ԫ腣��r C5)]k�/���j�j~J8;S�_�I����xp���:ȉAC��{5?]��m�e���~������Ķ��#cGw&R���� �B��8Px���DJ��p�}�,vԀF<�=ծ�9^,d���HP{c��9mrm���as|K��%���˷Z��h��鶕�19l�`�N~;tk!۩I3K�M�TL����֨\~�%���`!o�n2��3؏X�d�_Ƒ����	o�ہ`A��Ʒ#k�x�WR�5J�˹��?�J���=��F��S���C�9���.�jAζ�*��W�5R�J�L.%C~0Y,��t!�����)�^3N�
��n�̇d��A�G-��Q�$̀�zΙ�I�V�s[��9Y��U6v,��RUn�z��ï�{��r|��70RI�5�c��Wo�WnsL�K&�h�w!g�VEn �,��1�0<��it��x+���,�X���c����D�{�E���s��z���3������R���3n)�G~��hi���ၖ�[ 3]�3��$�UC���B��_�!�n�Ik��X�@�g�4e����S z֊�CK�`Qu/ȭ�Cp������ .[��O��D��Bl^$I��v��Qa���8�uC!�9d.�V
����e]�K+���b��ԝ�pی����I��m�"�������c�=*	�Y�����O��mCa�ݡՄ��j�Oj��- �F�p<�|G��l�i�բc��v�n�;tΛ"�g��\�LG�.��_���/~�B�~2�= �w�Y۔��OO���+��S"UL#ja	��ݦi�i7:酯��R �
��pG.`8�U���0� �4X�h�����ാ���]#��1����}�\C֗�ڻ����O��j�]����C�P�����q$�<w���*��F�|Z�~棌�؉��R����wI�������� �ǈ�+��2�=u-qJ�t�S��gNe"O^{Ks��l�z��ҏ�,%H��r8"��� �m+1�A��ή��jL��9�j�Hd�aC�Ҳ��}�������*��k��U���=�6`���55�9���Y)����l&G^̫D�õJd��CB�T���Onl[j�ؑ6>C��K'�"5��Ѻ��EBr�x����8�޼L�Gߒ*�᭧�@�::�szL�UK�����d�>��a�����~������Zo�����/�%7��g1�.�������1�7=0�l��c��q�Kh߉7X�W�Bto�%�}"Kq���`i��"y����}�Df\;CB Q0�/2>9G��Xva�=(�㈽e�8�$�KJ�GҤ�E`�)��@����0`A|f\I�,����-�G	��!u���o��2DMyT��<VZ��вLuB$�O}h)u����s��l�^pݙ��;� ���$`�����{��Kbwץd=HM k�&�*݈z�KP��<��+>|+�q��k�c#���X�$s�M�'q"e�����)�^��®S�7�䓎��w��i몳�ޒ����L]���v	^*_J�J=�}.,��=�X�^ZS�1ה��\���X1"we�N�}`�؋g���%���9�XH�Х
�u�QN���5:*r�j
(S=�LL���q�DxB�Q�����7?�k�:�6�e��\��`|�X��19F��j�����*�+yi�۩�ь0��-~cd�ée��K�;�f�ɺ�\N�Q85cd�� �N�XBq�Q{�Ґ*��?fs܈���|�QW���D�a\A��C�;BM�V �ώ�w��8w�Ƹ�6g���c�\�����&������e�E#?e�㲧�������D�.���a��~_��!U^��_0/�m$��I����JD��C�X���\~���傋�8^��L�S��K����䳜�A�]��0\6w��$䲴fQ�@ZzJ&�YF�;3����,N7; ��J8��A�(s��ø�8�ڀJ�*z[��8����+��fq����D��wݲ�q�b����^��5�L:F�"+�M:�x<E��=�W�j(��
�O  g��h�=p��+%����G�j�W,V��6��$�*e�fpm�?�C�c�ɿ<��3�}Y� �Lagz��Tjl���;�E���Q�a�G�մ����D�2�tEa��ϥ;��E~�ε<N6Fr!���oxnҍ���q� :ĸSl9�|�Qa��ʣ�N������e���DC@�}�^��S.~��-���,|h��D�6���dMt5@ ��F�D��Y�I&���Ò�.HKS�� �SW��Tc� ��F�Ȧy��R=��%�'�G�T_������Q�7 "��#��r��P�xI�%P��j�!��in����W��
�x���v���=�2�M6G��6�t�Td b��D��΋cڶ�Y�F�E#ǲ$��CԄa L(������|h���(­HQ��[-����h�"d�`�,y�!j;�t�62"*c���t��E7�ⲣٓ�G�k��Ji���7K꽟?h<�cM��:��l�������h���l���"�ͬ%����PB�� �Ez�����|�ŷ>� �����#���`����g�΂��"��D�FK�ךᆷ�1Ŷ]�x����-5'��,M���+��7"+�l��M�޸K��t�	/,�	G�X�F�f�����@��HEW���r>d.�ǌ���G
ú/��z{k�3/)���\���|�z���/o�zR�F~��r�<;'j���A��۔�v0�A�4�}#S^�xXm$��b�j��=uN0����Qd�,��ˆv�Sj��һR_&������ݽ�Q�ҶK�c��D3��U������|�!��ȋ����e�H�w關Aփ�O�O���8�VJ��!/��l��P��](��x�7���
��;���O@�A�ՑA���Ӡ��Vy��:m��}hן{+��u��w�<%�JZ�������'�,G�/�h���.c1�_�s箝d�e���P�>�.26,��P�2�E�������4%�X�WMԢ��5}rI�4Ì�(`��|��6�t�?'��&��j,D�>_��s���w�K��6����q��Ά�cI!�~��ȝ�Ie���-<�Y� :��Ht����S�㆜�dt�b���٦�@���� E�60&�DLi��;�XZ���R|tl��oۯ�p7�Y����q�x�`�D<�`����f֠�)kp'��Oa��JEѪ��o�W&	0+��Q�r}��K��6v�F���B7��1rc-��|�s '4�	�u�q[=vhX7����z������4A98a�=�	�1F*bp��v����6o?�u�{�Ga��@��m��"�Z��{3���/_��ce`L!�D���Fr���h,Fp;#sl���K>�&�.u�+����V�o����!�!�o��Rg�!>'�Ʃqn(HG���ꦃ|��S����]�L�6�w��\�{nw{�]�t�z�f����f�וT$A�3����wO���[�'O��m�޽�'������B\caa�L����E\���7j=����~Z�Ѓm����
�K0uluL�c�Y�g���2�Ec�^͞qy�O�!�pz�o���ނt���nl���`	��oP�,�� ��G��ذ�}�$����NYm�H�]��ϯS��uӴ����;�,�b���lո�Fnv�L�|�K�d��:�Ga��y���"Y����0YNn%�gx�G��dg�"t/�4�R�=�d܅�F���֍�S��f~zN�S���i��.۝�1q ���L���̎�Hh��/��r<*(Xzj2~z;�,�U���O;Q4_c�.�L�y1�-�2���8���/�����]�n܄X��ӱ$�w��:񉳥�?t��dnl���$Ɂ�Py��|���B��G���9��Y�� �9O��n��68�#D�U| R�;����̥[	tR
a�=M��6$�ΐ�dgի���o�EZ�R�d�`�v�X�>&H�U��F�����c���rgLNSc�Y�nʲ�.�gت�Q�;
|g�Rӭ��'A��m��F��	��F�o�k����2x�2��P7؁/#OͰ��z +��WD�/�?[���^�*�?c�ewQ�b�&��Ow���͋�i/�J�u�wpU�� �ï�U���41:��J<WGd�ܚR���(�k[���K"4����LFsF9{��#,-X�>�>U2\��Nw���m����c~�I�jŰa.'��J�\z��7S���D���z���=ŕ����Qb��v��p?�3�@����(���ϡ��=��jY���j	�N%#Ӊ��_,L�
�/�����3����9��ɏ3Azֈ�E���]��S�<���[�]D��I�e*���H[O�n�����t~�2^��TU�rF~Bt�ک�ˡ\`�6�b��*�XȥNC.q)�/��X���S�����
�!��&X�<|��?L�>�E�	��}�ј��[��� :fŜ��]j����\��q �<��k�i�#���>��a��Y&��em3����\�=5�[#
�jUF�����끎i�N�Wg�HbPoG�%(���_hҹ��4\��.y��*P�?ThJq�#jC�j(ʴ�ǋMTL�B�8�2Nj�r���XB�t�
�x��ձ�Y�_���.�'C8c����[��no@���+�?ҟE3V�Gu�A��T�#�൓�V[:&Ov��p�*1�׶�~�[� ���!o���4)��U�22�ļ��?��Q��-�jt}A����|�a&|�S2�sA����.�j�& ����x�T�e+`{	�¡CX�&�q|CS#�dG�'j�C6��!,ة�Qt"MQ��G,�Ͳ�T	ڷ$Fײ�j3c�-��w}x�3��@P��O�PeJ��x�)ٹq���X���������3�L�SLfl/�6Q^�o;)<�XN�k�)������s�ԙu{����v��fh�-H���Q�S����^��']#���^����E��xY� �:W?�䄻{�t �fE�㴞�NmǨ91���L���S��)x�i.���Or���s"��+�@��2�fS ��+]�C�O�����'�2�Q[�\m�z
Aƪ��cN���_Ȉn��d��pIk�7"�K�İS���i��_�[�q����0pr�� R7r��^�8x�1J��@C����T ѡ��9u�ص�d�7Js��7ZCg��)3��=i�5Ȗ3�ly�Z���E\L��)����ǭG&H�������D ��5�֬N��LE�8a�\1�h#b�9�~��]��'�Is(�����u��U�R���ڌ�7ybX{١����}E�ks� v�EM>̔��ǖF5kQ�`4T�.��ͅE���eF�*���f���2�o`�P��Z�i c��ʋp�&��I�;���(��m̕��N�>��=��-q��6ڬt�Jci��_�+�N��-������Ocx#�rzܼ}+�I:�w�r�#{�k;@�C=g ��˝^�[Xy��IL4�+e)�_S�ZS� �F�(�vq�w=K��h!z���dco�g��
ɮW�8��ڐ���`&�-I��ਗ਼��#�q�x���&([t�Q�=�Nn$�h�nZ�K�n5����F<�Ϩ�?_3�2?���T�9�䘺�?���Q�SH-wfk��[5�gf��qv��yP�<�ϖ=�s'M͘���=D*����+@�m=���P�QS�➛�`X-h�e�ã�鹊F�V��$���Fv��P���t5�)�f�~�x��/5G3ۜ0`�ߎ�h�Xl�������� �D�������4����!E��h���C|�2RsN�=�G �,�,�?��%A�o�=�L�(��v�6V8Q���ٕ	�dL�!xj�Sa��w�@���t�&H6�G��ϰ�;>�Dr>��J`v�����6������������� �����g%���E���	ځ��Į� �����=�ws����������Y/:����8���:kwN��UF�* ���	<������]����d܊©�[PE̍/�).�0�:����0vlH+����Ù}"V���誴W\��E���,�Lm��Tj�Ã�m4��e���+=�sF���t(�cl�S~?y�s"��>]���[B�m�!>��W��SR_��Y�V��f������e��%��}

ze%��P�m�sY�<&Y����/�^�tF�������?���}���51���P�Y�L�G_i:Z�!�)e���I�j���~o*�Mڳ����L͘�1�������m9'^
���zZ�ʢ�[(���:	bIo�g�Tj��;Z��Q��2��ћ��P��RLı�ThX�^�;lk�pm��&#�6���Ym��h3��[%��.�wL�>�ǒ�����=S�?����z����Nb&2_��o��}5&W���l&���zr|q�J'�*z�?<J�;>i���@�O�io@���h�+z��_)Κ?J�X��?HY�B�2��s��W�8vɄ�~��]�i���p����Eۓ���K�Ho��6�lL��P�/���v�����ӻTt�?�[����3�%a�q�[9���l�D�~t
"��/Aw�7 C�?Kl��(���C�	早]�\螁��q%�}~{���b���RbT�ᖨ�~����i7����Q��Sy���臁�Gn+�KŌ�-�A���ug@��,�Nٓ��z�x�'`!EͲ(&��� �=wlSp9�[�&�����Yo&vK����w�~Ft`#o�e���)M������j7��nm���{.��D��H�a�	-]��H�,7_}p3����y�2�/ݾ2jm ��]s��`����:�+ܰ-��p�$$����l"Y�~��\l��@l�l�E&�D��pO�VPN�S�n��g��wl�ݫ���B��D��_��\�$�?O�h�t�M[����X��љT~�@�Z5�c��%�a��AMƍ������$��m��h�,N�SL��2�E4_�)���0���G�f��4Z�41n��f����Qö�#m�P��6�Y���+�m���ۏ��Y�����@���Ab�YJM���vb1F����4��?���j�%=��$}Si��z���0g��&5�˹�F���d�@g�^Ȼ�˚nh��0��^	M�u]N}j�2���&H�fS𥰵l�u��dKy$�Cj_`C�&��gA����d?�#��r��~�V�T�R`A�:��{����=�X���N����D��b⌱8b�����k8O([霸�<V
a��fv�؎�k=���ډjomgg��{��=�-�׸��nwg&�fs�o�;������*7�Eȧ;Y�m,x7�=%JOR6�1�H�Gq��MWi�z�Ç�}!�g� �m��` �;g���.J���*�y���H�EQ�d���2��ӛ���]hș��2����L�U���4�n���]��!���yB��M�6�=?o9�
z��WR2`��Ƭ��l�/eb��Â���q)���4�@ԋ�hb�"h���8�CA�9*�]dHa����uW�1�X��A���4-1����|`�4�Ͷ� ��X����+�V���S뱭G0�	���m�)�f��K��� *�+ZGm1V��E�r�q�DQ�Y�}�,�%ڿ�2��u��Yu�~�����-i�zfQ4��ۆ�0��/�<yG%~�U�{�J�8r!���=	���4�C	���P�%l �j�I�&�ש�k;�n��7�����$��F�o�R"�����]5	B�W~U�f��r��&�O/��pL]�6�
B���ռ��pn�r��@���\�<t�ñLA����������o�ZS�9f���6R�Ly���K��C��|}�r��W�����π΀�D���+�0�4�U(�C,-1���'�>u��Te��Nv�fn��Q��Na^լp�������C<!���_���wI������o3:*�|͚j�K)^|0D
��"Lu��T�vX��{v�Ւc��
m��OB��;�_H����2�߇�?� �M;Ͷ����!��5g��&�Ѡ�2�Ԗ�����4�!ؐ��Sx��ƺ.ן��N�M������$���a�7��hܥ;x
�KVu(�.(]���ȝ����������K������Џ.5�<�l��h�y0儫hoЋY�P���T2�4���sn�u_d��ݝ�W"g��?�S1�����r`4�꾎�n3���=1��3�"��,����G�0-t����x�0h�i��ənn�Fy��m�qB
i����@H����Q*�*�����3q�/����o��^B�r�=�ɣē���������\��v� �j�a�%8�CC��N`,`����a�Lt����@�2��B�N�WvW�ȱ�<6�����@I��)e�=�!2G ���*�t��}��jw1��0�*w���%��8����y������Y��k��@���t��~�)1ш,��7��
w���"k��ߡ�"28􋬋�;0�q+�Ht��v=�Ry 	��בW,A��=�Wo�X�����O�����}���\R.<R��w4���.��H��3H]��%�#�BS@��2��*�N���L�?�w���v<��LÖ|�Wb�k$n�W�rE{��ߑ�5�h�{t����TN��nx���?|�"�wL��L41�
lzd��Ri��E�?���ؠ	*R���#����<R��TJ+ʮ4O�A^EY�1:�R�- !�{�%{Ա���}���)w)���m��lQ��c<֗�D�  �SMaE��8;ki��
>���1x�(ڋ���&h"��JJP&�{���X�p���
{/�Dԇد��U���r>���_�w�e�S����[�7h7љ�4���'�`�֩�O}��i�x�&+��T1�\7I�&�[�-��a"��En��x�P��N��@��N�(:��u-�����@f-�q�%ox�>�����'!�5X����t�:���Z_[�W�$s�5+⃹�3K=$R8�c┻�ǒ�לD-�����t�V�h��!i/#όw��)��6Ň����D�5�<+��|�g�y��Bc�0���k����npmXs͈G�8a`�l=TK&*I
�E�"�C(���r���cxۢ��뤒p{�P1���*֎�INgD(/B��C,��<�r�Y�����S�.NV�K���X�=Q��8��"Yc@�i]��7��~�qg��q|�5��~[�~���Ĩ�7u���Xש�ɑ��vJc�]J24=�p{�\vطm#�^�ɡ�o��J���8�P��:Mo�V��H"�z�mO	�ѓ l�i�l��
}HA�[Qg�/�f̽�	�a�֧������l�Ѝr�WN��L�y�OwG��!&7�.���&n�~n����R"m"b��|�<��9G�L�-v�ug�e._i��l`K"�3ت���Q�����{���*:����+�j���Y��y�uI�[���\Xa���b^tƁ��S�R�ÿX�	W�L������ȳ�B���/������V׬��t:_N:D��j.���|���YHX4tD���WЫ
�$;5(��ȣbz?�ZIy���XTu^����;u�	z���:dK���`���@c�xI���VF���0�Ք��_UUFY�[�I������ZI��L8z�/y�s���䅦N�+��h�/̯�$��RڈO;=�5%���^�2�����Q]9ܳ��=�#�g|nae���"���F>1`8ξf�or7)رJ�hm����۩�m��'5��C�O���k��D���-�ʋ1�,g0X����=�i$Qf������PV��ٛDq��O�z'5��w�J%��S����>��`�P�ؔ���8���u�pK�c�Z��L�:�=�+����]?-Y�ٳ�