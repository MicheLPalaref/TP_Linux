��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z���$Gp̱`��@n}�D����\��D�]����x����@R�� D|�ط�8���V�����`kj��̢N3b��C~������L��A�T��c�l���~D�����ӘFy��P�1�ɂa̓��;R�z�tZl���k}lV���6�;v�܄a���ΎC�ÄGuM1ֈ��@t���̑?���$�$	xwj�}�G, uz� ��~����z���Q<NI����kN���pɎ��T'��ݴX�k�&j�g�P�b/�`���(ڤq\�Fc:�o���R��cYc<���G�E4�엡���dW=�{�7j[O�oo�\�#�xoH�����	�ib��;I�RdkR8C���F�W�J�	�Б�ߺ(��gW� �'P��e)�k��|^�y]VEgHkKR��-d��t�i�ׇ���%�M�f�R��s+��8{	̻�j!�G;|���Y���FR��5�l	G�m��-�k�4#��[n�X3�ѹ��Vq�<I�(�S�a�{b�91el��ϭ3���a���sE��p�����B���������	�|��C�ҭ��r7캪�O�F�A�0�-o�U��ˉ44��o.�|5�i�+��]��ʠ7Vf�.�Q����i���=�JѠ��k�R�Έ����g��be��9Y�=�3�zG�ozቔ⺗��JJP[�B�o�6Գ�0{�Ul<�6��*]?L�0| O\�av�-����=S��d�o�n>��D�W�綞���Ѕ� <��@�r�������Bg�wyb智X���`=��)�|Yf�;z��J�bjX��F�x�� ���K�؀�1��:Iu~[P���YJ	�Q�n".��N��/;��
H/N�BW��\���Qdl`T[]��/�+V��.� �gS앿S�\-;�����ճ\�ic_mӴ-�j���tݡ�嚑��Kv� @���iZN0J�)c��f�`D#�4s�*�$c�����j%_  �o����2�Zkc| eHF�����F��;:8;��٩��5��)�!~TM�ۚ�� 0.1�xfK��V1H���J�dH�k ���7?���?�9����ԭ.B	��d�w��-U�v^�);�-�4@��w�kyjo���_U�6H(z��<�}X�w��JN�L�Z���;�ct5!��zwV������%T��P� %:�t����@VV_\��Q��5"����Y��EܹD�U��s�,C_1e���?�S��>W!J��@�K�7^�V��}�e��8��+y��H54dze���t��[:�7-9L0�Ϧ�w,?��[L�h���g3x�Li��}�Q���3FO�:З���Ro8!�Y�܏������xKH�2M�%Z.��{���.s��_��n��ol4���cc�w�5�(�o+ю�]XPZ��E݂��ȹ��ߺ<���a�'5�������_61�8��\�u���H�;q�7��X#�XBȤ�q��Oϭ�0��C��%d)gʸA����ӕ��޲����]�F����)�!�h.��6����p���{�5�f��6������Z��m�Kə˫�2��xk1h?N-)����.��]:)l��4����e��.|���K�ݑN�IN��M��}]����8Z�P,�߰b��m��������+��?5jmRll<#���RX�5�@��g�'�Ҍ���֔��7����-����n�&>���"*|H��V,�W�u>Ӂ����$��c"��5���n�Pc���D�Q���6��"v�����8m�zf_�Lt�ׄAK�f��dV�4x�0Ǔ߲\�J6J.�Q'��0��8���B7�E�:���E�ɸ�y��Q�1��w����/��4@\�LXt0�g����M5�ۡj~��S��M�734Sl��W����d�1��\gu_q���h��r���Г6��@sݨ��Pg��}v�r�B�\�y�f��@���k*z{/�M<�����sC�4v�Yݤ@NbL��1�1Kr�uu�t��K�	�>w�)ϛden)�Y����$?��w�sIfݘ�Svǖ��{A�c�q���8��C��C2�*S7��p����C��.��o��Q�c�^�'��>� �D"�r��R.�1v���)��S9��i�B<�����&|�%��:篮�kCV��Ik�m�����uy�'ZW��������디ֱ�	��y⾟$�=e�DU�	�ּ}n?�ˆ�ڶ�#�C';��C�f
�9r�0݀T(p"CN��$X�D;TA�����U4����(3�n�㪤���."��W!�n����0�4�b|��6$���(�x22t�Z�!{�q��ݎk�y[C�9�M5��\��o��v^�q�T2쿣Kc�i�c��G���͎�԰ގ'�0$�X0��?��k���&b9�����U�1���~ ���r�2oOڛ�[�6>r��ѹ>5F�A ��Z�/�{i^��A����4�`zg�y2�]�{V<p������-�P�^�0:^t��m�D���I��<����u3���^	5�Z ��BM�U�l#��@b��l¤�TS�����B�F�t�_(v��O���m0�x��`Lb\�;r�<Ȼ�<�7����&qJ���e��^��E�߶��p@�&�w6���u�,�`���zE�|ũ?��c�DN?��m �����[t9p3����!���q�qc�~,2d��_*,�R�5�1��g�l��&�0�.�EЃ>��)�3O#�V�8Z��k(��v�I�3�(��񪖳��G�79�g"�V}���5��6��O�cOH���efR!ٟ�;벟k�f���?>�e�-s�vlq�,�1�hN��r�JXn�r�k(f��n��r��ă�!C�tf+YUG��b;����0���AT��V
2��cT���lN{�:����RCǳ�|`�C嘠�s�NXC�Υ�6of/���'�N��>�J!��c�&�yr��0����'��H��{&�ӾӔ�����A�i���t�
�=}{C�^���v�J�z�w�V��`�Ph\_>c��0�B��{�٥�ٛ7����o�Λ:)b+J�MS��۵x+h���sr�R��x���Ih�d{@�ed���x�d�*]O�Ea{:>梺�����H�����S����G�V9�}�Fw@�ŀS�Ŏ��g^��|�
N�X���I���]�K�3f�tf2��8[4���R7���_r���j�$�{hd���$�R��g��١i�쬍R$g�����/f@VDH��A��.�`�D+Ɉ��U�c�h�tk벿]RD̳�� �(�(j���X<3{߅w2���N�,���M���"*���c�٘ '|*�ک|l���_����x��c2�4���K��,��i��ǒC��ʴ��,�} JoP��ɍZ���Z: h�/�Jj�U#yڤȃ�ε��ϓ\g�2Z�Ͼ��)(C�<c�b�L:z�q�(c/�y'�=4�߿B�t��혗�p��"*�E�����σ�w�CV-��Ԏ�H,F�I�\�	�͡&�.ԓ�?�W��@���+`0�*1��	� ��;�g�q��aJ� �h�I�ř +ᱣ�Pe�I����M��Ў|���e������塄�^���kARt��T��mh��Ǔ32������aXU�����Ԭ���k<q�t�"c��=X�B�<e��y�������/nե=��>��*�%]�9��V�~�	�`���#���2�}���}X���'XM^�0�>��h�MQM���D�ysmn�0�Dg��"c�3a,��<x��@9�Gb�ĦP���@�'S�����Y�jq���j4����iހ�ýxLD�3Cv���̊R#���
����{���z�NEr_�{1���HV���(��	ӕ�]L�U��7n[�B+7�� �ً[bCwi!<i��0
��a���t�7�Wr-��o����Iiύ�R�l�	|.�#Xw{["��u�J��x�+7G	2Kڅ�G�&i)��ɦ��g
��<���+�$��'��v�ˈ^�!�Ǜ9Q7�ɛ���\�n+X��Ϣ�=Wt��K��O/��Kr��OGK����q����-��wgn�{�u}ّ�4���#�_�{-�/�� *{96q�R���C���*�.�i�]�,p��"��P�T��VS�\���ll�}cA��o���,l��F�1���3���W���8Vg�\aA�~�Q+9�V>���L�S�m"G��D�7�[Gc���C����2����}�S(�V�Xm��R>�?,lwʢ��2��̀���o@	i S��R:��������gY��h��6
E��;��S*��ϐ���?2%Y]�e��@޺�%t�5���&���w��rc��:����v�{䡩2w������B������vu|�lmݷ �R"�����d_��-l���E�W��InX,��6�E�Z��mY�3U�ީ�(���'��U������o�]Tx���y���9.�Q_e/k�������`���n&B��G'a]w�^����g��#�6(���]8�� �(�W��J�z9y�]�Hh�9e����Zh��P��@kc�g�	yq<����6����Yu�Ċ�}�a.����'�����������ƬҁU�K��~�(�g ��8M*�k��j	"�A��Lڠ�����P�.��>@�U��(�H1�{����+�D���)�U�?*u�F�+>	���{�p=�97�d�s������"ko5�;�N��Jr��̇n��S���1���Ӏ���J�l.D"IdgI�3���ǀ����G��81��a���j��6�m������`�N�a�Z\�����V�d���;�r6/)YZ�J�<�;�� 9=g~���0��%p���i��v��V{���i�H�ޤ�~O��D��C� Uu��fΊ��UC��WU�zO>C��gC�>bz2�&���\�K��x�Db �C�9:��t��	�,�}��(X��g�� �s�-~$x�� {�*�����o6'�Z:�J��&�
:�-��N�"8��G��w�@�Uљ�:��_8'�q��ޣ��	.�*�Ԓo��3��}�yۑhz���5�S�ؼЬ愄�����J����>���g��ЫZ�;�2���B�]e;�x��0
W
t�:s'�}��7>cUۄ���=�|V�� ����a��������)-r�g/����a��j� �9�:���b�˳h{U�P�N�����v�{�0P����[�N�k1�jC�A�nq�S���f���u"�6{.t��ڗ�<S���%���.�е�G
�"H"�ղ��F�V�&;�2{TʪP�E��݇�� �`�0�X��)�J�����}/;]�X�C��!�V�&# ����[h	�7�{��j�JDN@g�d��-tB>a����%$]dC�h 6�A�;@2	�l� ?�S���-���yѝ
]�B����o�������?��|��J�����?�ʀ� s���x4�
Zܠ'B[��/�;��������B�������=tO��K(�]��KI]�GL,%���_lt[Z�����#�b�� ��4�&�����r�<v9?	y��IB����8O���[v����%����U�|@��9����Չ��	�;�,
��g�*�R�i� Q]N��S��>XF�΃��7�%����5k�{'���Ko��pD8�?{��z�j*�J��h�:Vn��;(V�\�k �B�}w����,=#��2:�v���g+��P�-�N���g6��e���g�t�L�LwE�V���5(i�*���^j�T_̟J���o�z���]A���e����D�*<��S�n��:����<?��9]���C�0KA��D|����v���}=J$��l_7mM�P���>I_�4�	6Q�nw$����B~|#�@�%ҠH���񟪈k�>)����Ks����U��-�ST��E���u��:�د1��������� ��o�2���'���/���e��c" �?�R�U;P`B?ku��!���e�yҼ֗��\��"[:�_���b�Da?	v��F�N�3cSgx�
9q��S���'eל���e�Ξ�t@��1����ό��D��R.~�QX��$�Ot�	���m�kR�w�?�`������`Ϝ��4�P�3ޜ=݈/����j�&\�#��"4�]�ĩm	�M�d���Bm�✡r�V�o-��L�q֒3�$Q~�h5+$H;D�i�m���h�7jU/��[	38��N���٦.�����B�!y���>أ������d��*����������/����V����pˬ����iZ��\�`�<V�8���o�1��HP��0�
���uJ�hƨiE�c�ٞ^9Ԋ��k2��z��br��������0�YYS`�r�:T�� v�>�>�����<��RV�:�G{��_M-�H ��4��CL*�?A�V��t0H��l��L��-�F$�l�]����XثQ��9{E���w�t���c�$��|=#�t'q)��g�G>���&��Lc���i���o5�����3ށqO���x�r��I*S��n&�f˪)����`�L8�~�=�j�j �R�Sh9�\�қ1������-Ta��T9^��NxdN�{?���zcC8[L�ue���ߺ������x�^�E8�}j%h(^#���:�>���!R�|R�Í���l�Iޝ��*/ӄk���]�& �`J)�F)��&���5�!՘D����蝰T�	��5!X�v^��^y���1[7��*�@<��O��®I'ƋF��Ě{���%]��/�F����vQַ�j�>���]?���k��&�Q�j��֪y*r�?�2�m�ƘﶣL�Һ��Eg%�Ķ��/У�'T 8�ٸ��u.z�Ճ�l�IF=T��_#�|U���޽�g�?V��J��7��W���;�6�Kr����=�LW{�̋�"�W�mi*����\.��
G��5n=k��,-���7:��=���MO7=��z9�
��bK��]��9aC��(L9���1��a�*	Ȭ:��~1�9K/+�DFW:�ݣFs����X_U�$-BW��H��ˆt�A��F&͡�"�g}Y���(�K�[I����ؒ?t5�z���9^���?��b�V�	A �l�Hr�gԩ�v��=_�fV9$°�y�%�*=�U�����q�;��E����F�\[���Aw����:�-{����I���v'>����g�,F��r��H M����7�օ�܉� \Oa�Y�W�م�},�4�EFo
�����������[���r\i���r#K0=ã�2��`^K�N�ь{斥��y��d��Y���y$�,�+In\Lk��N���_$Yz��n~iՉ*�PXƽ ыo1�|�!�ޑ6�+ξ�#fp]���}zm�6�=} �J>;���&e�Ui����$��Ƭ,&�7'��>Jv��	���S#�$d� ?m����><}$�s�B�{e?1ĲU3�s3=w:�l�s�'��0Ā��|MM�� 6q�5�d���&����G
�V3{n���3�t /$�Yâo�}�5L*丹1[��Wpj�s��F�Iw3'_ ���K�O�pSL��aG�\�
�������<�.�x�ۀU�����
"? �(6C�D��1�;�W�;�v��,m��0�Y���d�Y�ՠS��S&�P�ol�����J5��M�0�j<�Hg�A��Y��a�m�.BP ��Kɍ�F�E,�aVLZ��V�JI
~e���MS�H.��#Qb~�t�FR�w��p�	���c$���*B���&��껪�)�F�d����7-tQ��,Ȥ�e�7��;��0�B�իLc-ߋ-��W�8��ހ�(XD�`���`8�hB��I�~�`�b}��"x��$�݉B���)z�Pҽ�������W:����gW��={o�}�����-���.����4dStö'z��߃�����7�
<)!V�a�I_��d:��$-B�&}�i;���������L�}+�OTN��n�xZ���s��7�%/�S��V���7�߭��=R��̖@E�I����*�Ȼ�8k�U�z �����_d��a�
���?OlV8��F��4�w�8��@S�\�@(���;[�lk�nC�	�F��䌹���&����J~��z4���)�,�H���_NΜ.���A��o1�#2�����KEZ�g.3U=h�Ŋ�����a�,���B[݈T�9]\�]W9���Y����Ǜ0�^�ҕxp�ۓ�>2p��x�e��C���!��u�>�]��z�2����vds�l,�F2ߛ%3;C`�F�wL2��h�8��7�mHz�-/��lR���>8[�K��f(kh���n�t�F�������G_���!���8�������z"X�D�h��U_i���#y/m u�uT-g���ݚ��}&D	(����sc�?�:Zr4��6�],�=�~	�d�I�r�*� ��4�%H���:��x�]ITl�uwS�`6c4���7Ē���.��bg��-���b�R/
���K���-&?����ѺB
jEb"}E)��������Sv|���������{��x/��`϶TJ��6�a�glm��"�9�uoJr�9�:���V�45�m T�ҧ>���Ns�Cμ3�.�[�ߙu=��ͭ�|,l�#��+@����L��Nπ�R��I������-2�	֖"�>���9Q�W���"������]�2O�i�;�,s����ۓ��#s-�g���r+&f�n�[�g?���7Om�r���q�Φ���	4�}��l����u�	z?v��J��u1Y�7?\�������8���Έ4<H�K�Ǌ��{��vDȉ��?�����'~� ��%~�D�wX��{���	�E\�w��k�0�a�ڪ\�~Ш�Qw�p{Ǻ�dM���1Qb�%5H��"p�MA�%R�k�ʕ(�4��g ��5�궁IͿ]�0�}!�l��
ҙdƓL:�-B3�-&�'=�e��J<��(�[��8ǥ�=���,�v�:t���(�=�.$oI� �|�N��N��3�4��7U�HBh��zc���z_�[o��G���Sf7��QF�:j��G���}����į�C�}������m~���n9��'G*z�*��u��c�t��x$X���\R��;�Jtc��6'�n�����9�Xi~G�^_WD쯑$�ԉ�(�E�説'X�N�C\�w1� �1fZ�O��В5Ţ�������k�}P�1ֱ�*�ģ3�UTy���e����·�*���q�bڟ ��QҤ&x~c��߿<-����S�~U�)q`��c`�3�f�H�"�ʚ.�3<�z/�彀��!�15��6�[�K���R�#|�s�8꜕�>��C��^�$�b��joyBR� �>�z��w�;"��2H&���i�^��\1)^f?9!�eWr�u��K�2�����u��h�:��6���T7x�@t'Toe3W[��]}�`�����v5HNu}�d�`��R,_�K���V�7˞.C Y�l�-mj��F�*"^�g	n��5|�QX명c�5@�MlZ��5'��	.���R�7v��:i��$���Q)g���m�e�:DƳ���#��wx���w|�#�G����5��L�3�ޙQ)]1��ՖZ\�@K�2�I6� ����oG�W��oxV�MYg�z�4������d"o�ջv���육:�-���匏��C[٬Xj@nu�!|�+��o��)w��E���*@��J�ѽ�� �L�/*)��?�& �a�ݽZt�,XL}�8γ�m$�����G����.K�6��w����b��{�F�3�.u)M	��jt�e	���[�8`n�6�A��s��h�1P�9��ŌB.b]�B�Ȁ���;������Uf�Ș�Rylܳ�T�(�3
Tl����{z�Y�&�m�'c݇H�<G��>�|�u~�X���&/Eg]����T0	�Vw«!�yh�����'�cEĎ�Q�/���Ԡ,���E���~�-��8��{	�_��`fb�R}b��W�a��8\�%v�w��wU_YоE��gPnܔ�{��\B��Ds�%�F�[���ˊ^���a����O���}�7�ULn'�U �ӌϗ�?j�zyd��)∛��lk�[Ou�+���E��=���ԑ$��h�T��;��lYt�C:(���,�f�?�� �����}?b�(a�1m��)lT�Xf��5VP>�j�t	��5S� ������H׬b�Y���,�����@lN��tkBI��3Lh`��2��/az�I%v�xz,w�Q�\!s^�`5��ʏ�{U�R��%3�Ԑ����_5���'ۥ����P�{}�j���{>�N��q�N��-\i�Âo��5l�aQ����U8�9�����:k]j��E$����~T���%ᣍ?N��X�泜f�@fQ���&��mF�c4j�i���ig��yw�;�NiC�ᒈ %�Y(���mJ"{�m�~M?{��/�u0�Kӓ����V�Dc��|���U����}lv�%K a��'��ZA�-d�h�ݾ����?�&xQ�֨ߖ��ݚ��l��ZO���Q�0����a��sNߓ0���p�.�����.d����'��z7�ۀ�JD�<v'���J(���"����D��$gS�g{nI�.`�p���5E��m�^��*�����A$�n���㌠T����jI0|�^-͉;W�;��\K(Ơײu<� �7Rj�� 6�ӱC��Lq�AVe��IQ���mXt;GBZ�]q1���\��/)�kk��t�Fެ�/҆9ƕU�Tc�f��m�)V���(�jO��Y����j�~�'�>@����:-�hU (�G���4b��s뮀]��^-m�𿏊=r���c��Uզ��ǁ%�����d�!�
zo�"jk˔zW����T�&S��rՀ��X8���[�p>Al�������hƠ�ι�����v,������<G��������|����v�tM&��]O�O�c^H��_՜<�/��P�v�Q��b�+�*Vݑ&�cD�r�	~��B:�Q_��w?�c�7n+yڠ�:�v���d�ΐK��O��\�ykNRS�
�[[���!�x���ʂ^������H��u���7&�CU�㘏�ʕ�E�n�Q��ƨA���9��c�>��hHg�����+]��L#A(�Nd�
����O&��<TDt2mq������杞�������7+Υ*���:8�M�d`�2�Lǿ1&u�7!�PZ2��OP=Z^�m�k�![یw���(Q����~�"2�EK�9O)�2a��}�Ϸug< y��P�
�x�yޑ7xn�%
N/���
/����WP \��E��J8��[�l����j�y�9�Ѕxg͵-*���;U��0�|)�K� ~oH"�	���s�����B�V,��)�S������g8GČ�[	Q#�jW��Dٹ�P�TɜAȾd�s�۾Sʩ��'�O���5�&#O�)7-�
z��V�?P��i�]5�ԧr�K����ǒ����*�p��G�;H}X�$6s���>� ���A�(;�̏Zzz��v�2���I$���Cڣ���u��&]��KQ��ʼ��PXn� �i����\h�K7N�#
��]*~0�&�ݣ9�bܢ7���}x�%)0��)&�|a���pT��^��
GY��.O�D*w8j1AS0�k�X���,�ڢ ��wRs�3H�V%� ��a^��Z�}.�܍k.bʕ��b�q�^�㙯}/Z8,���*?�����!��(�xTF��]HG|���+� �D�U�h���
m���w��=��nbv�8�C����QI~�`��|P�땃��(X����^�h��Έ׫{��V�T(u<���ۘƨ���M�����2�8�����e�pD��� =�6b>��S<��x[�K�ek��$�-bA�S�7z5${����������-�;֝/����j�ζ�7����o��vy��+4T���s��UCx�����Q��_���R�)`mJ.H�Rx��� >f-�Ԝ��-Ԯrf�,���� ]	l��e��^h�� �$��K|����	�bEWx2��Q�����J:�>w&=C?�,��v���b�L'/� �Ni��`��/�`2ZK��`!����ڗ�Qٞ��޿]��oEV���b>A@��Bj��������a�X��4�4$䑚!�y���eok��z��o�܅����UC�z|�����_�} �Pz%n$�J������n	�+��[l�Qƕ���"7�A�s����i��imQ��8i�_g*� ��n�yB�,��M�!��l��8�xd#"Pnf_�*���D���$`�n��+Wd�ח�GMM �\ٿN~�z����4�q@�L[�G3Rx�z����!�U�����S�saB��*��i̦�U��$��զ�{	�~�Bo�
ex�l׹{T��͘�ŧ�p�ء��mg &*U���J�� �Lxa����ĿgҀ'��ހ`�m?�V��/��@�f��,;�Jѹ�Rx����nȍ��䇡Ҕ9�.Um�����s��D_ضb�ӳ�yR'���T�|�b�G<>���'!8p�:p��_\Z�%gN���77�G�꪿��Q��b=U���*���?�_�eʬ�u�i��[���Iq�W�?G�r�;�O3����@�e<��|9��p/
Q�l�����i�H�=�l~���:sٗx�J����0s�������U����gXc֜PV�x�����Wb%���!�Dc��b�c��ʛ���4.k��:��#Z��Z�l�.f�tS���/�ubSБ���^Gw�ye\����F�
^�1w���|2ɺ@�*�]��S��~��~m��H;'-���ʛ�{������S�8.���
�ly�$�1��UOW�b��D!>�7����U�dn@o��vsƦ�|�d�<RV�+LI�@��!�K��\�jJ%Y����9hJ��[t�kQ�x��F@%"���k�W�#���_ x���W~6��y��,G�w���M��~��>��� $]����y���D����[)��#H�#��}���v	��
�I	�b1I�T�K:,�-k�S.Al1���,t��ö�8�����S�����?c��(�\�v��*�d�@�FBs# �y'�딶=)�7_�F�K�H����S �!�CJ��
i�#�-x�>~X��̨`~�+�p�ԛ=����~��H���2ť٬��(uN제�9��6� �8R2_�"Q�O�ǧF4F����C�M�3�,-.�Q�f7�E�@�g�Fs	rf��}��ʋ���%q�۟���9w�L�Fཌ��F�O��M/��5�BB�b{ ?�ҥ/��,�a����7�{p~ǋH'$g�c�0��d ~v6q X�С�|fbRo~K��$��܍�C�T¤u����x�̢�@��c��U��8n�jPYL'����~���w�M���H©��O�qyxBL]"'",�CV,��)�Z��G�o�T 0�P!�rw��gݴ$�h��~H��	���3 -����j"�Y�DjSw(��<�v׍js�P Ct�[Z�g���;��ڪ��'N��oeLq�0�MM�A`�\b�B,��}���E=U�a����UV"���>�i}���U����
�n0&-[	*L��	�m�i6�M�[F��&"uk%x�F>�j<i|o+�{�a�%{��?Ύn�$��B�d����%`�B)�V�P��g�=a4�(�%�:�Y|�����͝ጻ���j��V!�gq�t!�L��5��Ƨ>�G��o��1z]�@|!��3�S��i2�#g��)L�����
��c���l cV'��'��7%QҌh{�k�Еԗ��i�Θ��x�@Y�f͈��WL�R���\�	�]#DeG�[|P���f��/L��O��x��;����(�<9fS��a��N*lw"����ѯ���K�Cͳ߸�NU6�����i���5���M�a�n� *j�/vq.�L�����P��UO'���$	�B_J��2g��AϒV�9+k�3��`{i������ ������XW�T,W�b=e���(U?x��$47o_CM��\Iz��G��]�Hst-*�94E�$~�*;x�A�U��h4&(��o���z�;8��$����ٕ��WG�͘<Y��P(*��}�s1�9Lz�G�����E������gR$�(�=�;-������Y]�n�RL���d#?3BS�=H�>�C�y�ݧn8wL@F�頷aJ�Og���*�EY�2e9q�"�S�l5�=��u�����0�ٷU�^?C�\��O�S�&V��%��䘯�ܸ������N��C�@^>oQ�-	�������e.&J޿-������<]�,x�q�x�m߂`ǜ�S�B�M��u��x�t�Q֒(Dz��o�����զs$4��TOB��@����eԡ�P���1t����O`�����S#Jq��6����e%�o�R����އ�#T�L0��H��wYG�'���0�I�L/YEG�Xd��m .�[v��֭o�^f�S���i�7�cM��RO� �������_�|g<���l�vPm5ƻ!��U�A!�DO(D\��#�mM}�>A�n�B�2��WW
Z�t�{�  =3[�O��*������w�Z	雫vy�̏�05���;������[K>81�n-)���!�7��d��Yb������t�> �Y��k���J�@}��l@���3/���H	�� ��8?XH�u�-h:~c���$�ybC[�q�4�C))�v�vk��G;
��e�(&�zk���z���ז�"y=�ǘ��Z�_ Ai��hv@��wE���d��l�:JX��`�T�D�s�p����R�r�I4�o�
P�/fN6�V��q�܅H��@H����)��6I&��J�$�Y�4+4�Ȝ*5�?z$Hv(F�S�z��M'}\�~ȗ�-�HuV�liG������Fvͫ�uk��8v/C�(��g�x�D�Idd��R��y��+9�\�\�@|���ύST������U���$Qj� 	�:l�M���ë�U
_$����w����J��!fv&
MG:������_���ɮf�x�g�d�V�hj���y!}V�l��	�^��A_��T�H�w%���R½�54��Y���cNu�c����a�o�iʤP��؆<�xP��L���8C���
3�|t'�xr}i鮓��+�JWz�B��h�,���:Gj���Q ��9���#�
Ғ��[���E�+�i��{Z���j�QnkQ	/�X�ni�l�<��_�_��_e�T�=<R����g�iyr�A<u4��ug�	��E��B�	�Q���6ҿ��쳋�B�V����DDN��O�vc�i�­�w��?��we��K�g��1�<:x�p���J�7d�����Dp�6]1�tԦ�`�2���_�j�ʣ	�":8!c���=�֕K�z���i���k@�a��/��$jX�F��ΐ�7��1Z��Vމ%��v�s� ,��w9��%$̿�.F��]N=����N�3�q"�\^�7TS�rC
L��T�@]�y���3�^�+�ydQm�xr����eBC���2��q�k�� *��
G��q|#��戰~p[�.����ݴ�}kn!�^��i��kKu���n�oj�Iw���"⳵�84�~�]�H��D��pE�<C|����צFim�y�zF���md7`�	�Y:D�{����/p@
(���x8BZ�~���S�Vˋ�4/�7���c��9�Ӏ�A���4�h�I��?�3c�-�Զ��s�ʴ�m��x���{�C�Y��ǁ�G��V�pi���}*{�1N��%������>�1rG��Rk���[�rx`���.�A%�O��:����,0���0mf5@]��1�fۅ;��G"�aN��g��������J��빋Gb�~�VgQQ��H�E��ow�ؙj;���ji�MK��q||��k.�� �b��.5���A��:Í��R7����+hu���Cs$K����*�ݑ���+
<�|׃�p�}��@>ƾ��|�l3��������I?�f�iU:w�GNN��"	2 Ԗ��FGQ��y��� .�L��F�<!�(�@�����=/5~�O�~<1YQ �!�ĉQ��V(<Iw)B��#��2�����"�yXG¨����ܒ�<����ug������~c�ʈϕV/_*�*��jS�R|+���$۷Lg�ݎ)*���n�̝:ToU1�i��3"�����1����4G����@�[1�x�CQ���M��7	i)24�^v����Y)�>�;+� ����t��kÿ;i�}���YP�C�S� �� - K��ͩm��_�1+�3�,V�":��]T}�n1�5�/f/�l����|5x�O��H1-�����qH��:�3��Y�_����@�������ۺgAH]�,Y�̑� �@ܔ�*���9�`���j`P'��"�+�d=��/��+L�DI,�ٞT��$^ˆs+KW��:���.��QH)4�t���|"��*0��7�y�7&L�*b�Z]_�	��vjd�
6t�Ĵϓf��M͓�N~տ��Y��l��ܽYa�3H7�G�<#���`����8nP�'��Re���`W��& Rf���<M@��V202���^ca%�{P�ɴ�uk
�[��)}��׭Iª\���A@r�*q��٭��	22��5����Ol7 �7���4m/��ju&��x�7��3P��a%I�Z�4���Y��$���31����%5V��?bu��ϫP�-���M�CL�${kU���/4���h������IM��^�=@��R�@���_!���2~��H���q��{G$�*z�m�[є��G5*b�Ιg�&d�z	�&��{��j��ޚ���ɇ7�?�[���;��c��/Xy+wz��uuC��hS�����ϥ� �32���?|���D�8&\�$Z����`���$�*2�}�$���Q{�Vv.�N��p��۟ _K���ܰ[��Sh!1�s	��aP�l��.�IYs��Q�;��nVL�"BK�ue�1R���S��\�����@ZhHb��az����Bp*�7�<Z-@�����˸{��h��OO���Z̡�8B0��񥯾�p�pk� s�80���C��$e?_���6��ޓS�ޒ�_:7Q7?IiW��'l.��{��mi�0lA��+bJΞ�sVvE���Ū4�g OA��ʀ�����k�+9r$��Խ+50Ə�钔�O�!����;��<���Ͻ2��Z�g[1XTI�@�M<Y���EhMь�B9UY�4���T�����l3h���������j�	j�Md�F�D{_e'��K�"����s	9�#��!,;fTO)�N���Ϡ�	XՓˋ�\怲�7RSO�p=�	at,�N�.�[K�M5�d��-�̮�Q����)���əE|�&w��˿kJ&T{��5�}��-��\-�NZE*�\u9�U7���Z�ǜ��G��&N���ٕJ�?e�2�^��Yu�)�؃Ys�?!It�e�Z����]%�K��$k������g��T���l���%tJ�!k.�?ի�8*����_�A���	֔���&��H\���A���sI�H�={��:9��ȁ�f�H �on�E �ߓ�:zG�o-H���=ͽ���������*���f�0nd'D�:�X����X-���O���0���YPPp���M%�~�Jie��Ǖe������S���G�*��RJ2�v Mu:���Q"j�`5L��o���/EENv��.���sڡI[,�VV?%2�XCvo|0��	�[�jF��׊5�����񢺴Z7���78[�6K��"���~1����}�+�1�2����C��/����(�.���{����������P�}1 ��hQ=:�1]K�Ά:_��"#|�8i���[v�Ŕ:�f��u�ȕ5&W�d
�]*�ȨE������8$lKR�(2��FL��A�߯)Q�����.Ǚ�ǭ�K�cZ$е��_^r��G�N���C��',��U��{��I�K���sMH�%Qih�BH@$�����
I��Ni���5�`�ʀ��3d�W���Z��P\*�"�Nf~X����1��I�����{y���^v]c��JF����c:ڇ5�n�Ud��I{������"�a�_���jر�0|�އEm�cĜ�G�6����/�f�2kpz�GnR/�Q$6���T��x�������h�"�#d�|D"��N�`Sv	�ScvG��ӯy#<b&�� 6�6�ʳ�^���\V@ysc|zbu+�J���+B"� 0��A���g!��d>se�.��ڡ�p�20��G����_����ܸ�"�`�:H�n�]�S���L�T��\��|1Q���I�M��t��z8�"6ea��P�|3��h}�9������p�7B���FK�(�|�(�qU��B��!�r���>x���A���zKu�M�+�G�I��`�٠�|�;�
�ai���ˉ��J
^�*dgZ���x���'�}QR5s���zf��u+~!�N�{yF$��g8z�%T��-��?Σ3u�UXyTN%���q�a�s��]�*�Q�p��`?E�;�uu�x��N�t�`?�z�t�Þ�v�
Eyh�Hd�-66Í�z���Bҩ1�b�X�I�c�_F���|�m� ��o�1\m�1����}��j��-h}kO�<�ct��"�-�m#9�GP����|�����\�9��ZM���z�^���2�F�Zf�l��ȍ�3�bXw��t��Oc�ʘ�y���&r�,�w�G����ي���I��Xvv7��*.�$�NA��n��?��Bh��T��ڴ����0��"uc�c���X��ٵ�,[?�E}5�5� ��[�zq��.`h����B�cϤ8s��\ѥ?�g�O�=o��<�\\�\E�:�g�����{�]H�̡�_(�^��b�IP�n~�5��,Y��?��Hl)�m�j�2���.�Q��=���'�\�D��K��_�]�r�m�6���f��Rg��Y�Ƃ$�E��x8�82���'�$"���5't��h��o��ȿ3��<D8��۵�4d�#�a����67�?l�8J�����4��A����h	Gꆓe��+;���Sy'�-	�����F�t��'KӲ�$��f)/���W���8��ɞJ��B����e��U&�������=|��I�]��9a-I�z�~Zn��v�=�m���P�b��q�4�K�؉�p�Mx��S7�s&��cd����S��Q���wB�]�_��)(���:?��9��l���ms�B�^L�SQ��`����oe=bho�}s�T.��om�ƶ�p9Y���pb�'�x`A�s��Ky@�;�6B��� 1Y/ ��w���" $m_���mY��p�^��_���3�w��3�d��X��~֍���w%�K�H;��Y������Í�l���0<Z\���qOdH���׌���֠=-�Y��k������e��v�07;�yo8FtcdL�_B��Ǎ��(�a�����mኴ �t�m�����(�4If,��S��0��j7Ah�{����w%vA�m�����v��h��8X1ڗ�Rh� � �X�_�Y��R��ѳd2v��lX��/�;�f#�\tTmܦ|yEmYBY��`�¸x!��Bk��Ϲ5u��-C@6⒣��(�
~"��ե����H4�~P�6��쌕�C�:�jf�K_�U��y��Lz��H{1qe�(��]�Sd�6*Dt<�ܼ��ĵ�j������(�;��* ��<�b��ߚ�l�G�<�! ��kxݾV{7Z�8����LB=�-<���r�+oγ ^�[��t�$ʂޑ�ȖW`�3-h?e��c�#��&�����Z�.�P��{100�e��3��o��m����Z\a��.��c�^�UB�w�����+Z_7��'1�A�s�<a`�g�1M2���@���R'����U�8�Z�|8����?����˳�_Ïx��7fl�^x9�Iފ��C�z��h�(=��Ź0C�㺶�	�[��<��˖'������m|n��k�+HV�E{�w�x�c��P����Xbf��3ظ]�}k
H�\/�.���2���� ��F>t�N���rJU*�)�ݲ�l��.V����9��RR���M���4t���M�1-���O�T�y�k��P��&�����1꒕�{B����~�5���5��o	�Aw^s���d�Y{��2�-��G�5۲t�?ߘ5�˵�]FB��ih90�x�q 42u&�DO����߽v�]<C;݈=��ȁ����
��8ɣ��=�S�;�i�z#���|�f�e��(o��U1�"�'�Iq�qΝ��&tT�8�E`��QoSyS��qs���ߐD�U&�\h�=���̖��-�Nmx��w���U9�*Ō���-Da.�I�iQ�ҹb�]��>�������y8L[T~َ�s� .a[�+�n��!�܋i�(����y��^��ݷ1��Л�@Etx?�m!�J۴���g� K�S�W"�p�`֟�"�H2fu��ۓ2��G2y��W*������ly�-ӳ�9�\<�%��{��0�n���� ����i���Ci�I:��x\f|��5�L�cW�XGYL#|��1P��vr�A&�[�8�ԋ��U�S k�l���2�Ĕ��=b����ßU���Ŝ0}�\ХGlD�	�M���3�=��;PZ���&!��+�}��E�O�Yzp/���Os���*wHw �?���k�$���C��OM�ł�q�"C��S�T�N
�LU��E������|fك���ϖVZT�X�Fe���ҾK�*��LL�3�̨��I,�,�Y�-;*���	7yM�CY�����ȽX%�M���/�pW�f�`cmB��A!�3�L�X��s����ZJ�I����Hat%r'5�i��+�h bX��J[����a�[��ut6��C<ۼ��|�Za��߂�y�M��������| ��,�4JL�Uw�>Pc����i���]Ȏ`Iη'6+o�_�0$:�@Ij��r���J���⹨]}���,��O��'2�S����C��a|�SJ�� �XD�qeT�%�h�	B�0��m�/��4	��~��L,����i�v��_�ZtRc�Jʾ˶��M�`��@���	Z? ���h�꣤��%�g:˺C��K=����c!�����g��<fp��V�Q����6���8��xP� �-�M�t���P-]�&\��G����0x["ʪ�h��z-���F$�{�=�`a��#e��Ik�?���6�:ׂ̍��)�|���[(p)
�_��ʔћx,S�&�tv�{�H�4�
�\�_Y\���*�c�֌P��C|XK�
�3��,%8��J�å��,�K~'F*=k���IPL<<��e��w��ǹ�'��]�&�ʍ <5n�]��Յf�,�QK��	dC�w�mؤ<=�}�gS/\;�z��:���D̐4�l�4���z�TYY�D�M�)s�:B��ع��1l �B���0�:%�X�E⛚�Ŋ�A|�?<HT>ѹO($��r;P�>��G�L9����E˨\��WW:߄�����#Z��}�5w;)_jH�&��E?U�5�[��5�/:&CtK͒z��llԋ�)�z�*s�_��G�w*�0O`�AB{��Ι.��|�3����Q{a�s��F>o�����pI�[H�
$�l�Y�S1���[0Ͼ�.о�{��#�;s�@Z7���*!�a9�`�U�jҗ7Z2�����$E����h���f��tx>��6GY��¾v�æ�������a�;�`�CI"P �1�,f��[�o�E<={�[{1Y�Gy�9n��L�yJmx!iPәn�8��UQ�UyP�o��J�Z�����aH6e�:����t��6>��Pw/��#�[gk�a�a��$��^`Ŧ�*���Wmv&��m������d,߫����Z��ݚ%��;.����� ����+E��Fn�s�3.�eDO��yH����1���_��36�� 0�̱5�H�7�f;���%SUZC�) ��/��>�a9bzn:���UL�=[|Iw���vF�(�vK��v�
�Nk�A%��A/��c����u�˶���4���d��؈�Ԙ�'�ҍqw1��H[�տ�g�B�F�#���D�f���5�#P-P[iĭ��<��o�׫`�^>˻ħ�)����!;�ή�o����{g�7��_
�����57��%�b&�wy���{�Z�>`��*���7�"1��r��e����2�1՞����s�Or�vw��(K�[�Q��;ؔ	=1op�@��DH��fbLkU�dQ%* E�:��۵���p`�nCTBw�|w��lɯE d@wm�)��t�S����=>'�g~������Rz���Z^�J�ұ|�X�=ʻ�x����~����@601n�N�,�~�af��fa�p68�&��fx��fT�����ɦT��^�/��MyV����I���W�Dλí���B]�^F�	3'1��J gQ�������-[��$�_u�Y�h-�U�-�g��)�
�ѓ*[qnPe�y(��S����5�T�5�`�kG	?A��_D ����(��c�E��'Cz����Cz���D�m�Q���j��ߐ��k�v�i�A��v�⢾]t��,C�oE��	pku��,pP�^�����<�Gh�8��w��i>{<���qĀ��%Ł�k�)-�U�6��� ���Hlso!EWS���N4x,w?6���c��r��xk:J)ejAH{�����λ�ם3����h���x��KC����Z�!V��VO̕�ߢ�\JoX�J����4u��|/�A�G#hQ����|-�D�ׅ��⪃�A]�(�!�2d�
��T��^\$:_3�����}������HN�����.Gn(C�]�,��gbi�͚�]��L?��0�k�"5d��wo8u5�!^�F�$�2x��j��yp,����G}�O���^�4r/�ER�F�:�ӭ� F��-#5���'}VG�+�VQV-l�ŵ�Ui}L��[��j*�S�ރ
r�/=s�R�VZYR!�0.�w�2,X��o�CL�U%�rWxb�)>"YBb	~0�J�{�E<;���i8�<��x�QS��s
����ɪ��<��Е��GR��Ϥ�=gA0�?)�X��p�u�,��A�2�R���	��C�z_��E�Ԙ��Bժ���I�h�$T�]L�ክh������?�t����y��^��;p�|ıP���_�Gr&�a��
�F`0YOl9|=�.�3g�b�!s�3�*�%���^��baƤ.��eW��T�z�#��q@7�q^h;�c;��<�'��U���7LI�����w�ֈ#\*S��N���T�d�'��;�P^v���/�F�&]�磿������D���Q��s휓J�9�����v���I���w�p8�X�g�|��(cߗ׸��#��z"�'��(�ȭJo�ۇ˄4�#��Μ�O�)�S��1��$���ق���ⶆ�q�_U����߮*�⶛4� �N�B�S33Z�#|�o��5'�~n)�� ��+U���'k���Q�E6\8��\dݭ�"�-����#�T\�����66:���?խO��nB}�0&GpO�#����p�V�}�Q=>˂��Cp8��������6Uv%��T��mB�;oh��?-�USKm�����YDʣѾS�eva����0�T�]�tochi&�BD2���"t�Y�w��4*�x�]�)�#����[^�(��`m�+��v9�)8�0H�`������� ���R�<9���K=G�m�`{b6h��e+(`���ĥ�^+��dR+e����;I�z7Zd�U� ���_��GآwT0����8��6�%L�iR+�s�G����8��Ԡ��+���
C����m���\+uj����'	4R�E�rN7�h����E��"�g���ZS�~�D�������z�s,t�.�eN�E����e���?�k~8��>v�L�kMH�hP�7�OWb�p�^�(@�0��9�����R�����`�9�0�p�V֞e��=D"e�·�N����v�j��K�.ɭ:�59��{v�<A�Ƶ��;�x�p19�ӻ��;Z�,?�lb0#}$��M�q�W_ሥ$@�>}�G$�M.U��V�����D��$1�E��^Br	��[�\��;L�Nb|��#�6%-��髻����@*�!g����m�v,f�d���+�+�fx�a̯�ZU�灥;mZg�1>RՐV.|0T��ݺ�y��n�3
'���C�	<X?*���$��l���)o��B��9�'�v\&���n�E����+�D��)�K7�W���L��n��p@��9�.����+=0���i����2?r��c�
%�lMn�C��?��e�d�#,�h�mJ	92� ��Yi ��u@V����E�A�4�h��^H	��9I�*\����?�i��3�s0��ɺCS����/规͓S�3-fq��܎����:R�Ns�+�!`��oJ6L��eY&�&6�!bF4o�����Ѩ�iC��p�\�ҁ�'PW�wH�	�:�'��l�o��҈/r�`G���0d|�� ���;��7Z4���M�R� �:ƿ�� !��r�������B	�}���O����]�	�+ m�(|�����{�po;�"4�R�C�b�^o&:�tݟ�셩��Zҥ%���|
�V^Bb9�w��8u�*����,HX��,Ȝ��eT�?u�*�t����S}�J`e�/��%� &W�����;�-lJd�����v�H�5�Y�[LV~$8��2�R�sb��$����VN���[�G�0�LO&l�W��쭔�-*��0u��`��$����-;w�{�Sp�l��ξR��yL�0��S�tg4� ?�}�x"�	�GɈ{��>���_D�1�v����{G^|�Z2u�+�\�^Ҝ4Ч��)(�)�,a���!��Ą�2#e�.�V5~d���ɳ��+
J�y:<&��f�;��l�ŴT�jC����YO��|�h�rn ��6Kӣ-ŧu�F���j�e�~�q[2�E�7͘��Pq�64��y�|J�"/ϖ�O �[��/��תσ�&x(��@G؋���a�n;��t�Ӌ^\����5u}0�1��s<	�x�1W�j���C��)���<�;���c�ߺ�	Wv��+�5�h^�|C~(Fx��f{N���g�U9�̤�}ŭA�[�����
�9hjk���G��g���]��'����5.O�������cs�ss: ��L�;#�^Y���{���`� ������n��anm���������2w0M�ݹ�C��g �V:�+� �5��|����J�O"üϞ�K��X����a��ݓl'�^��n0��ac����ܘ�z�Jl�v�j�!�Yk^\�pގF���]����B�^��|[@���S{��>>y◐Mث}yO����M�&���N���eK�-Ӧ��ul���FL���h{9�����9�}��yo_[.`nK���ܴH�]+�|�}����D)װ����±��f�C����>I����:�X2t�?^N�>]*{��r�X�{�3:�5tm-*F��m+�u��������z�Κ�^T�i�Ĩ�Ê�d5�l���6��]A^m�%Q>� �ޓ��m�:���Ji?z`'`��u�g��1坫���u� �Yk�ɯ�&�����f�Ogwd�Ԅ��(Ԋ�wy���y�ip]�B4%)�/���\�}��\\�����k��e���ݏ��Y���	TV�L�78��<�ɗ��uP�U���j+���&~���b�R����D�4���2^i1q%�.+�����R*���r4@��q�����~'߈�*0��cE�F7'���e�s�Q;j̠�yӴ���q���OX�^��~�U�$OݪZ�\�^�U �?��FS�љ���O��o� b��ED՝,Q�=Tֈ��V��w�t�_8
-���b��Ia����oy��A�	5�;��%�=g� X>r�+��&L%��!�?u�q��R�7����2v[�!�����Ϩq�����o�;Ċ��ȀT�o��%�_�����L�@G�L����ܥ�:�Eh��i�4��_��W�kx���͏.���H/쫾�;uk03�=�鳮,I���@vW4���r�Y)�r��MF�j���;5!�E�)	�@��!��/9���kd�l뉸�#'K��a=�غ@mL9�J�����`
L�|�u�җ4��4T;��a^���t���A��ˢOj��U��b^l%��[6c��V �� �*i�"��DԷ�٥Bs�R�����%��@�U�#�1*:��Kap��K>M�.҈��٥�d;����jE���V	����5�CD�]f"~��:����b��O��b�P�	�R�Z�*:�����q!�v�Vx�/S<�j`�@
jW�4��?!̅��d�i#���0�ؐ�L��]�9�!�������]�{�Tv^M_��ݻ�U[^a?>�~��j�m͙In���S��'��C�'H�T�R4F���� �|���8�wF���guJ�b9s�sy�&��!�^L�s�f�E�\Q(U��H���a�?�K�7�`�	�)"�������.�]�9�Jk_Q �!�4Jx�5[���cL�F(y�����U��z?o"���ә}9L`D�m/������)5�ՌSh��K��H�U�0>�F��@����Of�����"<�6�y��uG ]�}��g��ٝ��ݿ�k2�ˣ�d7dUےDX��z����D��������n���+�N��1�G{�� #���1�a*�2������� ��[��*��'6+������ر���!P�F��qF&$�vr�{��O������C&�}e6��,CXl��|�,R��mZ�(��#7�������b�V�Ȧ��B]T��,8�m��\���cg��X Tb�)�����=P�Yۛ�8�v,?��z�k*�[r��#�����C^����JlN�Ԫ�ע �����Ė�eE�����x�s��q���3� ǯ��I�1w����:#��͂Rvq�M�'�YY�q�;G��!��(�0��7��J�'	��̹cМ�MM6�dCL�bֻ"��ڪ ���m�/M|�;�Uw�͕{儡�쨐î˼�֧���Cz��{c����$��wzl�/�����IL7�&�/ֆzQ0�^�\vA�T�|����EÂ(�К�f�L��&Fz�qhy��u$�XO�zx�G���b���K+�]�����}s�T�uo�� ='�uJ�׿!�#f�_���_�)�U�m"i4�b�q�5~�G�F8\�h@J@��*m+�A�2m.�3�:?-�Aqe3�J���yzl���3�6&�Q%F������Ї1T� ���N���_�4��q)�8�w����)z��l����q�ǌg`��_Z�\#?�����e:xI'g��v���u�1h'�lr��Ep��~gFZU�%1�L ����ވn:�ƾ�t7�X\m�v뫰�\Ʀ�D1�s�{s�@�ҩmJ���-�z��A��C��۾�<D9�/8\-&�ܦC�w�~|��;SޘC�1�����?[��N�]��EQ���E�De
�Gƚ]�s�9��tӧ�+�(��֜T�AG<�b��~{�1�d/��
��ELn���/WG���F��nڈ�^�4uc�)t��1���~�Ɣ�q��2w 5e�^d޸�61J齂�kp\ޢ��Hy	CĠ��>DKg��k��5�˳RA�`�˓����`�h"f����<��+qN"���U�V��`��V����v��sQ�6=b��o������$���-b
�g����qJa�o�6���K�C�*S����Ȗר�%�SkC0nɼ+�ғf�8�S��Rj��)b!�F\7	�T@�b�y۫jxӢe�\я���m�ʢ?Z�0J?��Ɋ���U�"���2�-�����g���n�k����X^GTR��
�+�J�^j�
dl��d��e$��������r�V�#+?���audJ*���5ݟHLa�[����#
���m��f��Tc�!Y&'���mdb�FY���1�0p5�����N� P�v�t�2ҵr$Ū`nrvu!��u�ݰ�Y��X{�+�*	��>~x�%��ZP�>�F�b�q�U:��i�˄���j *����a	�{�8�Ҩ�m�fz?��@k�9;����D�r�p.�&�CH�~k3�s�ބ&�\Ss�݃�a��wf�(��$�k\�tl��l�۵�(ڄU��m���*
��I����h8=_��֬�O����T�@���wAm㢠D��?j��1�ZH�"�a��a����.���љ���Ĭ[+&��}<�W��0��,s�F��=.}���l��i �m�q�'��Ŗ��D?iĽ�F��"m���'�c&ѹ�HF�߉.�}�0@���P ��j�t��_Q��_���,
���J9T�GK���+SQ���,�k���<�ޚ�O��f�^��J@K��켃�οXQk�@�q{�6jq���u�A|��ߗ��^K��Y�1;e�S`#�{v�H]8;K��� \�a�Aŝ/v�ϳG�Nid�4��me����f1�^T�!�������E�*�����q��̸w{>˘=h���;�`	#�j�$���7-�O ��� ��io�~��x�2�/�1�[�`#����S�l�K��l�-��^��6�#���d�۰x8���{Y�(��0��� �j�用��o��I�O��3�kw>��?~봹+�DX�f|S$i�}=t�↫(=��h��~������q)� ��L�#`iD-}�ּl��-�N���Оė}>�AA�:����^H_7
���{�&�[��rޞ0�#^������/��A���:�]��܉	�r�FX���'�ŏ?�����%�⎒��ZZ�i�Ķ��S�8�5$�/�H?�`(�I�k��eEܫ�DlE�������gR<ǲ����A�]S�m/.�5�������~W�5��
ΊG����a�	���<�Ej&k� ��;�6�~u�.?<d�|4হ/��Xn5��50c�U��Q�h��3����v��B�LU�a�������)������a�ّ\M Y������M��9����Y-�8#z��M8�ta�^�h��m���0^I��o���x�5�?b��]H��W��Ȍ1�6�yJ��ٙ�`{�����4�ݍi
��?4mYi,Ehp��q�nX��\@:���f�[��_���vA�仜|��+
�#Rdۗ�6���μIܱ���"l.C�� ��	�8$��Y3�	�G���y������>S���-3� �b��E14Z��i><����Vd�<t��n��{F�2�U�E��%�ò�Dn�Ҋu�8j27�[ȅ�4� a����#��X��PI�Iz��!�0]���)f�*�,.r�5�VĔ3`�D���v��l�F@ZܥBC���[���YK,��� &�l#"�>8͍sw�:X�*�w�b�D�u�X����XoWV��K�b��5�!L�0�����{��W�q�&en���`�y(�"��`��&���hF<��Ͳ^�I:S��;�� ��Y�`.3K�>���.�4pp��yz�^
,ބP��<�VZv�S���h2������4�$�pJ=��I�1ܺ�ȅi��.w�TU��1�反j�#X��ïNܾ�z@lw�
�y&���x�t珌ee�7�}.����y��7l���k�8<XF�,����%�������T����>5nT:M����eL�u�P�<YV�jq�o��u�Ҁ�_�����d�zD�Б�E��ҋޏ'3�P	=�?Ѭ�חffJ_��4w{�Y̥��a���N���{�]([�d%���+�b@��h\V���	�}�83s�TA
�O:��N�B�]�&pY8}���;p�	q)]�(xG[ZxXI��Fp`�w?��L`���RS��2c��Ҭ+Sc�ÁU屠)�#<��l1V�c��׿k����aa��j��
�G7;��<�ׅ8���/3�j�tu6��X%�y-�tP�S�a��,���N� ���vz�X*Ԗ�w�n�Q�v$)�@~�Wi"=�_V��p��Z���r	�3�D�yƍܿH��ix��v1%|r��IN�Ag�7D�r��_/�s����2�n]T>0�8�ǽ��<������q�Й�W�?b������=�vq���y'���r�M�.:7���	���yz�d	N�n��c�zD�剻�9m?�8KfG{(�4�w���#�<f�u�D3N�����o�\aH��F�K���$퍍��v�h̰{��sV���k����Π�qS��f���X~���^��I�!`�Ģ�;q�yaC�	"��T��#*���U�S[� Ф�~��O��$�DD��1ڲ�V�V��x�u뜏�����P���D7����� �~�L���;�U3��b��ch_b�c��R'w��j��p����⌱���N��h��.��ُ���2oӡ!6��������b~�W&hR�ڋr��i�=�յ�T��i�U�Y��&xȝ�mkICMFv��G�]�l~�1�Y�}�]��W�?�Uh�=b�|�3��gW؀��=.����� ���3�Q�N�y����nХG�'к��D^�ë�;7|���k���q~��G����-Dw���L<���;bh���.�������l�9D�Er�w_�踫=�^�W��r@�t���@jс0���Tq���^����@���
C��%�r��޴븅o:�->�c���!�J7��:�[׶w+W�7�vc�J�
���gXq�{[�=�V+����_��\�v~������'GoB0���/$�p�*D x���KbbN4��a� ��|������@J�U������&�#�q*��cև�Wv������Q���v��b�ǝ�}���g<�����W��7h:�_�@t��M/�TDfQ.3�Oq���	RZu�[��y��K&��㢀�U���ӷ[}G?����
�F���
	I9V�
��?��&��M7��g	�:��o���;�Z� ��dnd���`�Df�E�u��*�G�4+8���T.�?Г���"ٵKG�}�S@�m�M����M��1�$L�4g��b
>	�%J�_4�{pS���3^cO��j�	'_�y�)�Ŭ���Ak!8ٖ�̒�7��d�y��P�y�[��k#��R���J���f'��2� 3cm:�~=x��5��QԜ�[�:��p�͆~�F���Ʈ `� ?ȫ7UU��E�i�:�������[�)�x��7쎻	�����8m���wF��'�� 6Ql��V-�ծP�%{8�J�^ό'��,�kI	y�zW�q{A�Y?��2j�>�A[�<��'��m���}k�q�S�|9at� �n�2�y��	�4�4���_M��6|�*pG�t��~���K�YӒ.;����1Պ6!C����[�6�l����.�kl^���4��e!k"����3�tr��B/�}e����CG�s��t�K�=������ҍ��ϝ2����$��Ո-�Q\���֞�X�?%��=<K}��ͱ�sOֶ<���_���"~ ��0B#�>]�%
�FO��!U�^ͩR���:���O�%�:��f.Yl��w��U�b��a�r���mz�L>�hל���<~��7ԡ���5�dR�����U �m�'���Mȯkғj����H{���qk�\�����j�M�Ui�}n�o��36�wA����ʻ�#a�Z�نnc"�P��԰ m�@}����	:W8�%��Hm���Z����P�R,^��u���f���q �?��:F�B��^xү�~+�gulsڳ^�m��������g��C���y�1�V�������?��:�I�Yj��Kz?��c�8N��(�Ƒ=`���1+Y���8��L�j��q����	$A�Ĺ8�1��a�~�����:��r�Sf��TV��X|'���RH��֡���	��r�<Nƭ%o���)�~Մ��ىKQq98��WW����B�g��>"]#1~ϼ�`�m����(Iv����-(7�o�����o�lJ[�6N:Tao���/��ݓ��Ԋ,� ���	��*�!�6��cV{{��6�K҉`,^ɷ�S�h�6l~Ɋs�;/�x=�J����r �h�G6��=��ߎ��� �����d���c��F�5�z��JX��:}=Ɣ�� ��9^�o����f����M�=S�%q�����z�_��#���4��(�),l�������s�x��;?'�����p&CNfR�N/6pZ}�1|�+P���q+��x�n5�F�ᬬ�>X)y�lj�x��|?y���[o��7��b	͞u��[�#��x�8�������|#�����ݙ�_Iٴ�����L��`;���VY�ornM�P!�)��i:I¯PQ*�h����]z��
V�+����V�`�@�=�s��x9�B���wL��%�8���`^��p��#_J�~0�'
�<�H;��"�y)�d|��7�鄓�E}o. ���Y�:٧�E�v���3t��`(�v��q�.��*є ��ǭD4x~��{۾�<0F�ɔZ:H@G�C�����2C��~.�k`�5�P8��9Owe|���z\�&����>ѧI$�&1OѬ�� h&z�9���y1����[��g�7*!�`v��H����q���|��f!�po�Nk���+���M'DdE�J��[W>��Ҩ7e����sL(a��!k�����V>Q��a��kY�9O�e�ҍi�F�&N��̔�������晑Η���j��@��b`����#��j��lKIKwl�$�}��2�+U^[N��)��6�JC���I<���UsE�M"��lf�؞����g*�ż����L~�e ���(�+^l(�[E�1�<-[%b�� ��Sj��o���G�:.��(`�����].���Q�ZYf\�W2���K+b�ȗ)E�U%ZҎXaR0%%o�O���F�%Q�s��D+
2|6����Ha��f
����c���J�=�Yrm�;��SE��Fv�H�f�,��D���,V@��I�r�(�a�eB�X���H��U��x��E��j�JQf^��Sy$��<�V5�ޞ���J�u�f�ZM̄��V�<�n�ۻ�4L�'gh6h�;��%=�p�o��'Ʌ�ag��ʒG.��Z���3f�<�,��?Vg)vz���Lo�Dľ�œ�?����H���1� ����z������r	&MՂ�I�țH�o���gB�Y���N9��@��l��X�bs3�㫰m�M)R�1r:�I&�/�0��gD������XM��2r�s�\��+���e��ZR���.Lc�nǹ� )����շ'�-�CH��9Or8�nog�9�Բ����LB6����<<_u�i#��i
��Hf
�92��c2R1F��x�41�&7�7�@O�[�w��kE�ɾ��n*w�%z�	Es��Fz��~[;����Q��!|��L����g�u8�� �2�c�0ލ�� ����s<�K�/���T}�j�#(;��~VP�Ri7�qn��xi�����}�]p���b\�ڀ��XP�w`a���h�sv���B��=�R�� F��Y��QA������`^�����E�)�%�d/hz�]
���]h�1��R�d�EZ݄��1��G)�_�c�y�>�!$�Hwb��9���Zl��B�;Z���������؍x5���i@㮄K�/J?���@B1,=׊0�5��h�B|7x��gc�N��|y�h�M$¿������\f��~��K���zCΖo�Xx��΋d�,�D��A����2"���������^7K�Ǆ�fTe��=cO�1��?VaL�����vEm���)�����Js�y�C a7�t
�Iஆv�;�/����1����e��goM>3�M���◕5$s��sf�o|� �5^iR��Wm�=[��D��]�$��aac����Fk#7��`Ϋ}�3�E����/�V�B����2
�1�C�m�Y�wtZQp�WiX)��Z���w��[R�-��2�r�>�"���|�g�tئd+mg��S�Z(@-�k-��/�C�r4��|���\���8�}��C���õ�94c�Rw�'O?�J,���h3!z�Tv�裠�1��5�8��'�x�����v�rg�e>ä�9�uk`c\^c@A�O�Z�W4t� ���������4�ﵷql���ˆ<��|^��
`Q/N#��͊��$Yo�����8Aol�?B��Q�b9�n�X�(��%���cٙ�O��PH?�l�j��E7}�f�P���t� +�rW�*'^�"��k�s��E�{���u#Ŵ�����jB���ϙ�����ks�-v�Bb�Z�V C{�:�W%| �b����Z�u�����@f�����:�����[ k��+���ᬎ8EZ�X/��_f��I�	�!�^[&͇^�B��������z!�;Z��[�f�*�g�MA��e���I�!^�6ީj��Q��'�mv�s}hD~x�mD!c�ۤ�֘�j�蠏��[���
��2�'�J�Ad�:}��iS���CR���I :y����0��5�N`�����i���$���.�5�����8v���ϣS"��܆����rh!�rgF�"���0Lc��r�ӡ\�q�qAP����)��IW�f;���e�<0�s�무���!C3�<��>
[Sɥ�v%�V]< �n�d&�Ĝ ����N�b�t�؋��/T� K�wlÇy?LM�G��`�h�����2A����9��Y���s�0�{���\(�$7mJkϊ}��Wf7T�/�OPه��)��H�k@������-����7$sS$ӃD���ٽ\J���O�l@m�L��wb��Tdh襜0�Ê�b	ش�=���1pܓ�B�XK�q���ش�z���p�X��50�M1��נzUd�[([1�78����(��?r��}{��sѕ�V�ފ�yt�ʎ&摌�I���lt��(߹6�~��ct[m��/ƧkZ9�П6?��#6��Y�;F��+�\q�5s��E�ɻO�S#S�/X(:q����B�sCb񘥾{�y#lS�٪s\��q�T��W�C)�Ke��~t;PhP:r�<(�<�<	k�&ܮ�LĒ�pR��-�'�ǵK��$�9�F��{���f�CF#� @#{���n���/���㨯��a-�!�{�(��U2���ڑ ���
�vp�`&������i%
�9k�fc�P��GYN�	��<g�?��$�n엵�<-���F� ;��$�Ux��V�G�rP�@���=��υ�Ǘ��}zS�L]�s�uF�.?Pb!�2
%H,�>lL7�Ց�	B]C�E|�W�X|9�CO����֋1��&/ڈ���KV�v��ȼ<	�>`I}�+�Pz#�|��0P��2�a�,w2�z�,Y�R27���fF���;��9�z�س#�ÖoQ�Gb�lض'5�PM"���lg�uբ<r���k�����%�}�B* Y:�`��r�b~��X���,�|�%1-���)�2����~�D�y�yO��s�+%��5?�Uu'p?�FKPζS0��u?X����spz�B����;���/iS5�,f��y�G�ʣ\����K��S2T۵^�+h�HI��� XY �.�0����!�L���� ���[�q��-v���b���[]4�)2N�����KIV֨�7��3ֹ0��@�7$@t��	�{��m0i��?�?�Q/�e��/�͈6,��HKzt3���#ŏ��T۴�c��yV.&�`�T�N��μ��ky�Ps�2{�_Ѽ؄� M�]Wdԡ�5�y�r��2�$-L�F)���?U���$�����wNY�[�E�dW^�O ���R��G�^�m�x�z�ǔ�j昆Kp�C9ధXIܷĥ����L=��)�t�H��=��z���Z8nx�s(���w8[��Z����2x>�4ι�`o�6I�O�R����$��6>�`�l�ud/9:hѣ�
��疣�2q���7��ŻQ����z���=C}~��Ն��������	@�V:B��U�R�?p/��C���k6���m-�v�pg!K�-�4s�^�͓�0~�d�M�/5K��T�,S���I#)���c����Q4��oG��6�y�&�ƅ�Łu@8nŏ
k_v1��m�*p/��P�ٹxMљ��^�����n!.�aڡ���?��)Up�eXʧRa�=��SQ�����P)� �D���e�j���z��	u���3���2f��c��/-@J�m��4CQ�VY_�0ʰ�A4v�8&����i�V*���'w��P�����Ǩ�t/��/�7��F�k��D��g%
���+�h���:�akG�����3�����)���J�/`�+��:A�B�T��?�#c���m�]��'��N=}E��b#���K��Ř.{1[MG3ɓ��U't�tz�}9��R�luJ��v��
��A�خ�y7�b2��>�t�c��g�(-O��� P�2Gi�_3z$��� ����˯wB�:�}��p�����9�8�H�IX�u��\@��t	��),�3�s�K�ql8K�E�GZ<I腘�R6�k�En�R�~�S�7�2r1~�ˉ0(Cͽn`$�\���z���٧"6�`��Y�7W�r$UkXܤ\[J����ӊ{1���5�� �O�����˴jw�z��Rr��s,��v<g���i������x���A�?|��4ڏ�wXd�K)k=��,:�m��պ찄G�7~D/tb'%�����Ή�L�q������{F%��9�S������h��]��{y��󬖦Q)��?�jy����z������F�ͦDou��M�����{c�G�֐5�a�`�D����7?ᴨo� ����^NoT��H��(�J˧���mOm�M0/��^A��SK����
�&�	9Z>WHƔ�`x� L��2�ؘ�O	OZ�����#ɢ�xUR���`��ճ����Q�.�Bo=�����8q�!Ø�a�����kTu���K�i�*��+��l:k���!��Xk�FQ+WP.�De�R���J�܄O���7<X�*�^��6��C��}Bu�C�ӽ����%��S���S�������:=���S>�,
 S@�����QX�#��/ƈɳ���-Y�l�*͡:�
L�ثE��UQ����0��HX�]�����n��ӝ㺹���d�b�9ȏ��i�$��$�߾1��Af,hÃƯ8�jxf�'72���)R���Bʃ��\\�A�o�[n���m�"FIS��+�ZD<�P��ɏ�:U�@K��}.U�?��T��g K�"�^�_{��.�TL����T�,��F�ʩ�)TV��S�ϷK����s��\DFmX�̎��4m�1�z���+쟓�=����K�D�$��`ꛃ��<p�S]�-P��c�(4�^��M7���^�l��L}&o�ĭ��]뺫�!W���W��>+j��o��F����8�AڠI�K1��.m��>��Dh3��5� 5&�jZ�m�w��xQ-{)�(����������_\;}Cj�Y�����X���T� *x�*�[�x���H
�n�K��VZs!Q8�.��JH}vzz. ����z���y�`�s���r	�`�@[fK��mw������K2`q������o�m��x	;B����E����Z�{:�iZ@�M��h`Kv�V�J<����H,���d�_�j��ͥ��[x�o�}���Yf��@��(��e�����q�z.��+D9Į�8��L�z��T=�w���}�4�����1q����h_R-���I����:��2�bI/�<���8�(gl,L0	n$���j\��Jᄅ�Y��H����i#j̘r4��B�Gw����GU*QAݜ��0��r�'�Q�2\�g�vx��٬.<���BW_0��7��<l�N悸����'ѻ���~��d�?C]�i��#�<r��[��ʱ���D�h;|@�t���]�^;��;p�:b�&����bS��LG1���+�i�6=#��{����èoM�C���B[�?p�A��І�a�O��Ֆ�����K+4�?�'�[���� Es��i0�;�jŭ�:���2���j��;�al#���{ݱ��;�ϑE����C�	v��7ɭ��k&��wV����4-5ƙ+~�.���Jw�	��&H�8f��&$�|]�E��
�K�"� ���I|@OR�c�N��@z��!�O1�!�4,�#���r�i�ѷ��EG
�M%v������J�|X/Y��NY/��f�0y�W�Y�A�gu�v� +7;�s����&olޓ{�{h+�'"�+U4Ì� 7,L�n�)�6i�R��hs�߲xv��?"�!�ș�H<�Hȃ�n����j��F���0b�"�P��᝙~��H,��N�����ӛ)dض�&���N�A�=~�={�l��Nl�` yR��#�q��c�S�	� �\* ��9;Q�����c�el�n�Sީ�(5��TqR|�kqvLg+8u3\�[���ac���4�H(�!�������x 'Ǌ�t�~}��Cj��4|�}���p���I+�Iy�9�x��%[׆^n���8yk��&�fޑb��PwF���aO}��Q��˺���~#)9W���y����� 몴�����9vt��ca�ħ6�f���kW�a�������1�Q��Nۺ"�JJ�=�$���W�l|;F�d8E�<2��T��>��v����6��ףE�"�~�o���>�g~۞Ǒ���d4��*��&W}U⨞�<n$��d6[ݸ�1��}vҢ�'`��������	�<�E�:X��*��?�yA���̖�����|���tV��@S4H�#69��ȥ�jI�ʼ0}\3���{�
�_Q���8�T_��~��N�� /ԯ�J ����� �y�H�x�UxOY`�F��6Y��\���e�U#��Ek�F����(�(����RB�A-H�pmבk�!��FJ�yV\�{��џrvh�/z@>(�����ޭ��S���(���Z��W��~��ݞ�r3\n����^����c}�¹F��Q�h��n	��Z(F繋�b�;u꠫UXQe�w�������P��5Z�g��-�RKI�|�G��Ku��b��<xv�����6�v��L�j����5ᰈk�T�n���B�^�U��0��+�;2	�?x���D#�b!P�����~�u��Z-^�R᭷{B��
�1�i������'�9�"B+��"L�Śv��D*�+���ֳ\G�R�K�2C�I��]t#^���Ǒ��K߮�s��[(�r�|,�W�a�x1�}_�i=���WB޺��^����Et^`�;F-	���	s��'-��F`@a�wZ܂��7+ԨՐ���3D^�UW0��:o�xQ8D����N�`�42�@�|���U1\CEAMt�F���'�o��y�+�y]⚜fS)�m����f��5~I_OI���ǎ�W��WP%e7HPut��MfvO�pqr�a[�?��w���r_	�*ݒ�a��ppl�?���̞�w��6�3s#}A&�nz���ݩ;��X�&s���86����\G�.A��ûXڝvGR@L�϶�K����	`�(5�0��l!�k��Ґ��W��Of�7DN5+���\��Iϊ���:���y\$��0̦αZ�g/����3uH۳�;R}�?X0�8�M���cG�#RnP(~��R���5�<���{�y��Ev������ �m��o�~ޡN֧�r,�*�{�ɖV禸5iU �A�,��¼�l3#�3w����oN�+ׯ���XEdS�:�a���d�~��@�-���l�%gxS��GP��:gD"�D�Av� �������� �Ǌ����L���Qd��s���sF �z���;�|�O��>�9:'�����ܤJHIy�޺_.~v����q�	<3ZeXHE}o:����0��a�S헼�NC�� S�N����`Z�,O"v�GK#�����/�fp6��gN���VO�6��A���o|��ǜ�M1��H-��d&����o�TR7���]g���Z�aV>�pj*[Km*������w�t�4C�q�^�R�GKu���;]��fe���]�͕r�tE�Y�5��m�Z񀙆	�L�������~���������~���9iT��H\wl�t]J)D]�V�]qQ�4�U�V;����v�Y%�<H����qw���K��.I#G���/fؕ����5���<c�>Q�f�h���@�=!pa6*@�-������yXRQP�uz���i�� po���$w7�$�0�{A�<����
Rݩ�t���}�h�#����-�z߶�!��@ܯ{m-�yo7�GLsn?-��)8�]C2$ω��`c�.M���OR V�������E��S�+�Hث����S�= {M�vH6����߿P���>N܄�Gr��Z���y��&cE����/��	�`�v��cW�T�kCPB�pI�W�ے<��`?����BD��t�si
�Jy=J�������;��L4,\�$��,�����t���4�>O�d�l�� k?7���N:��i�K=��0�z:����n&����ҍ�����ѻ\�߾ٚ�m�q\�����&q�& �ON�o���OX��Ӡ���?H���|��w#�HUs(M��@nTQj��e}���O;�P�vP���(Ò�g�{M�To��c0�}�-m9I�����|��G�pr�[��`�@�	q��Ɔ�3���ն�h564>ޗ@#{��o�������c�����.�%/ ��VUf��сdD�T����p9&8���1��ŊՁ�6+d�t �Cʙ��>:�xs:�a�.��U�i<K9�#uJ3g<~�^Q��c�4���I�9���3u�N�TΟT�`��c��,pzC��O ��Od�8�b�2o%<e�����M~���p?�2��4�@��3�(�,�2 ��{|;�	��HoE����2��7��UW	�Di[�%�"C%3�:*oJ�)���T��u�#�Q0X�[��hD)46�  ~w	y$�h����I4b
��X�W+aN쵹�����M �}��ݎd�"')?R�����*�^OJ��
r6�D��v�)��)�.Ym����� ^�!^���x!���~��ŷ��G:��Kعk6W�DA����#��������q�T��G_�����6-ݹ��X6X���E֘!��؃��|�ӧ�\��r��l�*�k`���7P2w�q&�ibda���U�$��po^n�a����j�喆hH�����Es�-?�֪ d�����8��t���x��U`A�lWT�A��	�&D��\����c�q��{�quќ_h/�rK$`�GY�D*�~����m�fAK!��l|P����ސ�)��t����yU�N�������2)�C׀�"1�D�&��<�g�%�AL�4������s*Lݫ~<��T�Ҧ���-��-}`�Χ��o�w5e��-��$VORK9Q���__���̯*�>7���9�[��(�)��V<XC�f�$ƞ$���i��i%����-9W�+R�	W �<>�� ��N?���]TE��bM���K���Ơ�/<T�&��;��#bc�h,�u����\c�bp��Z�f�fjY8��w���&�lQ���
X�ׅ>���ѐNn�#@���M�.a{7�/A��t��9� ��H���jw,��Dę�a��X��#�.�t��s�/���*�y/q��:'CٷW��$$ ݊�Ћ	�Q�\g��J8tqL�u���Ő@"(Z�2���x���Q\Au��_��fn=�*����*&����K���Z���U�ܼu���#߮�@X땓�.-�A̟U:�BV�Q�9�ry`N�(#nwc�3��(6[|���C	M�1��(��`C�����)I��P|�'���Z��"�dNYG���;�"+St>��*n�c!���pG�0ky�V�[h�x��(������TAf����r���3�ȉ�8]�5�;��#l�yPq'w�K�C�Y��c���}��cW��-��Q��ru��0��o���*���1h�B'M�k�e�@"S,�4��p�892��
d��"�ĺ�ԡ�M���!{����.K֛ tEZ�nG�V����\1�PCc�/#�QQ#�[��� �?ca�+�
�2�������@�����i<�ھ��ݟ��	�,o���&`���㶚�)⸋� Ӆ��#d� Ly�*"��T��}��W��W}����
z�����W��k�M���@l�ok�&�"�
�ICЕ��I4G>	^'��T2��v���`��A4���tx��G��	��t-��34�E��b3��5��Q��b�x7�b��<Jԍi���a�[�7\
�ũ�����4g�@v���!��&��.F����_h8��G�g�Y:ELޙyG�:bf{m��w[7�r_�X��
��)��'D��ևA��*���Mo��� �9�G�i�����lK��qOzF�^�g��h�(\��TjY���=�=�{.;�v����st�����4��6�R�8{Ĳ�4z/���r�$P�P���ø΂Q��ē�O�Jv�9���WM@��*�"Jz����L9��l�}�M#�4�����%6|�O�B�Rُ��U�؞�������:�����o��J^�$z��Sچ���L��$�Y6AB�m�.�Zs�ȑq���O�<��*���=�O�an^u�}KBkQ�����Z/?���5f��@�f���PbS���Z�E��W���ƿ�6)����QM��@�1��2���9�A�~O4���t=�h]��*�p#H�:SͶ9����V�|[�Q\��N��f&A���{���o��r�t�R�)��N�G�l�Z��|�"��������߮��)k���F���z���rT�F���C)\����k��}��-���ju`��u�&��u��I��n����m�T6���1`�J���TE\�Sr\c�����d=�m+����D.���ɤ����[��җqmK�,<S1:�7��k�z�"6h����"��=U�6�a�B .�������_�L)(����r{*!�ք��4����́ؗz(�)4ګc%�Y;��K��3�sW*��N-B託\jʄ���Ω�U�!̖te0�O��d�� 1z�R���#��=���F�(rN''C��	��v�ݡGQ��Q��U�4&)`�A/�9����H�w�5z���T�A�AlW�p[���� ��,�r�#IX{o�eȄD�B�
�N�Ruq��"��L=��ڵe��[H��i�B��9�*?��d9z�@��}��oN	x�E%����Ml�����I^U�yXo��y!�]ɢ�dLbץ�C����8��n?�E��L��6*�
Ʌ$��*�-G6ݡ bI,MUA���缺'�5J#��g��Y���k�:��b*���J*p�v��dwT��Jwӝ�c�LV�伯0�;7�4�[�q �_#�S��!�R�����W8���x�PC�Է�c�_VuH'��9�ϔ,T .�@&���bم̱�y��+����Q�!�Ш�нS�EO�.u�x�u7����WG\�՘�~%�8��qgL�.ְW_Y���Y������	�\e�oɂ�J��
�l�C��%nr��4]Xz>C��Odo�y�UE?�hx�#�GJAl97�:��,���P]�K�H�+��ǵsD(�9��Tհ�'�y�e9�2-��Y(�����6���ـ�a]4��`~N��;R���-8C��R�pN�`¾�%���=�J
����z��]��� �UD�#�/	�ڽC>��b��&�����E��
�4���ƁzcO���w�g8P!�M��-M�j8����0dn����~%�ŵdf�oЏ�]�+���(Q��?{�(�D�}_�ܸ��w������ۦ�"]�3E�*������d�;
��G�7�����FW�xׇ� )fo2/�q��e��8�Hl4�T�" ��AaSRm�_j;s� �}�vk���:�9��X�\?���GtㆪL�Xc�a{�Z�P4�D{ʪ���u���	�-@��85�k����6rY��d�8%�A���hS8�VӇ���y/�N �3y���ǁ0͐�2��݉� pf �P��:10����w(4��A��bcHaH���{ͻ�	������qISJ�[b�F�6�
�[��0�j����P�Ț@�0�	'�w��eM֭�����^Ƅ���.��=���J-�U�o���`���d�t��!�~�SW�AS����k��y�E�RQ�+8@���vC���W�g�V���74�rT��W�]�__奃-W���7�Xm�?���ӓH�ȧ��ù��R�vƎ��)1'�-�A��/ŗ ��1��0ӑ��=������)�!���u��qS���zPJ�Xúq �zk������U���еx����O�F'�>i�B�jG(�3�M5@�y�y�+F0 1�������cY����;�vb�kDe�n*�=	e��J����JPzw�Y�G=|uo:�N`A��_���K�@���q5����/�V�];���,cir���=$�M��!V�g��l���5������
38����F��i-׵����5��-)�����16�k�N�S�����	��YOI;�P�2�R�W����h̪K��_l)����$�p�e��9��b@t*�g��ͷ���M��kM��"�:��K"�	��,T��U��{�� �k��U��A��#`�d#t���8JL��m��c��`���?���H�%�fK��n����K�$[�'7P��.��������#%nhU�C�,��Oް���Z/���H�Iq�%���`�2�?�8+��b�G�7��o�*��LH����rh�q�ʆ�o�G�^>����址�"Z���U������ʂح<0�F:��*��Ũ�b��'��PKg��iu��NAC�,$7��c�8Z@�Q��Bl��̍9�9�0?5��,`�����H^��6��`"�8]E\�:�~7D�$`����z�I2�"Gd�z=��XS�D!R�S�P�X�9�����ja4����]�#�>s���ja��c���L"k��5�C��+t�L�'��ӝ/��H�Y��Y.��{����r�l%�i3��w�4�|�_�[}�#�S�R��,�D5K�?W/��75l����Y?D��p2z��G���JӮ�}Q��H�%'���������Hz�dz�ab<?5"E����d#Za��$}$o7	u`�֕�s�p�v��:vв;0 Z�݁i����ݳ����s^�� ~��,�G
���Q�^d+_�ę���9c�F�ߝajGN9aƝ�8r���*��nF���92J	�;��i�8Y����J�x�bKB?�AU ��h=k�����A���ͼ�=�7+�_.O��O�r�Z]I5:R���3�"n@�:D�YR�z�8���},�ȝ+1m}01@0�M�e�9m%��XCr��ް�/Ds�ִd2M����Apu�q�w.a��*���^!��]�	�Wo���V�	�s�������9�8L���V9���	I��j ���-�]]���8���'������(B���h�3��)��E
�.�������2�Y�'�[3��AȜ��}Λ�i���3���ߴ�60!Oא����ߕB��Ab�˥L��uz�jߖ�r��ִ03qS���f�������f_&���A����Mms
N�ЁQ���mO�8a��x8-�_�r�d���u\��Вꦼ�uz �ޑ�5�M�6��O�������7��uD�����-�x�K�����X1�oV����cST|{��;E�@�SbȞ�0 =�y��j��\.�\N��Z��LD�b��$1�#��^�������5FD�5$�{Sp��h�L	���p����h�5����)r��%�rW�nX�E�s5Crk���[�\.����NX��Ǒ��=�"��,m�V��FWj�&i@'�H[R���Xe��	��O�Vb��v�g���b�*J�� K�"r���N���x�ϓӈk0&t�L���$�k�fr/���eՋ�]T�����;=�a4��#�xv��U�\�����5��G��ɓld�雏�fV���U��A���N�ඹVJS�eu
�' n����o�,G���@��`fd%_����Z�?��$VE���O����_��>�g$�.H�=�dϷ��ag�I��Q�v��ƗC���Xz�{�0�sjI/ ��E���QOlz���x��������؂��H"�}jQ���pTN�ؔv�g�5����1)J5W����
�Û�	{7�m^N�p�s�~5�~��1|�hl)0�b�'Ӫx�n@np-8H;��=�&��&�7u&��R
.t�{̸���¹Q�@��ʺep˰�s��W�l�L��+
��1�~�s���X{<ݳ0��G������R�"��pt\�ǁӟ:sA喔�镌�o<3�>��o�'���i�DF�������E�N�(w�^�vf��O����	�I%G��lJ��8��l��G�J���iKk��PxVFd;ux��4���
��H��Y�j#�m�H�?��gA{Q��h����Nd,*aW�U>/�n�^w%l�VU���ex�>�Ͼ-\^XX��0���l�w��0wm������t����d�8��A@h�ѝ̵��M
��Wg�Dw�� ����oq1Pߧ~�T3�坝���됬h����p�l^�R���&�PM����V<�f�\�7�� 0߆��5��z	��	�U����Y���_��A�d�2Q)jp�������zP�.���&+-?��%��'�O��|qW��:��Sc�W�h
W^�p� �'�yv�s�$Dzw:L���]D5��V�h���*�a��V�w�,�O�|(�u�ʈtK̊�S��QGAc����g?�a�����I��P�G�v`q����p�?��˝�VK�����{w���_nɧ3��ƪJZ��b��9qcVT(�X(AA�c� }j�T�AE���ȫ��xw:�HQ�k#�
A=0�hh���20	bƫ�n�b�%���S֗�S��	����F4B�EO��6x�5s����q9NY_)#SrI��ɋ*s������7��U5C���#Uz�˰2����OĜ�Ct�f�U>E����`^M���`��j���Yc%I�哺�$,l��@t� ���I���VS5m���?�x���֙�Hb���Z �В�F�O"�E�eA2Zp������IW��h��D9��1_���h�c���D���^;��o7���`LY#r�>S}���NW����i�Js�GU�о��5�����/Ӕ�ˢ�-b<Ȗ�N�3D�����*=2V��s���yU�\V>�5�4���<���������� �$�����2<���?=�@��F�&�0}R���?S}k���y�?ϊ��d�P��r�����3�ivQV��[*� [Y�&�;�e�z��Р�Y�L���@t� ��jh-��r�e-_ ,t�߃�J������5>�D5�����*I�+[{!���R���K���ٞ�-7�uc+�C���K��F ��'��!�I�\��ű����Th�ёK9��P�8f-����}�1����ju�r���E�/@e���7$�o6l��;0�����TC��V����u
��qu{�
B�%���%�h�'�ӈ $�&!}�ߡ�B�N�x�%D���,Wx��M��w�=�f��w��7��E���y�XV�ꢫ�%<��2Y���q���7$ҵ� ��!��������\��ԛA�p��\Cp��]K�=1�pV}N��#P�b��f
s;�&�V���PYuz��|*��qQ]�*��h<lUD;��e�F�4U'��qt�ɛ�T��-��6
3F��v�,>���Z��}��_�|1��{`	���i���l�N�+�G��\���@q��b]�ϔy�b&a��Zd�h����J���A�����+rE�.Qi&��qP�85�{�D$�7kD[i�l ��e��Ci�`�!�/;��H�휍(Ƥ��A�|6�����m?^|vDv����Z��V:L~���&�����2���iSe{�D��Y�?g�mb�5A������b�� �/Rv�0̑��r�t�g`�P?��V��I�z/%�|<F>��󬲨��ݜ��i1:|���N?�a�p���?\,��-"�� 2�uK�-#��������+L,����΋Ƈ8��H�E��ޖ��X�<�0��sw��
��Lŷ�����FsD�Q/wt�Wm��莆�,z$z�b���Ri��biv�� ��:v��Nj�nro�9-v��5YJ�|Ջ�8������Q�W�t��F]}9�H+�<D!g^G�Ϋ�	^>�|7��>z/J���1���AT�>��5]5N��%p:�.[`I!cX�avŸ2ٹ��H ���D|ZN��t_E�-HCנ���@�q�J
2(y�@e�41a�:�����h�	oD�Rpʳ���ҟ�"	�)�>��̰Ph|l��� ����f
&��|�;��FU�*��B�Yxg�vwz�s��}Z빋=5�j�d�=$[�i+� �іǲg���9~"d���b��
a"_�v�;�U���Om���Q< �6Ď?�M�S;e;2�;p��"��Cw��6R#�̐��4�����_�5��v҄OE��-s�2溞D�V>Npm�.����ެ�,ı��6t�~6�V�<���KjBY5;'.A���n�n_89^m!��X7���5/!c�g�aj��ӳ���po�nD]�QS���W �&:)�G�p�/�[�Ϧ�W.�7[ƛ^�U<>��68�6�%k|��v.B��h�=����AX�)ԁ�V>��\	������d&�:�u�y�g��&��\7����Y��e'i�	���y��n�_����'޴�����[x+ܷ��+\(l�0�����7���*
Uv5���݁��Қpl����\LWA��s��N
f~��öe����oZV�5F7*�v�����|�(�ry�tL�#���:�t��/�Z��!}���6�Nr4	��$��M�q�/��x���a��2 ����CPy�H���Ü�����fK�q�5�������� ����B��z�$�a_!,����:m�_7�K�}����T��[�vi�.��b�^�w߮^t�,!��=~3aRT��sQ���z��H��C,.2M4�U�#p�m�'Ș��dq~���s���C�rv�/�k-��t�Ѻ�:�z�`�V��?�}�k�Xа$9��[�s�����X��2x�b �w+�)ǩ:�Vy�{���UY��J����^W�ؓ[;��};vl������b�۬���0�e�Ja��EB���wG3���v?���0㓘,�jX���4�<��A�f���$�A��XACP5Pځ㮿�gl}G &�
ka�2�6H�x��Q���t�� ��C���Rh�>���o��"a�X�ѷؙa��Ȅ�u�������x�i�іz���A�ձ�oc�[��m޾��sc6����d�G� sŘ6N��wGG%���+��rP��,�2ju���t&^�u��%ϡ�x��Q�v	h��G*�AHz��LX!��v���}0�j��*ş�Gn�_�z�E=� �H=0 �&���r���-�7���K��C�͆$V�|~*���`�]$�Ow��cٹ �ZI��#W۰Q�ZB����C"@Z�W'{F�l��-�Wz�"/>���$
,)=�W|$w��^d�+x(�2:�T�4�B3��qv�¼��K�DWTPT ��P�ɻ�JY��?:���9+7��-7�Ŕ�-��o�_����5$�+��AH��F[�*�R�er�u8_���|*�I�Q�l2�e�"?Z�8�(���D��O/�O](�ٯ+��n�f�Xׇ�Ĭ*���|�Z���@�O����|:��\�>��%~����炐uي{Bԃ�)�.0����J��Se6 ��vb8����)GF~!
f�����D���:D߳��Q��B������_�	���==�1M��4]N}������.�Pބ��rcq��L̽wI.W�|y�%m�@B	�C��/�2�;�o����QR�{��`/U"D�<�z� {4\�@���1j?K�3�wE��L����ڠ���`�乿ӭK⤉�g&�'��Z����`� Q�P�� {��b�{,
������M�%;b�o℘S`�<��[ k�������P�B̎Za+<��b�L�x�"��,�G��bȈ�e��U�8 T/X�Pz�,Fc�ϒx$��x�(�	&�7�|xŐ���y��_�KW���9����"��nT#���D�f=76!D��xO��B������K���+��b��*uR�Dΐ�"T�{�Oq�L��9��I�'�&7��۵�{�C�2�Ļ�0���-pl���5'L�l�ɜ��C"��<��k�/�y�>)�l�"�{s#���V�	,�i\�q�d�ϗj$�<G�k,�tþ��X=�^t,8�sW�Ѓ�Ip)r���Q��|�=+���"��0�ozr����:�p���������Yy="mϻ>�4e�,"t"6$���Nڏ��J��B'�HQTW|�����^E��ʡ%�I��i��|�2��(ԯ���k�m��.���!/v�� �e$Z`�O	��ѭ�@�=�9E�M+��@�m(4�H��-�B�h�Nt`\h9�*��e�p&��1	.�˥�cq��;&�9>�}��f�����V/��z �����AR�:,��1[�Gh�&�,9fFjNЄ?a=\���f ���AxeE뼑�D��Dt�������yET�(�%Z���yʝcI���>0�=WU�,!uO��;z7�U.�� �~aEx�4ÐIe�](x|p�D���b%�R�i�A;o���p���`�	�{�� ��|Z(l���X��;�kY�hKD�w�R��Z�ʍ�Z_)�2R+�O�B+��B�dǍ���|r���uu���2?&�.�E�=`1ib+�#���jKl�P��N�2�c�&��9���k���b:	�g�Fq���^�;��܋Q���u����fO��F�o]4^�:��f>�ݰ7*Vˏ�m�,m:�,Խ�S�b7#� ���Ռ|TZ@Y��u�X�]�ݦ�L���ā5�l����Y�2Gs��U�{���D�*-)W���go�K�b���g��K.Ò�+ ��s2�v�'�8ql�D� �'��#7sU�����H�z358�Ѥ�Y��V���b�H�jUd�Q�ޤ�����>+������BrS�*v� ����B���#U<Bx��~T��G�=P�1B\fu�ʭg/=���e�t�@��I4�D�;��i�h6	���|إ�Y��u�#�ԣ��ر�ϣ��V�S8]<�u.[p>3�!���\t	kkM�֏[��e4��H�ǅ�fd<G��n���#�� �K���(HLJ��Ĉ��RMiZ�
U5a��Wٕ��6��b�EҨ�U2<�NٸP�]o]�҃L��vog��
c�P�r����m�PS����宯b�s���1�}�c̮��O�]x��K���r(��QM�l���Ԗ��_kJ:��V�*�v�u���5?إ}]&T����O��f����Vg:�| �=��_t�d�[��Z�ESvnw��ѰEU/ifKɐ�k�Y���v�ߵ����}�B��d� ���8N�Vj $�eh2�&ϛ ����,+�ɝp�˄����*��xI����ĳ�t��:����Tb�1��3������H���'����#��i�t� .r��md#�]�` ���]�,AԀb��?�۪u�wݬ�=�)Z5�B^�7N����%�F���3j�o҇���I8^ՄWP�*-�pא^�8�=��Eg��`��ފAX� �2�g�(�k=��
SiK!~����S3�a�[�\%'7��
�1+����6zn�6<^��_�>zA����2�H�RH6��y��qVe�;,ph���e�PU�J��`n���^�5u�T�r4�L���>
9&e��HC4q�zi��w�Ӿc�Ax�5P�c�PZL*�><���8N����%ܢ��4vn9gOt���2W���@�q��.Q3-j]�I��(���K�2��WX
���G��/��B�*�x�$�ju��F�;�f�z�9e�y�ް()�0/�ٚ	I5�"��cʚ�^��j�7n�"���y�����M��^Ł��y�֏��`K��֚/�j]5�g�HJ��A��VxW��3��-_h�:����`��fpݷo�}���|]uEiMI�#�����Žm1g,�n�5��I�����<�';k�F��fM�(��6�g��挏�芵�١%��.���*;Z"
�$
��kM�»M��r$b�
1@��7�YP�E�K��
 �q�:Ǥ��r�ӭ��mԗl��}E�p��Cn)���m��i��Ad"�S��D	��r���D��{���K�p�|��;��fo��j6k�y{�iE�{h��3C��֥��5�OX7��a q�+nۚ�"㘫��}*�+3%��Y;쬕��cQL0�]�����n4_�w��f�?
�G1�O���r���m_^z�Lh��`�J8)�I��gy^^�z7b��{��8f�F[d�2�W�P+�gº���>�Kp������������g�DP���<�F�H���K���� � 1]Yx!z|��.���N(����D����\������PJ!� �+�ב��O31j�P�jyH
r?܈c���
�P���=e�Mk�ݐ�(�lDGK�?D��:i�'����4���@�29����"-[� ��[
�ޏ��nf,�.׿�*W��uE��lb6EűY�0V��O��-ீ�,L��m����!�d��h��1o�o��_��j��|�d`��k;_h1��ւR�dD���$)��
 ?+��UT�q�ՕQC�<�n�A���n���2'#����	�S'A~�:��Z|�?l�U^��b��i\��({ڌ>+�NK���k[ �3�����+~�k�7S���Q��?A,��VX[�|%:�����j2��O�e+Q�S^8�o����>WR�&���o<*��i�TY22a+��Ģ��g�z��@v�C��O&}����M\�Q��>����*�#���1aDi�"%���Px�\�?(����z�|%ݼ���s�E�G��͒�.w� ��>�,OЬ\��;`kmI[�/��w�%���W�V��Q9�A0�uK4k�C�=��̥<�������<���}�JVۇ�\2Q��9&`���3�0�u������I:���ƫxE���kDas�8����ݵ�=�$,�]Ѵ��#,�7N��N[Y̕�P�|O�,�r���ڌ����e��̭���t�X�roQ�m�m�$�K\�k����$^�x@cw�����D �~�s7e�˜�X��H�4�k��d<G5�݅�,ʊ7k`�
�G\�IU���\cm{N�1A�N?���Y\e�5�@*���p8}�nj�0��?gQ+��`c�-3�FY�/�|��$S���U*`�)�j��BKC�(U^�#�k|�l!#��U�:\��V1����W�qf��9�>(ד8�'7�h������ �ǣҠ��B���k�ӽ��@�����q+����`g���S�wHx�Ivѓ����W��<n����ŧ�*C�17��`�̊`8���-t��1(�$��c��"]d���Jz�+C�uz7��<]��f��|X͖�c�ܘ��Vg}mk�c&�w^��ު��P��yM�� Et5�`�*q�)���n�D�n��L��.�b#�?7tfP ui9�47Y��Yy$�̽*�x�y�WN[*T�Nɋ=�,Ґ��1c��!���O���]��v��'C�#Ӽ8�f\U�傴�	3��U^א��P��1<��~b3�_������^Q����Q�Lkw��oy�E�b*r'|x ǌ�"�6���E�9Ĺ�[�xdS��x&��I�_rL`
D2��P�+ �\
�����8d*�q��ꊘ&�r(v�#��7@#�m�����9o_���&{f�7��F��-��"Oo=Vhk�:�7/���g;��^{��+)��,�ա`��������I�;+�12C��^�Bq������ nٞ,�CR6�Z��B���5W,�J�L֣�¢����Ӄ��A�2JK��鸦_�\������k� �I��B�&�C�3��o�����2��QH���J�c�׮���B̀�r��?D���iہ��;����AU��F�_-�� f�]�KCl�>V��0;^<�	�RýL����U��rk����p��텷���@`�#CIT4�Z�~'"�pz.I.{9q���H���jP*D�'�{��Ϳ���ћ���N�j\֋��E��7�&WAq�)��<�s�ʢ����{�B�0y{�e�A\���C=)�l�북�z1�s��gV�u�"RD'�v�U^�����SŔ�����E>6<�)"9��c���:�pL�N����^��0�SO�T�zxs�0�7zt��J�6�6ܹ�[����$��Y0�J�ߜv!�t�Ңbv�P����d�8�Dw�_с�&��;CG�U�Ì�}�d��9��N��J���#�bC�>̃���5�v�X�؟$N2 �����˖��?�ҿ�� �$�ͱe*⧶<�s�D�RE�j���]����ѳױ+bv�����a}���;w���y��U:�B{J1W*?� N��������YEȟb���Q�!��5��B�Nb�s������O������rB�U^��M� �+��Ϛ�E�T���"�"r�$�-���aj�ϯ;`��d����!�9��'�nw~%����˿{��i2�/��I~���	h�w�|�^��T,`�#Ge6���4}ω�qp��.V�>5��%��ƢI�,2�+_�^�H�Oj��YFJ���뼃4� ��I_kݐ՞�"��������V�ǝ+�)Ç]���BL��;E��?�
64��#��tp�}_���U�h#Җ�$�o�:���/�bV�Zi@�ޕ6�N�{���c������\��>rm5Đ�����\�x���˞cq\�-����viL������#x�a�4Qp� ��A�m�y9��#gU$� �E��g\�x����3%���R��s9��Q�v��f�c�X92�k^(��@��J�y��9��*Y�?�+w�j�*1�0P�9���yDM�Py���?�u����`�U��Q}�OT��s�~d�R��	#��8�j�DLR�d�{MA�:�h��E^���R�͍c�����^��Z�$K����o�Npo�jϦla��	G�?M�!+3�!ڡ��y�R}��$�.����i�A�ʔ��o�T�'�l�rZ���|�*b����â�(��u~=����GϷb��k��V����;�pK|�F1�"G�Ƙ��?��0����1�X0F�|fN2��Q�zX�;  *3S��6�nJDe��w&	����ɉ��.bқJ��b�F�Y��"��Ǉ���VI�K4���c^H���'PCώ��B��1@������m,���T�T�8k�j�.����/×c��h���4�#.1~����)����v���HM��3�<���a��pu�1U.�������Zz��⼆��� ฽� ��]���aZW�\�a�D����W��c�|{��e�|�!:�=�k��c+̭6��jgm�#�O���
F�.`o4Q�|�Yn�����QM�<�]r͗¿�1fQ��^0���jv��閁̿��C7J�<���}H���q6H�\(S��h���=h ��3�URngz�qD6[y~���V�#�g�f�l��ı�3��B�����K���Ϧ9lر~�ޙ�a��q��}�\���o��)�u���h&���7?9�sx�s7a;�(�Z�QB�%}��d���k�R8�������iC�4!<�v�������Yp#Y{H7=ͷo2r<�O$ag|�U�!���]���ͩ�e4�To7d �x�P����(j$��N�U���M���:WO�k;��F���M�����#�)�c�:�j��e-$9����?��+���v�)�ҫh��0�k���@�B�ޣ��z�6�2����x܄'_lh	��(}�����O�[��TS
�w�XJ$#�Ƕp�����E�Ykiׇv������P@N�V���#�8	�������WD�+;7&'�4��N4���)Z� ��w��aU���}u�WS�� �����Q���C�>�T9�.��[?V)�h�q$��g�I����s8�Yf��g�
�w�l.
Χ���		8���tZV�ӡ\}�0�I��g}�or����j���9m2w�0P�|e��;[ ����_����.��Q�M�[����A��ʃ�=�a�y^�:�����9�HÑ�g��ٵR�P}f�@�\��l�����<��<1X�
^;�.a��P~$���k2S>�����7V�@��ϏJ9x�Ӊ�3j|a9P�.�^��J�Ws��t4ාvq�.8�)o�P�J�?�.<�g�Psv2ƳÝY�B� ���'�l���B�m�
�4C���>�C&΄	��y�Dh���B-�����ǂ@M�_�/@$g�w����F��-���;�D�wKݦi;`iW�MQq���Tp%��Ls8r�{����hd�x� �Vp��Y����8Ē<M�əpKA� ����f����eָz3`�s�	�h?`���g�ߚ�v�A���q�����5�K��(@Bx��d�b�ix���d�)9�aJ,Hw��1���P����$�ZO�5�����F��pN�Y#ʯ�,��X`�(����/f��-@�~r���[�XyK|����dب~�����%r���A8s�Cg��,�s1�<����Ե���p����q��é*�j���HΊ\���2�R[���zS�ڑT��{�U���mΊ�1꿍��b{Gu����^��v�a�K �X��w{�����:]OA�#�;6E�Y8���<�W�0V7z��ӳA.لA�/S ������Ͷ��P���A;�V��E�,Q"_��MGF�N�9�o�Wҹ=v�)�U+���cF�N�xRǠ��R�`�V���$�hˠ3[�&��������LP	eW�)�j0�!�h�ª���g!�L_X�.��A��At�G��[��s�,�Y0ٶ��oKѣam�-���c�AC�s��Ę|�sL\&���ӯ�{�C����8��3WA/�ߛ�l��l[S"��ExJ	���%XE툉>���9��Q�5�3οW��|�+��ķ�c���O���.̦3P߈��DhR<׹OZ�T�ĝ��_���f_����qgWƢ�<����W����K�.����:� ����
݄IS����p���|��WN���"���"��_�e��ނ6!K%��J�_,, ��\>݉�^��?�+�&]�A��D$��=k��]��<�{R;��B�����14	(����n^8$��ӶQ���3?��L�r��-��gN�֥A��t�Z��X�\Ap,N�^-6�7S�8�AI��}�1=mY^'^�H�@�h�BU���S[���MD�:�u�w���E�Nn2b�0��o9����|��|�$SE����奣����A�Z{���Lh��=�d|v����BO�Ј���� �bY���ˣ=]���xݺ�֭zIw,���]A�p�ϵ��C/YL�Fk֍=�s�����$�<�Pv��C�۸��'?�Mwi�%^7��fx&��T)j��/�cp�v��� �ƭ�R�*c��v�_�&t\�ͳa^�2�Qq�f�ͦј���`��V8U+ �Y䃡uE��B\`B'��Ï�}�?ěT��o4X�Ą�>���s|��ϐ�K�V��ъ��JK1߀��(�p?�*��8�[�l�
:�G5倭���&������@�G�4�g�s�ą�ɜE���ⶣ썡,��7��ئSXK���pN�v	��<�	$�gΪ��k}�#���;��Hn��R�f����
%+H���'�$d�}z�uẚ��E���i�hrG�N���`[��Fm��6 �jIh�gtM�F��C�fc��/���Ō�����o]�]�=Q�Q�g��D��x��z�\g�ϭ�?n_(��O� .C���+���u\+��pi׳|�O�\�Ð9��PIXY��6��EZv��C�YLm�e��Ҡ�*<�B7����%%�>�w1������.njԢLO�<�k(ႜO'���t/s�]�V�r嘮I������T}�M����8\�29<�Q�"�����点�R����K^:U����j7|�x <`ت-��Ɔ��o�G4냇��eZ��}��y�&/�؞m5�@���%��~޿���b�A����J�&����?&��E*��-�4��qY�A���ϝ!�ӷw�+�x �˧H�^C��Kp�F%����@�xib��\������Nz�R��<����Ę�����\��Hus�cE�B��B��JD�� *c�0!�C?,$\��n�ѷI򚧫9��(��L2�'a�RJ�n��?5S����}���h�rE�֑�*h0s��O|��T_�bp��8��o+}�#��e5Z��Ǩ뷸O֟�q�ǃ��>x&�X�z�6=g���d.�
���Y���T� *6�I��n�h�xV�����ۚE��j:�XÍ6�.�_����h�9Wޠ���^ҊF��Kn��T���^�e����u%bb˕�̧5%��,�R��9�s�)��H'��
�2����Y~~q?U�:.�u6���SYK��&�9��c���3����?*��X�܁Ń$����\fZq����I>_@������t��Zi�2��(R��w�TJt��9liȸ_�:4S�O#YIc)M�-�Fݶ!>�����[0�+���3W#9���_�
ܑ�{�����Źq>f�X\y�?y_`\m��]�O��mCa��uK�4
/�@1J�C����TY�Ķ��H�Э�|IUJ)�_�	{�a�	\0:c?	=W��;IC�%� �cBb�ܕ�TJe�ߒ��H"-�����X�m��{��Q�!��ͺB�a 8\���N��+�޶��I��Ȩ�>r�p��ôU��51�ן�W҃m��~Ř�ϸ�.$�E����X
x2�X����a����	�#�����3�mм��[�������j�W._\);���w4Xp�*J����Y����D��b��d|��oDgP�L�!�]L�s��ڐ��h�OcIU2'id9��LE�I߈85�]/��ۇ֮m���g�]Ծq`�q-D9h�Kr�a���#�q�Pn:��*^ZG���TU�Ǉ�ܒ��7�*_YEZ@;�ю3��b���q}��v"����%�Ί���f�M�른~?�!��C|߰��O���H����>��\�r  �^���G���K��H�:�vS��Kͣ>��VQs�q�'��sa�zV�� b�9!F��Z���jקSЂ�����Kn�!��6��L)=��R�ch�S�ɲ-T�-�58�*��	pS���C��N�]Bh�4+�}q���#�O��9 M���M�Crp�Wv9N�򔠣a����z2Z��5���L��CA��Lp���p����&�:���C_�2%�PbB��?�$�0?������䕨����Je}���/cy��}3K�� v��-�X���]��`�ZM�7��g?��T���} \fD�<���b,��ܳ�9Ϟ�L��4�ʕb�W-���C8����)'>�p6!1*��+=�Kp� L�2�\R6�,�̴ڝ�A�`\�C;����ˮ�C�f��(�`q��J�f2Qϕc�Ӡ�����(���N���v���#���/�D2?�iD��`�pna�:5�a�~Q��{q��{M~�� ��v�2f
Z��A�mٻI>G���)�6���%i�ګ�b4y����]d��u��e[e��t�ґM�h�S&>8���~+��?�U���r��E�y瞒Ôjf��s �c@��N���H�=%s �N���Y�uq��熚��D!`i�y��(�6ϥ^<׏�\L����z%�Ť���kw���\��P�������!�����dp�v1E�6��R��Ѭ|v8�K#itk`܃+`wb��������?�ƅ"&�c	&'����d:(s;�mf}��M�����GW�?�`�w��A�Q�s	沁�rv���+;d��U5�5�Fz��W�ٟl1���ȭ��m��ܴ�vM���K��9傖�&��|]
�9'K=ӽ�	�Gi�W�ƌ�@�0�5��x�������׎i�㙧:74?ٙI��
ď �8I�-Bx[�4aniB�X�L�*��v-f-�
����=�$�IFYWqC��Q��e�.v���\9�%������ь <�K�����+x�,�<V1
f{(B���c4lZ�������@�"Xf̒�X��ěm<Ԩ)\A;�[�6�g>�?��'�L���(�9F��b@�dd��G�cE{D���Kb��)Vc����>��E޼��_��� �-��z,o����]g�伥��e��&��=�W��Ԃv� �DJo�m)�0>��/�2�����.0�c�;�w�狕��z�ǡ�vή?�ʯ��s���Aɶx���NE5W�+�<-�-��P�s{�Jɒ�%*@����n�+�V�׍��Rqo>��x`�����AF�{R4�G�C{��}~�tU]ŷ�<Iu燆�}Ҏ��C���Doo��w����k�A|"��+�Uz,vT�3�DIA�T�x�6��O�N�#m'�-D�	���H�0�os� ��~̫�W�'QLoe��X��$����4�wx�s��E@>B�!��%�j�#4!��@x��V����V��|g%p#�,|g�
��~$V��h�V��FK��92줮�т�U%�'	���P�_���r�Ǜ�1�[�[g�$E`(��6}�3k�B��n]��Y��v;���9`{�d+|��V��
]�G�D�
�K�������&������=Q��3x��t9�}����
e��T"��7ل0� Gj5��g*0���Q��ӕsz���9�&l������/��CyV^̌���Z��\��_��%���l�|b�,�,���i�:��XV���^UE���P�5���vh��g�p���7?���BS�H���]��+�$t_]q�f �}w�ߧ�i�s!#���m}In��2���'����g1���%q�gc}�Pډ\'�%xl�I���[%hhH�+���&g��(D�֥^{rvZY�A@Q�xڌ�$ށ�Ak���%�S���G���g9��1�����]�<�,�����b����V!FV�T�o�����,u+�+!��!k����Z9�.�����قq!��O�Ϫ�Z��%���l�Q���i�i�?� ��A���	*��H��}�&���gv7"y/�o4����a���b��4ڀ��d�^��{�,�?(3_�|=��KM1K�מ�SR_�8�Wo���6�F��:C4O�z��2��^d��W?Z���	�	�{�/.G�jkNq����7�$��ߛf
%�S(A�Q�vl ����-r�c,��D�|���2��8���D����X��|��_�P>=��TEm�;�1��l�Ɂ��S�4�'����f��0f���Kڣ�<��$��】�+��0��>0I���:�����ҏ��Mfw</��s�&�ɥ���������E*�6GX�#��i>C�����l���4 �?��*}��ߦ?Q�\/EHJ��w��t�|���1��#?���'��P��&dGH�h��6�~4ؔvH�ľa��6�mذs_0גe'�J[ǿ���k7rY	brEkm^�c�X�����T-�;���������J1�J��e��'�2������C�<��xI�H�Z|������'� )�lioF�3��a w�dŷ��$�T<�2��s���;�T@ �W"�K}��Y &:<�F�J�5��DS�g�a�ق(���/.`��	mD�.]Hۮ�n-Sx�%t�{ϐ��zp �(ˬ����������M�=�a��@+ǘ�k3z2�0*�jJl�����<���çX�=���&ŧ8Y���,�@tC�6����c�˱���M|�����~Z��4��JoPM"��7 �O�T���yB�y
N�¨w��#�q�'��
UyC���2�����j�Jf�(���z��>�%����d�<:�\�TR�
��c�^+�6��n���E�����A�Vޙ�T
!������ֳ�؜5ư��P�$�Ce���Y`���P���x�j����8�K�tHh&�����kapɶ��һ����}U���?|ϙ²X�_�w��J+4��f�g1�dV�R߲���WUeA�������L���/Oj���T��[[?,�ebK�8��|����������+Qgl�k���x�슜C R\k�+� cc3M��*��!�٥��u:Ư�VS�F�|��L���}�ӱ;1���͈�& ���s�t�.J
?�L�A�m.Gw	.�qO�'v���[�?H�o�I���^��Aq�b/�9�e�׬i���z>#��zD�'��.ُ1i�o:i=�y]�T�]�g8��T�C�%7x\|A��2�.�Q<{^M�aP��QA^�|�S F"ݵ;]��م&��G�~q�|��QF�.MO�J�mH7ͭu��(�F2���	��
�IjW=����&��	�H�I�G�GK��t���f�ՌW�J�?�1|G��a $�yy�}�>�W�T�/�s�G�e�"E;#@PTz)��2_���r�H1@�7Y�NKW�����y2՛(]H�;�)�6n��v\�� / ���m���}����)^��A�-e!�P=6^�|�mK�̀<6��):!g�N�d��+PUE�@�K�[���@�]~����˰�v� ��gKہU��K\fn�� X{>嗰�r�.z(+y����R��3Bi�n�����=x�"���X�Х�����r�C/��i����z@a����`�y$t���}�e	��vCˊ�
�`��=qK�����]��)j����b�#�X&�k'.L���ta�bZ��i�
���[�z�j���v����:Kk�]x���@eBi߸L�@�� ����g�J�(W�f�7KsK�6z�[��K2�Dn��g�iV4f��cC��z�߃k�J�Q�t��S8��f�v\N#97V����I�Ƥ���z=[�aS��%�Nh����q��yK�Z"{��������v�d'�"̰�^�y�QP'l�K ��+�;����z@�*��d)p�-�&N�m��~|��*{ �&�Nt��>���#9�AP4�ֲ�l�+����i���ls�ٵI$N�҆�L�Q�%�ok��z�bs�f꠩`���Q�槙X�h��K�)�q��6Ϧ�
-y��~Z��k١��$xR4�c�˻��o /��\��3��)\x�6JfӲ��t���hD��<�z�m�z��o��ZI�]��W"3��|�EI��TSx�1_7�� ]��؂J��uCCAI���wFY�x��09�ƒ��N��*��~(�\q��(�m����N~�&����0V2�I�/����]*����:S��I'��x�C�vG�#��x}�P��.>�	�B��� �.�70�N^[U�ğO�@�⻅�z=0p6�����j�2:DG:��hy�@MU�8��eV|۪�QӤ�C�Ƒx��n%�lI,��-,�|�-�}�� )X�U�8���0Q忩��t����5���6׋�*d1�[x����7C���&_�0M� %��#�8QZ���'�L�ٸ��h�f�Ꮸ�?r����s��_���4��̔Dn�l��2B���|�I��]Tp�*��6Ϭg|{�g-q�������7ʶ�_2�<�ͣ�����M��N�/u"�1��J:��s�m	
K�9���`pu�Ⅎr������K�����k�ŧ��@���5�%���'<B�x�@8�S4^k��Q�$ a�Ҹuȡ�8/�w��n&[/�U��>���� �=d�^�-F��d���ѻ|�i�biWg5KsӾ��Mq�ɨq�o5����t���O��L9�P ��Á���3b*S���ig���im�b�|���������]�pՑz[�wh�L��A95m���/��}��g�l�(���j�q��M7�c&���nՓ���u��K�Aj����,�����*�~�|Ͱ;��$�������	�'	^�G�5F)�C��w��Í�L;�Y+G)t�8�o��#�	Z�?ؚ�ZAMe�&ُ����M�aZ�7�� �J.@((Vhx=����$�k���o����JXP� Tnm�~>p���{�3@�̤߈��d�	[��4�8;&{�1[A�
���[2��R*�6�5զB��V�f]���k�'w���mm� �^Y�^^�	�I� ��TJ3@r���f���x�c�\F���������i]�j{+���M�����~]��զ�}�<�~���S�+V^M�m�1�3ʗ�Ĭ��;�Fk�O+�,*�Wg���T�*���������&�w�DS�^���/� 2o�,��� ��{�/���HNNEHP�/V�Y_h#���M!��V�����9��樤5r���~�u��}���8�
9D�&��	��k�X*W1�g.q	�s�&\o]P1I��$Ӹ>h!'QPM�B6V�u玚��7|dH╅k������W�*���A">Z/]���8�R!��DB�*��;h��j���n�!on�wk-�5F�8j�K]�&���z��o�}Y�����=ِ�#��X�gjo�V5��׶{��>�OT�t��ɞ.>h@m���:�hp������T��F�V��i��̛,WdW���_a���N\qŻ�E��^��󕤖���`�ca��ǔH˪5ݰʔ߄~/�4���N�~(:���W�4��ȶ��"��Q!v�*F9�3(c���&��B#�3�� @���x���W�\h@�"R�RQ�:V��ڴ\S�1���(_dU@+0�J�!�}7E����8RJh��]�m�Z��y��xE�ŇHb5T-�rd+��yHQ�����K@�%4Ebr�z�f	S}٠��1G���d�m?��+�"���Bgb\E3u[V�I�o*�ATv)j\����D"œ������'�D��*V���(�HЦE�6&V��W�ݢ�=�(�W���b��!����K�e��r���e���������/��t�ٮ�$����H���,U>��#��V��`�%���u��l���b�z�Á�����n���&(kBY%{�Q�~6�雞�z���X���5��Ey4��@8�\]����b橮x�����1`Sr"�#i��N�P�l?�>�z�4�,
�����m�f�:�ИS7^�mnl�*˂9W�=PH��%qG�y��p\��M������mp~�X`0��=c���v���~�jO�o�H�<+�^�Z��G�ɂ_��ew` �V4}>�B�k�r�e�a���u�_ҁ�˫ڜcS��W���lVin ���jHfM���P��-]PƵ���NibJ�H�d?�O�z�a�J�9zm����ʪ7a��YM��r���*�^�{�M6A$y�Qp��2ｽ�
nҿ��X%�Q.B*�;��g~�I���
��mG�*?���#�g�g�*d���+%)0x���#S#�:�[VsH޺�!q�}|ă��$Tv��$-��Rw�m���N���� ɤ��l���O��	���g�.:VnH� �����/�������L���
e��U�����:(��5M�d�ۉ��m��.��D�.`��1O��>��춻Xl�<� X$Rn�����V��h��^l�Rop�_=`�-1{��i- ���C��=Ԫ ��bz������-8�E�BO%�;�iK�H+�$���li�ɇ�����H�G�&��m�~�VYT�T0
��,���O��'p�JP�s����	�
������+aS�
޶7�P;g��di~q�x"Y$e�����#���i�g=��ӌo~�$��D����T/sY��EAu������*Ds���%&�u�4�8qi��>���1�:�(���\(�cظ| �)K	���==��� ��7 \���3s:�W���$Ԙ
!�sKo/^(g,K?C�Ɍiw\7ӡ�;�u��r����ɴ(��N�����������l�4�&[6�,`��_P�d�����oeX�*^vz�  .Ľە��/���=��s@�i��Y�H�]I�Xk�Jv&�:����z���\�.⫘���ǒ:�ϫ���x��8�#�Z�F�6!yf��'�I��~��o�Q����+Ѭц��y�!�sa�{��"qI��o,�	�	l�Y�d���c�ǿX?��0����Ȱ�c���,�^\���Ή4���E�iW���6@De��Yͨ�z!�m����ܳ��d컥�ATN���9g�*<���]�n2O�$PƔ:i��iFzq+S��?�곈��-�b�b�0VZ�e6K���{��H� 
��D���s��'��T��s ���W��9�
ڡ� L@8��侵��
�y�>K�u������%M�ۀ&�Sz?��Oy�z��x�F����QS�z3薶�	� ÕZ>��*}�'1�5��.�T��vq���d�S�,��C�r�iDzؓ���+m>��'�|�w0�uՋ`�"k��0 �3_��l7^Ri�U���v:��S�o)�ؾ+̌X�?ul���p�Ƥ�pj3�C+�떌�\veAO=ci��\��l�`��h��3�V�ѳ�KԢUʰD����5>��T�'ET-���J�RB�R�{�B��w�R�<��� ���r(͛��44r�p��.1(��&��� �1lA���$�₂��R�'�`n,�D�Q�	u��6"�<�5�B��ya3�����w&�q�V�k	"ա�=�y\��~�	vU�$I33�ވA��k*�=»����x�
���':�b�c�T0��ߤ�Q����=�5L7�{��h�;O9�B>�؀̀էX���,�_kVn:_��m�!�Ls�S��Qy��\�E���)�h#I�y���z-��c�c�E2���(B;�t�(:��V?~dn~�!��WX%OK'��g&��MR��'���P��Ի��mC[¥������1�Δ�Do�o����&>^����.��z�=B2��m��W)b�%ƚ�8n�3��ß��[����@�'	�4�����:HXm�)Íf�ϲ��,�|���c4��X�Q7ܗ*qM� �r�=�/sی���+�ʏ�tQG�= ��a�|��.��r�Ɇ�Sߣɂ�,�=��=��U&�A�m1����7�f��M�g�k��z��[�����Z��`Z6I3c�ؠU��aޝ/v���IL$#��̿}��/R �s}u�����a���ŷ���d5q���Γ@�A���Z�]�@vXA#0��KR�P�$D�	��G�e�	�\a56���lhV�����P���
��8��2?q��3t������
�N�����eU���"�G1;D����/֧�r����tG�lx��{�E�#�;���K�H\�b�Bڡ�o���P5:d|���i\�u�$ax��eq �:Z�H`]�	��0�(��e�=&p3��.�F�*�b�{��TH#خ�)�YW,G?��*&������a�w�μ�8/�շK���b�<%��Hk��O��_N��/��u3�/a���'�e�B~ˮĻ���6�81)v�W�L����OK������m���!ho{	>"�ґp��Jx���\z���"q��
��	��8㎽�f(^h�����۴1�D]����u8*��@�)f�*���`���s��qL���2e�����˧3�x���C��~4R�e^Zѧ�����	�SL���
�T)ڔ�8�Ii���d��ƽ� I��n-W���1���D��zR^��D�kW�Qݳ�kE���@X��������*O�Ф����/z��錉D����B혧�e
e�]:Eێ�E��@=�/��m�gU "�Y_�;��XK�t@d�4�0�Ew�9����#�-�3��W�y�e�{�P{�_��y���^��5�Ql�Bț�O�����X"Le ���!���t �"6�X&w�K�����8
ڵe����RX�N�U����{�R�W�5�>�>�X%p��Ҳ䓉~ <����I2a���K��P����հI�I��I�'A|��?:�Q1�W �ޅ/�Gr,]{�->�c[�Re���j�����	�O+
�vI6���ø���be8�%�*�[u.�C������zp�9�4��~���ᾊx-���fH��]K�Zs�q��܉��k��9�x�"��(���3 k��^ ���y��O�ږ�@K�?x��A��B�y�ӹI:@i�}7'������i�~X��x��@�$�̺�U�NrP���v�е��v���Y�X��(*�2w�6�"���ӯ��;�μ|�	��,�p��t60`���b��R�&�S�Í�JL� 3�%i��bkuF�@�S
�Co]�J��ޏ_���j9��N�Ƶ4�9���1ɹ�k�e�d1�*�tjr���Z���c�c�D�V,B�_wbٴ�(��h���q3e������۷���2mlρ��I��{jL�;�.~�9���쥛:�������N�J ��|3L2�Rf�O�Kn!�x*�%���"��)��`n�&�3���C�J�j�P�����.���w��8"eM1��u[��o�`����
���Р����8�ع?uE��u�!�["���厏�_�*^�(3�[�Y&�>9�$՟O�N^�\~Y�iEΫ-��-�o��v_�D�k�ߤj�,S����q9Q[.d���*��C�b:��O[^�I���5��;��n
G!�]R$#�+�T�!)#�P�K�_>�i���^̜Ϡ����׍| �u�'X_x�]%{�;{we2>���)�_�c&�R��:�Tu�B���*�Uf���&W�B\�f!cF�"��_�<3='$z��v�@�<kN�,)����.l��=�K=��b�t	��
l���X}�>�q�?Y�<����t�	��G뗖�n�ZW:E��7m��W�U�*cy|Cϸ������d�Z��I�-�q)�H��K�T��[�LB���K���82�Uf���o���;%޲��A\��_H��