��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���jl�7�x�֫����_��aoY��?#��#�r�m�"R^F�(hb=��pt$��e[5�v� ��n{L�x����o�x�+@wM�ca冐堏����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A���q�	Oɇr���-"Nlp�-��%D&�\�*O؈j��p^;Ջר��Ƃ�b��![�Thxa]w'�|�#�G�0������fp
�G�9+�H}�$xT.)�P}�u�-t-H��}�c�U�H�#x���7J�E���6GJG��T!G���csp~��"V�:Q��e	�Ʌ����(��-���>hF�/8W��7<xHRwf�Ӷ��#�B�O�l�6�� Τe��}.���M�lF�W���}�ps^�{'�D�.-�r9G���:��
�\���+0�����:rm�no�~>�t<$�a����zs5�RШ�Z.��m{�� =Ge��P�j{�A���ĆS������g㓝�&�FA"��j~x��ӽp*)�:җcC��m�J�Ѷ��n|(v\'��z7����N�Q�@�	��_'pr��ZK��5Cͭ�u1l�՛���T�q�@����,gv��K2x��.�p8��Yi��������X��*���2�}�t\s���ު�>i�7��o����e�µ�i��l��S�$B~iL>C�ck�>C�����ܭ��%���S����LG��}>�-mG㙤s5S]�K�o%�I���W��AQ7.�3���Z*��B�Fq#�g2�m7�?�sLT�~�r�9��U��tϡ�M]�q��o�|j�Q��1��O*��~]OU��ǟ���2����w�J�8CX�����F�R�j��Y���C��X\�p��_��bi?���w��u+N�?4��r�쉴�};�	Ðݍ6Sò^���˔%|8L�ף$��f�Z�i��;B�4]�1+�Tt�Hڔ;�d���.BĊ-�)p!���Ty`���%����i�E{���ɡJ� j�M~�r����{%�3DK�f�	�dF����6�k�EWv=���}�yvp�	�)^č�+�(�����u�,�	���,7��3���qjM���T	��/<Vj�E��)zw��3��$l���[x��zW�0��81��{D/�BV��!�̆c8�s��G��I�'f�Ĵ����bШL|(����V�[�,iYNE �*̵�Kx��M#��:A�{��t~�G~== ��Pر`�.{�t��~�sԧ��9ަ(�_7En�J���g\^Y�ZY�>1B�_>	��qH�����(���G>@�]pgm.�ʾ�6�Y�s�!
Uf�L�{I��*�Kk��P)̓LG^6�!p��#�d��q�7�:�J= �xK�_��q �r�B<#��fR�'}J
�~�r�Vi'R��o����J5��>�
����n��x���p�_�"��ǰ'ܒ gʐ����(�%�,������Rl�թo=/Q�qbY�:�U���u62�����i���y��w��z!�q��ݒ�ܩ� �P%�9�$�����`,����}���1�D��O;�)ױg��cJ��P��Fu�{'(�	����KV����@�A�`�Ǚ^ؼ���Q�:��bX*��U~��W))���(�X� Q�05�Ǆ��^�,��2xD^�o�)�D�6�f�ԯ��B��=���F���@�����CQYfh�����b��cu;�M)�yDlu�P)�'uzG�Mc�����˹���Kn��2�{�J�v#Ҩ*���^��3z�~���v���H��F�ex��^O{sM���G�f���9�%Y9	()�yq�[tx-'G�*�ܱ168�>X�_}��� !���9���siP�] �o%&LϞ�C5Ŝ���^�2`�;4f��-��z�B� wj�W�d�&wt �i�O$&8�*��I{�j��ɨ���$.ˇ�H���`lc�KA��:�����(�m��`��qJ;c�o�1� �R���0*Hd�{ŭ�?��Mn걲� CM�����c�@�d���#�i'Q΂BY1���ӬQ�(�uoL����b��_��s��i�8�*~:o�*._��.��4L����$�J����i<^@� <�yI�tth׫���Ӛ� ���%Z�dس��yL��D��
]�Rq0��T��.�,8������ڰ,F�*�:
�{��V[�@�ۅ� f��+R
�H)��플X�X�$�S:A�ڦ�آ��ǂ�����o�������*ó�F��-��F�֗Ψ�.듿���w8#&���:���K��uׄh`�R��{�c��a�bT�V�����K�h�Lў-B��~*��<��/Wr�iEE�İxe�x1@>|�]|"	(?��!�s]o�(��� �(ܤ���J��뺰՜e]��Ű��&; L�"A� �f	�PŰY�2*#�`��+�ܭ^���4w�'��E��Z��Sج;�o&Ǔ�VbX��cK����΄�hI6>-��ĳr��n�*��n@���зY]	L�	�|��>��h*g�&k-؁k�����ᄽ{�"�d��wo�Hu}�������w�+K��ͩ{��P������t���Y�)���ݐ%��4�Y��5��S��L+���/p���G
�m�X���FR�0��X����F���̶�����A���7����.Z��g��Q7 ���i����LHXn��>���z����6:�X,H���R`���:j�ʦ�D`=�7ż$V���zp0�e��r�(��aX�ܧ�E�c5[V /��Ic���\N�� ١z�	M^��2����G��X*���+k��`X�dz����Έ�{�/�o~8�|o��Q���
V��u�-���Kg�?y�͙�.��Fn��]�s�W!5�Y�`<��w�{�ڦO�V0�;V\�%����,@�H�����4�-��]#
���[Pk6=�x��ھ�k-�#�����bp��ӿ�@��Sqw�9��T��Ӄ��zi�v6�-�;kU�g�s`<�"��,�-P�t�|��0V͉�0:�R뒿��c.� 9)����l�}iNaRC���!����&%�(�)�)HM��͊��-*dS��%	}����*�[ԈcGW�F����"�tG9	
#H,��a� ����e��=��6�#ؿ��9�8��̺�}8��?bϢ k~��朹S�A�LN��I���|��j��t�
�j}��,~A]|ȄWC����N����sǀ�ئM�0�!�'!�W�b�{�U���`-��I��b�;�u*[aC5Fm�D8��]�0JBaM[Ue2H��
$�n��V�B����[j�tEt���!���r~d+h F,欋sSQY�m���*���)X���!�?��g����^F�����^g"��&լos����'�Y�ޢ��|!�l4��o^l����y��K�AG���A%��k��Vn9ϋ�US�V�Fr���u�p7!p�z���K� m�6��A�Y8�6���$��D������~t_[aɽ�{0Am�:���}R�5[�y���V���&})&7&t���=K�A�W]�^z��J��[sJf��[e�Dm�	\�f�?�K�Ga=�<�����|�K�0~���Q���"-�R�����S;e�� #�|	5e����~�7�Yo���/�\����cq[O����{Joy�Ac��/<p��H��mWi!BLW���a�w�M�קa㸌�W͞��G>v1`�b���W{�L�#����&!���f,?�^h-�fF�2�8�����$4!_X��v��0>3.��)-��[�*`���n��\J�pbTg�j�ǉQ��q�%�t����Ph0]�ht�����i��G0���h����c�npn��zE�n+������)���]1�&�ğr`H�|�A���}���w��O�GD���Xܻ����~A�� 9�30Vo�(���?D
�g�D��/�������%bܹ$f�zɔ �x�e�L�<.�s���l�iσ�霙����DJ!6P����y��n>,4l&4�ȧFb?�Ǎ3>#���F�pv=�~�C��ѕ�^�|�Ee6+�P��M���I*2p��PA��w,�0�8���,:&J�� .�y3�p��bx?��S��(�$��I�L�Y�l��gSP>���tW.`��{>ӯ��&��z��6�/ZV�+�^E����8'�K��)N��T]>�j-
���rC{T�������w���㐻�e�<�X��ڍ9G1���J4�>�S�[wL2���Ѻws��3~�X���N�JSQ��4����g��a�>7d���el���2_��!�%pv�����:cƝ��Ѐ_>*���nI��Z��"�zG��]o)v2t��EM�=��hP���E���!@G�h�v�F�:0>:44�1ɝ	�a�Ş�����׀*^3����9J4oqB��w�v������C{C@�xZA}��P�]�#�0��d|�9�=��\*v=�$}k>h]����x6(�x�.�^�y��� �*��q�"�I,{B�>��cA�郓 � �@w�XD�TݍMY�D���B1Ӧ��K�~F�V��K�����Ŋ���X 2꘱T8a�������d��i�09��h���I���ξ Př#'���#`�
7�;(-�?6\[GI����O�ˁQ��;��WA���%�����D!V7٦"�>F<�_"���B��-^=�y�
^t�A��~�TT����0�K1[H;.Y���_����Ľ�N�P:�L�� ����:�K��|�Oy���Y���W�&g}3�}~�zF��A[i�[oTգ��e0.��W̘ZMƺ�<,2�Z �������ܿɢ�]�$mm|8OFv`W|�!�Ay����i]ܝ�}�ܿT��`C0{�or<��"�٭Ky��<�]\�'�B�Mo��I~W�3S��������x0��
o��⾱/�W~���=�j�,��0�	$�۪����҃���%�_s;��Z:Z��G���Q-)f�I<j3�n��aj�cW���S6f�S�xᬨC���
PZ��ޠ;1 �u���������C$	�D�fot
1W���+��(�Zf������/;,���2޴M�O��蜇N]�8��� ���L�w��}ى���#>��m�#*"
�{��������	Xz��혗=��o��$����.F�k�7>��]�'���Zi�=X� �0t���=y`+�F����Y�-
����.� ���l�YI,�˕�����b�7iC��tR:;Xv7��t�!$o�ە���y�=�S��$�Q� �a�� ��e�#m>hs�u�T'��fˋ�������78BR��H�D	? &i���=#%�]܋�4�_�Ljř��&3:�{KOU��B\�+l�C��P癚S���{�!�ʎ�ę�>��vo����|��~���H�ۏtF;G�(���
n��P�x h�[QBJhITi��⾓�E�E����ˍ��������7*�-����Yl�ϐ�@��2w��(��
���P���~Xߙy��E�$�힃���{)^��^]�������s�3���o�6��!����+�~e�'� �x� )v�H]X��4�*� �h�e�����nŢLC���&Z�2<��"S���!��ɇ$�FN�9X��{�H�5w#�v�����$���،��&��;��.�,�".�B�:o�uh�H��"��(  4�Hq���菼����ȑ.=�#�� Ƚ����wo���J�g�W��o$,ܛE#��~e<�-�B�ks������_$�=�TsP��&N�Ӷ;�	��S��5�ZQq�ꢺCGؽ���
��sh^!�CIo�n�E��cH�o�S�ώݲ���x�_�S��d)ʾ��(X9�ŮL@Tw�I�CA|��Ο!�^K6����f޴��d�VD�!�gk��0ˇ���-e������u���8O�;S�p�i`�l��4�v��h���13�)�z��ϳ$K9J�;�Y��n��/]c�Z����G$Bx	� �0����=�$��6��&7a�ΰ���O�ww�j/[X�E?�����d��H����"���}%�v�`/�x�X�!VX�b�Z���л@.�J�@��j���[��ϔ�N�I:�a��/�݃C|܅�v�jC�v@�����A�m�t�+��o��x�����ׅ��^��N��PT<�T=s���)	�~o�E;�^r"n��z�E����x�{�L���n���#	�EZ^C��9^ݘB������6$��3�5{RS u<���&�i��v%_��]�Íd� �S��]���/�Z�M5��HmW�JC�<�i1Tv�:����{��}�oz*�����ΑiF��l�Gо�@sRaT��?�Z)�X]��m��z� ćZ ����:��~Em�n���x /��	�Z)%F�Z�,��U���8+��AK���������a%��Ϲ�d�I�C���z�Χw�&=�sF�|�	���hs�͊0�'�(Gi�Rg��:�a�2 ��6h�w��7Ŋs󽊇V3�S�y8���Hf	�$�t�v��4E�]Ç5�P%�/d*��d�]t�0�+��4�ORTn�T�zy_a�'��-P��)9]w@�K�=�D�R����rX�����wd�K4�ԇO�(.5��m\�L.}{�cx���g����arU��ĸ���g��P�^�:���^�C|;�`p��FQ���B߲��k�)>R��f[�i�&*�|"|T�\�OL;oU0G���}ŭ)`TQ,j�yP]�0t+Z579u�\�����¬fZ�]�L�B1�Jn\�Iٞ��s$vI�g���*��3o�_�C���k�eP7�x��+��%8��RL��e�8`��b�����+H�É�0�\�bm�]JBȏ�T�&+��6{{d;}�
3��ߴ���T"��?*dg�� �Y�e}J�Z�I �U���+�F\�R�����X[=�#&Rޠ�Ǉ�ag'o��jRF��ڜ�Y��2�(TC94Ȓ�^���|���ir�L4&w�=��@8�$;ɛ��xWZv�9���b�P�8
<�����!p"/��e���q�M���h�Y;� ���s�6���B-ٗw��x#����;��f��<]�5��,ԝ��l�����$m��G�$��жO��>z>���]:i��l�u0%�k�a�,.���e�oΟ�0A@����r�荍����9�L���VO@5���;���7ª����g|�K����qQ�,h*)d�/ �l���q�f�"��m��=�R���S�c%�AƸ���E��xg�9�܊n�ax46��{Ї'�w�E��v2��T`�%1{<�us���λk>z�\w�6-ݏ��M�cS��.���w]��oGӠX��H\��W,��+�jÚ)s�G�A����yG���_��i{�{eڬ�,Wi��}���f�0�l��q��9���/���EE�L�hQT ��w �E��.���T��=I���tbs�� �V�dqNp�X����۬S�?��ڪ�ɟUuhA���c�����\{���B.��#�!���M�G���gg��}����L�7�h��ZA��ث� [wDhwd�XhL��8z�����}��wz_�����\%<�P�Ѣ�}��!"@g�"���zP2�_���	����!����.
���]��&sn"���'|�OHZQ4f#�d,���K�
"�t��FN�`�VUP����5�,�.���=9�fcvf�b<�9Sχ7�O�_-=�&���였��*b.��X��VW����kR�%W�Gʞ��K�of8��\>T�}9)i�Ӳh���ҊF�̷a�����r�]�B{�v�a��ڌ�%�����O��L���p%���*�aq��-R�:_�7g���2:5���6jՔ;���I�z��b`CAX0�S o���7���N�U��7��\k6b.��${��U���%�1p{�x��C.OZ�b:׃l�>��q��-a����V���Q'�h����'�
O�vT�aJ5���y��J�E��0��BmP��7a
�j��qU����Lwhko��[�s־5�R��(�vM�?�_�{���O�_�����Ҏ0Ɯ�W�҆p��}-�Q��p>�(��v�F����K?��0õp44��5�ծΞq��/Cc�Y/��NP�uG�߆V:�t��ͫ$7���@��G))�Jc���f?��+ �!0(��Xa��� ejC$N��o�A���폟C�Oe��� B(!�t@�5^�:�i����pFq���po��������Z!�'5��o,��g\�/���~�`�0~k..����\�8&&�r��\Du׃��ѹb��F�U�����4L����F:�|H��ح-��p����=�>\�7���zWr G�W�g�7Э�Xc�\��[���1)��z5����K�HX1m�y{gܡm"��FUa�B�d�sa)H�@���3�4=�5P6;���'J��m&��c'�'}V��� g��n���ע3�9���H��tos�)ao^T8aml�b�'�a�sU}@�4���5'���F74#�9�HA��$��3�N'ޅ8��������z�c���নhS!q\fX��dO�����js�O��NA���bU�_��[k���rU��t�<)�5_g�ƞU�5�q�3��o�la��*=�̯�B�oU�:|��'Ǖ����OQ�A��^D<�t^�-��u�;
U	�L^>��p�!5���u-ߍ,� � >#2"���^@v6p{Q0a�C>��F8:P݀���hl�n���J�=!��� �p�$�oT�%�T/':Jw��7E�6Y�e(�����5b�F��B��[4��b�0�Ø�Ϧ����k��QZ�	5\G�y�Bvl��:Q���G�O��h�����Qi���)k�gt�Y��p�	�`8UoNj�R;���g����K7�%�l��}w�w�2�Co�w�%�;�D7���W��"-w����Y�VL�7�ڧ�C9��F-r^��p�󧰘�K�^�Ζ� Ӫ����ٕI/��
�D��3�%���@p�KͶ�͠��=h��X������ U����A���w���h2.ЦLO&�V��zXϐ���3D��� {jD���3�3�6��}B�'_��e9�N�^ `���)=�3Cѓ�C3�0i�}�jl�����������w�Z�Tύ�Y���2�{v_�pZ�B�L��"�4$���d#P��͇;T����2&�O+ ��([����iJO�F�ߚq�y��BYUM1���T�!J͓ѽK\!!��^G�Q�����R4 N�w׼Vc/R���"s��=����91�zخ�[��7�:�3)����2�:!��E����?��o���.ƼJy9�y.9VI��|H����!^=J+�Y\����r	��)8[1��s��Uk��L�P6xl��u��
��@��D?}�YyLP3�
U��yND�;���oKω]�Z?�ǒ��7�G���&�#|i��M���,�,��gYN�o��lnn [���L3�;����
�햽¹�[���N�/��� jXt�@�q�U��t����$�I&�ۂ~��%9�r��屑����i�g�f<d��n��D�a��_T��0
xZ��Z@�)ƾb�:;��ـrK��O�r�=|x⇍H	/�6�9�yM�9Z������c4P�S��щ��[�#�9�7�T;e����{>�X��u �8�wd�3 ��t<�?��5b�j0C~N۶4��5(�k9"-��p���_Q��:���4ُ�-������Mv��'�cI�]1���,�#�^%Yg�Zmd�M�Ȕ���}��(%�ñe��-/E���3ǰf xO�Q(��޻+�(� �kq�C��
�����%&0h�!���ߤ�R��8�0"̣�"�tɸdx/���i�Wkb�n�i�V��V�3bM�r�=��ury�z�8�M�P����*K�iRp�'^��k��������
k$�%L�ѥ�9ȷ�r&UeY�J�YߵG�Ȳ�0�J�H��ȳk�nN5%�������z����?ͦ�6�eA�*X�os��4������lU#w/���������&�%G��̉��%�%5IC�����1(ӥb:ȥ4!���Q/��� �b�9S971Bts~�\��������-�1b�NBS�]���`	"c���L?DA�g���% �s�>�R�E|�1���h+0O�E�J�Ǚ_M�΍l��Y�h����jO~��ԥ���w��� /ϋ��dF$�{����O�o����N�lX����59��0�O1����=Z�?��=��N��-:��c����V:X@�����k	,��҂��yS�"�#;t�ee�
��&�zVgG&��i`[mg�Vw��#a:�O���u�����a�5y����/_�%[�N�̗}1'�1�d�e�$���q ޑ������C$BZ�gפJ�H�D[��ã?�8��;	��q1s�7:ኂ�[/����C3�r��9(G������j���j��,EDK� UI�D����5���g�v��K�}*ӌ�"lT�昧܋�,��αf�!�sO��E+r��_��{4�جU��^����u��T��T���E���V4ԍI*`�a�]�1y��#b���#Ʀ	��Wy���7�@w���h���GQ��@���ǔV�4�3����M5U���n�Z�4��I�l�,��w�C�(H����X K�Ey[s��@���� �H����e4��ѹ.n��yl��H��_:�Rԯ�{Y��+�Ů��5��Ez���:B'l��ЈH*6�[��5�
�%�8�*���C���-&��;.qF�c o�!i��#4�����A��/�C�0_��V��&�d"^����+���1-8c�2v1���΀�y��\��D�̙ݬ]l����坬���v[�cO��tT�5L��8S��q����Z�J�&���Q[z'�M�բ�P�Dq��Di�}䑘�����q@�u��K ���dwpiLFĠ��i�<�ۈ8��Zb[�����6p��r�{0�1��w�EH1��Aʸ��S,ŐU����,�W����Q����g���FWҏ����%!���1��ǵ�|jdo�G��f����]6��B^E��Pa�	���<#��J�/���R|$�����p52��Lư��[�y�l7�5	�Y��A�~�����.���hPw5�Vz3�d|����/�p涅QN3���K
�8�;�(�"��d4*������QY[h�/��>����!��]�Q�.X�Z+��W��ZA��H�����7���O6<y�&Vw�ζ=
lUh}5��?M��?�k�dP�3b�r��L��!ז�Hw�B��m����Ğ�9K����p��c��0�'�P���V��6?��?:6��v�p-�3�6)p�]snP��I^Y¦	>��Tq`�1]߈�4�G,��w���}�{"�i�2O设���@��-�.GK��޲�Rf�g��f��;Q9{
�l7����p��,g�Oj�R����Yk'��A&�N��-�𽌪Z�e̮_�}���q�@r�w�V6�h�ܿ���t��t:e�{��*)�����8O缁*����6[c�{�p>���|�l���v�ޙ�q�+U��%���Ud�\�7sd%h��v��!7� 5 SGlE�����]��9��=ךl��9p����lϩ���fM��҇8�NoO���y(��RM+���Գ��m��<�����I�h�O'' ��m7�&Ҭ嬐��i����8V�՘�kBۖ��>I�8
�x�@s_��_�^����#V�K@�H���>]�D��	)@#���fZ��s<7���_���;	� ���	���)���y]e��ւ~/9���������n��I�ZW?Ҷ.��W�:x����ܝ_�0����3*���ک�oќ�xEot���y�E=�� I���U�Y0�:gZ&�B��Ӓ���s���p�?�"a�=2����OpU�&����D���%��/�ڠG�k�S 4i���c5G�=|N��"�)>�w)�����ˬy������?��Q+��|���/Y��Q�#k����8�r� �(pE�Weצ�eOO?^�����>�����}��-k7e����vt���I��=
�H�@��W=S��l�x�7خ���c�˷[���/3=Z�2����\�]�4C�u��q-aZ�-��^~�r��'|6�K߀��ֻ;�&x�dj�Obʷ�UE�e5�|�+.�b�O�C/T{.z�u�7�<v�v��ru�ݙU�������H�C��ќD�D�YX�je��?S�-�ٿ��:c�=Ʀ:)�,D�YDxX3R����+@^I cғ�;|무�z_�[!���MH�CL1cۻ7�Ľ*�Y�4�E�3�a�삂�9�5;��ôxé���d�׊r���4�YG�L�P�ƚI7��%q�VCR>�{+7�8<���f��Y�.>�Ʈ)�[d��Iw�0�X8Tù��P�-���7naF�_���������)B���.�v9싼t��ޛ���Fٖoˁp��5�@���"������S��?�OA�A�Ĺ��q�*��v0y&���\������F���.�U�����h�E�;�Q�O��'��S�cѳ���_v	�SxS�e�|<�� ��7��������e��뚤�MB�j�P$�}(#�vއ��ߎ�~g<�������q�,��� ���5���v���h�>>Kҳ���b��ȅ[6|H�ƚ��	��U��S�XK��HK�/ʔ���y��8>�C���cN�o'ݠN��S�k�2�X��ޔ�W���m������ޛ��<h_��K܋b��pd���Q6P����Kל�;��]%͸�:㾚"!|�`��=^T�+>,H7�r�A������z�	I�Η
��%��gW��<*����6-:߈�$���a8��ܧ���*]+���o����n�����~�/cj�6�uͲ��B#>�E����`�
�=�F��7���mlP���5;ӻB�Ũ�f�:�6!�pCH|6����IS����u���gy��÷���d2ںN�]�(~8�Y�wJH����I*��7�á�|N�������p��[����p�{`wo�O_-G���H�}�ѭ��	V�܍�d��h������M�ٳ�ƷП҂�7<�[e���cP���D]}��D%xG=}�[=R�J.9�IQ�[��)��P0�|D���c�,�y{�G��@>j���P�Ć��j�k5�oh�9�l�`�l"��m7~�%��[},��.�c蠓J1�6�ch�r�����.D�$��%MM�mǻ��?��?ג�Pn�m�R�&��v���փ9�W�-�x}�	-�A����~�;v1��p 4������G|�s�+[��o;�O"���I@y=.��}���i�7���HV�ai����-�1v������6r�vqZ��5�Y��(NPY�[G�Br�[#7�Ef�â�γne�Y1�I�c��C���� J�G�Lr�H�Yf�F�hGJ/"���E�'-?ʷ�|����R8W���w~�D�Q��[6Gr���k� {��Z��晅��WA��,��o=��U�e �%3�4��!�]wOTݺ�P�0��)�J1.��BN^8X5�L�y��ʩ�1�$i/��]54p������fQF����| ^J��o�Y:G�=^�((�
DV�D<ݳI�e �1?A��Ie\��Ą�y|�{1���Co�P�t�g^&Cn���9���d�����(`}��I��)�g���n3mO��莜>V�׊hR���{� �z^"$�pɢ����V��m��Ml�J;��,O��3�tV��`vQz�]�?v�
���P|�P��E/~'���-n����~�ۅ��f#�O�e�YޠI2��f������%�J9Dz!�z�/�S����xҩ�nV��JuR��� F�#��c�kT��D�8RZ����Q� G�룏T��L�Y�$�⯬խC�{�Xw�[�|����C?J׊��#����o��l�����9٩"�s�Y9 ׌Bs�";�6�Ƿ�[~K��#�?O�C�X��|p��=�%�D�H?�~5q	MGm|L^Lp��V~9�uD��=ȱrL����Q`��:]qQ\�HM���T����i�ֆ�|`��j;�x��+��QHi�%3�Ep4�c�܌aBA})�S*0��o�f"��X̻�y~���Ih���f*�| �9\ s�O��:)�Ж���ؚ�R�Vq��M�#���'�\)Z.:����p��
����K8S�+PňA�j��� #�2�8"�v[��bܼk,{[�Hi5����]W��>SmV�D;�T>���=oO� 1��yŤ�{�^�}wť��!9��Bd�2�)5�q����s�d�Y-�ˇ ���L�E!�0D���$	<"�	�Ni��y��}�O�f���X��rKٗ���e���=��f@# �%Z�W�y�l�J{a���nK�H�<]��p����,s�p�z�� ý7���+>�:����6s��-q��Z>/�=C�}�ޔ��Ln��t>�C���M�b�Ѻ���J��PC�T���~��lV��� �o�=\�.����BVr��E[�}��Ґͥ�dS�$� F��q�E�7ߞPز��@�R��
'�2��
<uN��v\�������p�w[5h������-U��=��ɍ�V��l�zV�L�5�&h �{/<W6�B,&���1ٰZ����{�j8dT�C����"�m7JC��q�@��%Iͦ<�
��Hfl$ɬJ���gsb&��ޠP�K4�;�U�3���l��^��h��瀫b��'A �� 3�r��'O3,	���߯�vƬ\���8�ZiOl�,��,~����'����Ƹ��G{��,E׆��k��e��ɥcd|Ǧ�o#� ��\�Ӽ$k�?��}vʊa�n��&�)H�,O�i	�?(С�{�D�1�V�)o�c���(�	����RTyW�23��K>k�KS��Z���C��AGfy�V��}�f���Ƃ����I��%GTr�/4s��,�#N(�(�IczΒ�o'�1����9�A=�`]6�^�J�R@j�X��Ua��H���6���nMջh�q�n�,�qu���m�oX�f����	��-��(AWi�l�g8���U��e@���h�ʠDX1&K1H���IJ-�%m�.������Bʿ������m͌��Q�����/b��A-�� ���Ԛ� �l����,�#ha�y)�A��X=aH�f�o�ٷ05�yF����:�n�9�xnS��:�y�ל�3�ޛۡ<�+c�$���1����3J'\�˚�$�Y�ґaÜN��S#��������Cbz�|�dt�e��DA�ae�1C�����Oo�d'��Q��-܄�x"3i
.�q����j���00�:���;�&�L{�
��YƼ֯z����3��4`5ZZh��(��*��������Y��.+:<WP}{~}1�iυO���g/Oz=�4E�SXq��D��.��B��\X%�8���(גqU*���.�^O#��M�6˹����&����Bxr�D����eG�\Dc��Y���C�P�+���½H	��"�g�Ge�@Lz4�0��m�ņq��$a9����c�g_��d�!�r�*T�[�/��3k���ZfL����O>��SK\�e��#E�n(>AX���ځ硅$����9��nR^���*2�.�*P&�U�r�=�>o�W*��K��#;�K7o�_ϝ!�<^+ ���LK4�lB��dr�1�����EA&>�2��t&��	�`��
2e�7Z��a����o�_y��4��@W��<����
?�����/eL��� ��O,$r�#.Z7�(�<��2�?����yЮX��]��?Wr�P�ې�b̺=�+W�Y63����{	�6i��>��Q��������oł#}�l���W-T�c�Q����&"�:*K������4xW.V��k�����P�Y�^��_�t��8�L�nz�$��2��(���p�C+=4f���lJ�S��1�����p��K�s���͜ce�z㢔������2�h�>�5L{+Q�� �KtE�m�ς��O#5nĺm�q�Hl�I#
�T��}��x6��sݛ�1�s���;��/� ��ȸ��``�ٮS����Զ�II�[�x:K�&��m5���c:"��}��v��|�-	Lv䤓�H<��$���h��\�r����wbz
��4�)` Z�ݸ�tCDp��YYKw�4c����/���V����ua<l% ���%�WY�#[��0�\}nYdk�����|��᠐|u��~�#���HTg���J�06oR��G[�����zW��D	��/����{����g�2y�%���ꢟ�Ɉ�<@��� Xg�Y���mdH&��v&qj���u�<���S����Κ$�<U~�(�ْ��HA�3�E�#�۞ȁ�&� �S,���/t��uH��`�)�/�I��U4�:�;gi?��I�bENH����ah)t�?��+��Ȗ���Ws��l�?��8+0��/�����T#zNIʋEz��W���%0^?�}�3�fD��	�@X� ��޳Z0^���kKf4��@s{%�y+������!��T�iL���U|�����+Y)�T�RLӧҎ��M�?ܮ���A^>:9�(�>�c�j#�o�ns�aO�$��7��%�����K���� \_��id�uS���ݰ-�~�_zS�@��'��$jN�A���ʰ�/a�����"(ԁ��1u��>|���q�oc��ES�ӦI���F[��*�&���\���PS1u[̈́;Ym�J��V9=� ��uט<9��V𼒫2]���H.���ʲ�,���!o˖A�z�at?�p�x�U���.���YF�\[<X�D������7=�xr6Txk�������1&��%I)gE�����u�הD��ҽ0&��=	�7���Ss���ߴ(y�ܱ��AM�eC���	��iw�'v�ZP��~-Mdik��ܤ��O�R�~	Ո�-�B�8Kn�K�����M���<O1Uwԛ=\�3Ԙ�Q])��KK��:�i�U6�,�K���1���=�ϥ+ f#"�6�83�1�_�}��W�g[�|�Z{+/�|��+��!�~O*�i�����(u�˼�'-�.+�c�!gE�bĆ�+�7Ms3|O��ǤS�	܍nG�(�����5����
�7�E��0r��"�%���=�ℿÆ�oA��0�W�ȷ�6D!}% 8�x�F7�Di���E�q��ě�d��H��X�����jm����g�ȕ�R��sZ<�g�i�Q�$���p�b~Z�?\n�⮩?�l�@j��D���n>�������GU֍�OE�Y�iA�(�a�&��5EZfá!(#�L:,$F��F6�kՏK��W�~�Y:Wo�Y�b���rP�o�<��`=��L�U�=�wG��Y@����:�&c���dT�P�]&n��V�ܴ񝽣˾׉ߐ�H�F!����I�^$r�&Zy��+|��3*{�Tu+�\L �਒�r|�KC���9|����T��D=M޷@���f�Q� 3R�Z)�|��l�5�� Z��V:*SAhc��|s�&��X�@<� �g@<>}4��b�~�x�9I����{�;b�e�d�\������TU��h���(6�	�h�����biWw}[��SO�x�^�yqw�X)���#[�!?��K#G�-�Ww�=�6Iu/�%����o$�s9�Z��c��l�6�pq��6y�-$�ꐁ z ��8f��viG(ѝ@'´G�z/k�_Q�=n��2���s��h3Zq���@'���]�l�A]NkDg@O൹���w#5.)�[./�K�SV)q7�����{�b�&����d$.��5����Տ�ڊ\m]�n��$�A�P�ɓ����ɴ��`�cr��u\�d�K�Sq��o*J�j�9�)���Jyz��t�2	��7S��O���ʿ���\��/n$�%�\}χGȶ�qp${�����1�Ĵ�Q����8b�5Ȱ��'9s�w��u�5�q{��fd	�7���e�܀
�+H:9Qm|��rw�C����;�h��&�;̗����n�he!g��4�"�'�쩓�5���>;�XL�3� ��+y��_���%�Z��|��~^�3��q7�K���u"�����nt>�vn4�Q�,$�	�Ix��_/?���1N�SZO�X(�\EN���9�L}���S�U��m���w���Y���q�\$?,B��~�jf��R��[',��v]ҧY�=��HF\+C���v*�d�f㐃�
�.^�o�Q�wy��J��<��M8x/+�; ٠��V��V`�hX�M(d��74��n�.�j��]&sL��@e�R$�6�J�âD?�e\T���U5�2��/M
�z�����s�{I��p��1"�*��FgH�))<��n��A��Z�$=���"8kt̃}����9|'��_�]Ҡt������+�;oU�'�I��aS�8Ӯ�8M ��ߋä���h�"6�%�нD�"�:�M�q%[P��"s\�o�EBm׾-~J��;��*c.w��MR+4�cbLC4=�[�S2f�͟���]Sv&���L������S�!�_���(,Oj`Ev:�y�� T���K�AW�;K}h��i��bQ�u0O=�����bK �ɂ�K=��'���~
 ���a&x��A���%|�1�[/c�|gk�ٙ�>���"&�K�ި�� 	
�`���Φ�z<rq~eJ�����[�\C:sX�j�.�~jt��:g�8�'��uV�S�.�2���wT�fX�j��}گb���*x~Mv��Z��Oǧ���9��x=r�-C��Fu���.�e���U�]��W�s`���DElo��e�����L�/�f�w��U��l�~0U��*�/���y�x1�h�:���@�.[	$u���*H�ʄ̒����(�H B������[����Kſ
랇�Z�_'����,A�Iu���V�U 0���`KbLl�ʱ�"�}���O���LO�ZF@��DX�
/+O�^�����:ќ�<Q�9�ֻ<�#;L;�,�=��b�,��~�prO��p1�Gz�� Q���{��Z6/1n���6�ȳ_S�^͒��+Q���]�٢`ӊ���r�Ӭ���;Y��a�o+m��Y�c\����)mh���K�Ef��S��o�L��Е4hZ� .q��u�x��:���*�D�ko�r`�bS��y@���k�S<��N���x�}k�JK{CZ���a�_<�ˁ�7�zl}W���h�D},��)�X$���l���I\AuAd�����욬R����Or<]:��MՎ:�9r�l1�=����7� M�Y�$p D�����K>��XF�<d󲜧��>��Ţ?L�3_ָ��F��%3�&J&e1�=��I��6�	|a������G��Ղa��w���W��00\�x���RL�h�`�ʩϊ_Z��I�Q<���W�s��|��G�>V����^���8x1C���a�u��}p��{}&3a}���*Fꘘװ_�#/n[cӻK+`��.�XsG��~�'���5B�-Z-pqj�Hp�������x)���!׍�C?�߮|Y�S��s��e\C>�郭T�*6�3T!��ۑ�ک.j��ت����&���/e���:�-���6�3��9CO������4�� �+����C,���g���6s��"Gu���`�qS�5���Q� Fn�S�-���a(9�獦�������c�ى �[.��TT�'�6}q=���ȭ�$&�M����ߨ�5�|D���������B�b
ѥ�>�1�V�U�W��2����RE(#���x+����bh�qi�'�頨
��B�DpQ���Z�-2�H��)��e���C}��2���[�4�'���L#��w���"��T��:�qP���F�Q�6w�'E���^��U�~�$e����duqaz����r�Og�h��v��u��J'���EH���!'�2�C$̔���E9�ȥ�~Nk�/��T��6:~���$h#bZ���F�����K�q:u�=6e�'�
�
��d͘���݈�d�_��$>���B��/��+�����(�� $�=U��1�NuX�A(�>�6����@���)&�������J�`<:9 ���d|��K�C
��~,�L�?�ZB8�vf$�������,�K ª�Pt�Aq	O��Ǵ�����?����M0���������u}MrN#�M��u����O����۵{膞��m�/�����d�Ap����@x�Fc�&���P|cݮ�Nhj�I���eU�h���'�-&�Z�H=�G���p&�^��9�,������Ġ�0�l��Sx��Ufw!Y���zb��
��������N���=y�!�q;9<�O��-��ө����K�{O�K��B�򄳘�J/���!���_R�EP����F�Ķq�Y��Ê!b��7��;+�Vj�Uڕ�|(Gu���J�=�ڲ\�賷������ &��o$@�aw�\|8�hq�)��fE���V�'7a��=�u�mn�
w{M�sAO��wzmǣ����0NF��e�<{��	P��AVԪEg�P����H�_���`[��? �PѩL��4JRv�i�	t���vE�+�ʌ��$����e�w���yx�k�e�����* ��Kt����ۭ_�6�6� ��B��2]Zֽ�{�"���:���/
[�ϖDeVވ�Z��FTK�X��p�8!��vb�	�A+�@�T�qR�7&�#9�z���*>�3"���H* ��Ґ���K�E���]F׼�5���������
����Iz�%R��Qn�<����j:�b���8@cHU�八n��?h�f����uV�o���m�n-�cp�
��-���1����F7�-B׋ZJ��oS���UW[�/5K٩
n({2�t ��w�2Dz'� ���1���?�����IA�^��#fY_c��~�{T�z���k��D8�ٵ��h>�k����9b�&I�F��눕�P�[I���" l�VR�B�i��TD��eH�y��E_��3��lT>h79*[�7�۔%-_�~�T�#�i���R5�ո�?��~�7��ןul�\'��x�'��S��:G�&@�ז�@�j[�0����Qɦ�j�C�j�O ����7],/�����g�z��Nլ����<3*7�R�%c�ӸZ�kF`���Z\�;kTs�����V
M�o�����GQ�ӑ���Y��&6����Ű�k��0�Лo�W�D�X^�_��OW6��������H��v�(0����n��㕫̷0�KZE��k�/>�?� ��t^u�a�v���8�:�dh�����!�q{�1�c�E��Su�|�W-@SMx�4��٧@�D�T��]&��B��ݵ_{�ʇyK5��$���յ�mL~��}�^���J¥�u5��M��a""r���ת� X��M O������i�k�t^���ߑ��^pP=�p��:���f�R�.iL�@E�&<9x�Ͼ�6���� ��c����>eAJ��e��pR&�xc2�O�;����p�!j���"�ЎIt������;;L��+��N��������}������ƕ�p����#j��yd�k
�?]r�'{�l���J������e1��!2�L:��o}$�n{�SY�_�|��_ϕ�R�ɤx�����F�����*T���s��,Zl��W�|B���T2@p�1�LW��5�҃���]�|�/��BZ���3R������"�1�AP�?��/4֬请2G�r�?�E$�j�1v!+!�$6�H�J̉�T��T3!��J�M5���K�>�|+�K��- ����[�����w�F;�Z��*�xq�W�e�9I$��<�ګ�MT���\0���!v��g��BZ�Q�38����`l���{6��¿~}�r�0ԅ��NiGx}������A��6�F�ެ'o�Ď��I�R!��FŬ�{>������0��_��x�N�[�/{~ "1�����@߳���O\��[�&U�Vfn>��uv��hK�6��2OjBB����"c��o���N#�5���8K�h
𸥛�pZʛ�L����d�7�cZ�f��Q��-ULç��TD�>"�)4lD����g�X���`�	�g}a5�!�H���;w&y��{����Lh6�O��E{罈`�8�vD_�3����j,���"็�3S)���9Do-��Q|�V�u�}=��~f
��Y�\�b`��ɶ���<��U���R�L��a�1��>�*�d�Od�[~�r���� ��0����d��C2����j��D�f{�Lp}����,��d�}���~D��	r#F�
Ϯ��J_��Cg.�x�^�K'��7��/��dU���K�L�d�(Փ�[���I�P�uJ�����(Gt:x甪�j�葪%���:���KJ�ռH��_C�-z���o~���l��Ww��%M�;����T��;3���}�o��7�ݶM�C�*�L�p0-?<���{�xCͷr�;�cߎoڌ�m�&�ȫ�z2�)#�/	��W�F%.��ӝ'���hM�rd뇥|�z�jʎ������2�����ȝ-�k�5e�g^��_��S5��\��f�F�i0� ߷���� ü�#p�����>��lo���2�k
�h�㶙a�rY��x"Ov����ڸ�d���<�k�[�h@^�ݮ˩I%���tUs��M,J��B<�H�� �J�@#f �w���M�_��ߴg�*������aƩ6D��Ŭ��(9�+����e~���mX@�x�N��b�4����r&kK�&u�?��i��S��6����u�J�����<1M}��������G�����c�d;&|j ���/���P���*ُps�u{q���v�i}���k&L�P?��FǬe�1{D�3��)'�Sh%U�qj�0ǣ�o=�A3;��g=�g=�ү���q�����x��1��Uv	�8_�+��󊮋�.XALzė��}����u����k����H�)�b� �4dp��2�C+��M�1�18z��fO���B#�*�l���ըӰ>c�@�4���\5`Y�"K�}fa�3*Q �ƶ�T��"j�����.ш�E�5a�D�@ڃ���9F��.�"�63��f��6�4
���P��;� �E�������V�$a�_��.�e��%�;%ңpV��%EcXF�����O8���߬�����f�r�ʐ�|Ѕ��l�;�|A���q�;�E��V�Y���aX=;/j�v�Nx[��S�h�)�h^/�F���[��>b��:V�P&�^p3aBM]��d�ytg4��%�L,s�� o�6PȐ�9%�ַJc!��,oؽW� l*L��r/'���`x4�NA������h�{�
TGw�<�O6�8���<��2��j�k\��e����I�\ ��MUS���;�JQԶ3A�.4�@��vEe��?}�D�%fK���d�b���n�o�Үyi�q�2\���j�^�!2l:��Kwߜ�B�K�)��m���M�ms�K��a�A��>S�v:R��q$R~ZZ�v(`�aҤY��ՑQ�EF������������w�����7&"-Ϟ~a��y�݆�%�sT#��@7Ǡ-	@�QS��0�K��CK�#�)9���B�zK��I�Xa����!Զ�\�>R�9AÜD�%�?��Ik��oWx͢�3,��@�D��wp���p�DBJ
�!�5�$u��:4C�K�C�t;exY%;�)�*�J��*�(�L��؏E�Ktq�9�n��D���W݀�Ę�
���K+��q0ݯ���<��CS�M�Rj�j´�@�¹ͯ��t�nM�����V[lO�*�$O�*2��֊ݪ�,��5$��F�-=c����J�tLD�Q8�B����i#�<����
�qߚ�zU{g$^��h4t���������;�u7'��2,���D{Q�T�� �D�4��"�zn���tX}`g)��τO�pi���y]@�����ow�>(�m�#�`��c�d�s�h�UI���=8g�Ry*}H3ox5|B<a�5�7�����|�	N�C��i��6��,"����p�R*bQ=�)��U	�wiy���j�^�v��cD�ԭ����E�t���'���rq � ��'}LӀ����\K@�>(���o� ؉5�
���@��OL��{|>����R���f���1���MLQ�#v����k��	�0��Hx�2�3�1�NT�m�2���
h?�k�"����p)R˨�eB��u���-��i1p(Wڣ$�A��n�Z~�@��0Hb���C�x*H����U��|n0��~5u� {��**M�ޕ��Ӭ]����Y�!�9t���]fL'�=Y"��z�;��B{��Q�+�E7�XQ��ط"I�O�FV��	�VQ=W����R�SP0��g_�vsܤ|̹H��/�?b�1�2��_�ї��ˤ�'l�ʕoF����r�,�HD/ğ��4[\�&5��e-I��sQj@xC�ӂ��,6��UX��&*_ 녡��[v�>����>���>A���P�:Ԛ�S�� z��lҊC(:����v���)�,��?�p���U��pO�g�]κ�*nNۢ��U���Ny���ɖ�m�&x����(�����,o�i=/����+���QH��M���pW��Z��l_��T�晸_uM�xrE���\��r���i�J�Ǭ�{z?`ÄqoF�8p"ӻdL�&���⋽���h�?��5q��rz��R�Å��7�?3����1�.�nN�a奢vӥ�K)kX|� �UT��~��Z�1��/��'T5�,�j��`౞������b�'c�o��Miݓ��!۔)�#9$(�o���o�AQ�݇ѢüvwĴ�:2��-�?K��O�ÝP>�6����=��<���E�Fw0<�?I2@T� �!��v9�۫.ʂ�#�~ӇnO�d[�r��G�"��`���;��k�>��k�JO�`H��B�=�8�/-f/��Vr����^;.:q��ex��ѩ��_��n�KY(٤D�" 떅}�xx�b�����#W�h��?�Ǯ�YFX|�[j�ق+R�wx�fYfbt�wH��)�{%�Y���W�N� �n�Z}��_i�~ҟܐ7�7��G7�s��M��p%,I�0������6�|�$ sj��I'驎}�;r)������O��P,n�X;*LŌy���k�{BD��N>�O<n�jO����8=ڤ_w���xR��>�s͌�����@��MͻUk�+h@v]8ߋ]L���%���Or�bG(7����did �t�h��i��݊��%�u|��ZdN@������P�_w��k����Q�0TV�pB���ˀ62������܅	�/;��v�����?�l���Z���j/0����Orh!K���
�DS��O��������Q(�B��:�����V�q�S@u0�A�K�2G��[G�W7�&�x�c;aHTl{E!�֎C�_�#+�~��;]z�@�N#s�����.@Hl�y�N�qYL�9����#�G�ir=�M�7;k��u��	z�����H�"���wTJS�)��t�eRu��|�N����kQۡ�c{�$a�	��==��⮒h�=9M����8�6��o�p�65c�,6�h.Ԣ(G
}	�g�	��.*��*���SLlm��B؜�IY0�&���g��6[R�c����Ex-��p+ްU�<���j
���hl�o�9 l�:&��
�?��cN�^�ޣ�o�0�)�Ɓ����P3�<wߞNw��c���[%XRؼ��y�\F\�0�H>�9����c�k�B)�n��\�7����8�� 
�ų�/0�Ƚd���X��'�JF�Kʢz�u=��ϭ���].�7�s�D���ܼT�CD�a��=�ߗ���L�'�6����<g�� Rg:�8�q��)E����@���=:�5ꭸ1T��#2�TO�T*� ٦0P�V�^��@��ra���{'+ X�|:��~�ڀ��dY���6>���/&�)������R����R���^v���>��Duo�%a�[F����jxK�g�Y��ē����c�S�Ļ\k<̮�Q�k���ѣ�{�Ǵ���� ��D~)�4ݪ����a��(�+a܎9�P��gZ�K�� jGw��t����K6��{/�	w��L_y8�����/>ְ)��6�r�v�+.6k��H�ղ�t���L5ƑЀN���1��� ئ�[h��}	^��9�D����[j���)��k�Ɵ"&�F'�`��Ý�R̖K��N�
I˪G'�Å�g����2�-;N��j��ޡ!"Áq1�t�U��i�'d�-�:�T���t�B���-�p{���,���dJ�U!�.kx��4X�;�����ӿ�(T4���FΙ9�7h'�P-f0A|��}�>�&����,�p|b�����==˧u��u��=�����UT/N�]�M�!XF=gC'#� g�u����m���ן�+���_�U3&A��(44���*��ʘ=bǬ�Qֲ�����uy{����i]
�����H�¸�7X��t��'j�v$X��߷��n�s'˶A,�/mW4<!f,܂�`�Q��g��M���_�̮��rK�SƵ��^�3�foZz�1aVD�S��3{�L�5��������q�E��d�e��cYе�C9�K�1}�'.���_���t^4�T��d�W8N(��5�!��|L��_���F�XQ�^�Ο�t|VD
:�V2�c�ׯ
~;<9�<���5t�p9�K�����(Ա5&�f00q�5�,��8~5�>��\�M�α�?��j�$��{������u���L�wt	*T��L��5���FWv�/�5:�P*������Iy��'��n0H7��HwW!ᦟ�K2j|��^e�H���"(�>�a�D�+N�$<���>ࣺE��x����a�DgY}���M�3�B��	�&@�t�:f��U��`��@�F����^$��T�\���1�8A��N^S��,�k�X 4׺k/B�.	���4>b�-A�����.�p��i����*OkޡVj���|��,�ה}���}2X.b�_!F��?�+f���n�Yɂ�Yo
=�܁Q,5�q��R:�;�_i�ʎ��1Y6������
o,��8�H��=� �h��eqنʕniX||�4_n����e���#��D�͛`����zPA��������W�S!������/-���"��%&�S9ٯ"�����]�g�0�[n�|�� $C���?de�����c��*��]�ꗻ��`�����[#GFKH���X�@�����H���9}�h��Ծ;��2�G���w��e<�+4_8�'� �����	#�`�@���:���MH�~��������m� �S��x,Q��]e�p!����K����*�o2L��ೃK�'�K\Կ�b��,����M5����2���<��b�Bh��=W����`iŘ(��|��Kȉ�|��鰦ϼ8�(��;�Ӌ�)���:�����hшж�aM��)K��"���/k�_���&�/�2A�]>����fu�d����+�짻,E�诡 ;� Ї��@KN�z���H�rǍ�敇��R�zCt_�ꪂ�DW�~�D±��$�����J���eKe�cX�w6����t���5��$��g�E�:�{=@ aa�o����qQ�wը6�.Nd�o�ccV��k|��6
�dB�/s�ՀɎ;��J��� �k��'~)��9�,4��4�(b~%��R�ұ���d4a���1H�p-q]�m��q�@V`���"o��S��Ok��T�˰���.ڮ�Hb��fl�>Pqj764n�c]�>SS�1�F�������A*���T���w�;�11k!��w�*G7�K|K�	!�ޠ|a4��-��5s���Q���Kx#��8>�#C�� 7�z�7�F
h�)��]��Y�L�g^���OrQ��]�Q(�/�`�q�<����?s��ڝm�TW�s��k�T�\7�����f��.v��y:=3H���x��b��������3�DYP�9_���U���T jn�J9e�}f �R�d�a��p��Fn��w�#q��cP��3��v���Ӫ����CX.6�s�a���ED_�s�������̾$X!t�l�����1r�o��v���u~�c���W\Ų���؇��Zx�"ʹ/ʭx�,g�Z��f��b����7B
v:52|��s=�;�]�0;	UX^�u��l�>O8��m�/qRj��<�͋�����k��9_(�#~���
�a���fuFrI��ID�R�x&��7\�bDz�S}E�ۈ~���Ұ�6�i�����'��^Qˋ�,�	j�EҤh�:}�zPE��7� �i7�ҮMR�v��_]�f>�%�9YUiA͊.[�J�&4�Fh6F�LA�$��l�
$3��h̞T5�r�J.�?��:�F@U�xVgK�q��P���3���qC�K��ߦM�hi��-:8���>� h]k�L�����Wڙ��+6��q=�������N���']��n�	�Ɨ̋����U\^��Ȳ�-��5���[2IQ�mK��T���X?��	��h�ѥ����J�폿J��i#!0�G� +�����&�s �I�c"��`�C�~f�Ӿ'��B���-�v+�8�$���O�V\��}�c>�xՀ���a��m���a�So�oC�5���ŝ�ȹ_0Ͼ.��x�d-��Р�4raX&Os�O���vg ��{�����E�L&�dp5k�TZz^ �?���J�Ժ"Z���ƟHEQD�v���@,��2�.�<�`m��+ފ�2�Ԝp���ц3϶[2��d��gE�H֢O�`������+p�cm���{���6X���F�}��t��Kۤ�,+A&&��6�����]9��sl�Y����/�fXW�r��v��9�'g.u�Y��&7���?�'^r�a�ECA-����l �>�Y�*L��
�Q�!��n��|C��(� �t$Qa����\W"Emhj�B���6�����@W�dF��JY���a�{U�r~��΅�$[kb�"���.��v��� �u���Ф_�0A}�AIQ\�Da��3�j߿��fH�,���%��.C}-���G}��Xw������/��Jr"�B��Έ�v면�6-���VuٙDR�`F�[���J�f�ag�R�w��D���AiW����)�^�8��Sk9�^]���Aj�k�O���+|���	��oB���b�ɯ�^��n�l�̏}�:4�i�����l�w�;�D��ѝ݅̎Vk*�M���F|4���kj�3�:�:�LIVH����LM}�YX����j�2ܓ��	����aߍp8خrV�eW����8�!���.α�&,�S��c�8�f���mBbA���`:�F��'������";`����R �5�8����j�x'H��z�t\�[���Z�ؗ阺��lo\>��g�"�7�92Ytc^<��X�.��>��Ut�\�+��C^��#k�U7ť!:��,י����ڧ��2W�\ �]����Ah�B�e�d`	��K��Y��k�E��C�w3��|���{JW�9�+�1LN���(�J�� ����i��}��^�H����9ǨN&4���~���5
����X,�_3LIS���؁�X���$QȦ��vAS�a�6�݉Lh�8�[�IE��8�TR��
&iL�A�E��z�e����CY���y��L�2h���*"Rq݃%d/C�0�D�11�6}�,f#�c�/�B���?�����k\f����%�,��Ku����s�hDUg@.�|��(k������vyS�����!&�e�}s�&�Z�T�޷`�����w��B�]lk���>�7j?_�x
_xEj7UM��Fv�^cf�&�r�X){�rSG��z��_�e���-R�d���3�\���d)[~h�*��E�?f��iOM��4��!&���nk�����@��Дw5����gg�P~�GA�O�'I�T!/��6����:/��-�ۏp1!�I0������� 0k�*�������z�G^̓�߱��e�)�:�V���U��X;S��	h��U��	YWs"=C��N�:N3����$�N8�1��a�D����3A� �lF��t�FH���I��0:5r�c�[�kY'G�,��(ѣ���$��sv� �慓;�SO�XH+Á���dՊ�U�6����bY��[OF Yqw[�}X��1�5X����W���h��Y�4x����@�3���$MF��N����_Va{��&��i�uo�|�%~2c�lw�2���=Y[��<^+�0X��؄��ue�CQx�ot/h�Ǝ$J-:9Ap^�q6�_�z�XS�]�1�Wb��F����2Z.<���ԎÓ��/6m-P��h�&*E0f�-1������a��Y��z�A�f����7|�C�NQ���2����@3�HY�E6RM,;���g(�MP0$j ��:������7�F
�l�l���ƫW�V$q��h?�א�%�+��[}I�ǵ����N$i���MZ%���N��� k� �-JR��3�Y���󥵃s� �TN���uZ���e����Ato�7���5�lj�Q9(:cK���wA��]n��G���`�_��r�:C�8:mX��e��\�P�g���� ����rk���%0�=0�c���	�0u&&��%[V$?���8c�ęm��������C[i�g��Z�6�� ��$�~���V��~:��Φ�Z3��)��������Mŀ֢̃�5�9
���;r��I\��TYK&�
=�pAȭ�0�q�o�)��܉���Y\D>���+&�����wr�Po�M+@��| 59]�i��]P0�$�7pE���&ɦ��&5Ě���D&��08 ^��bFVӡ�UNBЫj���ݺʋ�0����uS������b�c!Q�k+�U95�܋oj��$��MMJu��b"���p���a8����FM.4�:+����ђ1=N�5v7��̹:�~ψ�ک���] ��񒆬��!BR���)���L��+]���D�c+c9-C�`��l�p�n�F,��*��#�1V^��<\�����&���ʼbֆc��K�����+2�@�a!P�"M~��X�6�}�N��Dw�2uȘĬih)��D�61ǂ>��%w��� P�%���,���Ά�)�/�-�AQ2�K�0d����WsI��Sռ�U�|_8&���o�E��m1>�Y"�hT�j�4�-D����&����T�b�7%bj90G5���R1���aQ0 ��%�Mh�X�z����E�`��S��d,�/�y@\�Y�/��=�yH:�� �.��֔$��]���)�'��8���[��
�
�H���F8���:��u;m#��MM����a��f����m�w��]ƚ!��h�g���ۺ��ײ.#X�v�c��#��s�ǘ�ʙ��\�/b\�@�v��([d���|��	л�lO��������y����[�c}�	���k�!�Գ���}3�MZS��/H��o��||���Cަ־ R��-�����l�{�[�$���e�O�t\�7��HV��r�V�g�3Y�����B߱�xOQ� ��2�O�׭��i�W��X�~�funY'�����B�F'v�~�����و1��̓0���\��_4��=1?|�>,�nd0�i�Ss�n=,x��G�JᲙ�I�_�2HC�|%�ݮ~r��'r"/�q6�W��]���Yf��蘯ʒW�Ǭ�W3pҔt�Eec�#pYV��y��S�>��AlpKuW��$o���q��Q�pYG"�j�,�R��XP���b��Τ��DD7f[��'�.�6>������f�l����w�畩�R��%���LH+�zrOx��!��-�;)a�=%k�,�f��O)�RW�����R+��w:�t��«���ݦ��?���E�V��z��
l��OGM��@�����SŲ1^�L�2qͅj@
D����
���f{xAʆ��kk�2�ULs�=��@X9�#�\��t��rI�AE���	�پ��˃�Yм<-6�P�xu ����#摈�K����Ǒ��v`��!3h��w����z�`RH�'��7���Z�F\01;��v~
?IN	~�S$�	�=9��l��Wj';��%ݕ:��1�&ry%�@�aW��v.?]�]~qf��9BW��F�D�M��U�}�a�gތ��~4��� ;{��\�e���ؠ���F�����Q� $��o'	�çz)����>.�^M���Dn���2�Wz�$�W).�l�>��5��:�0��b�M����ȁ�T�F��Ń��~җ&5�y"V�E����\+��f�}B�K�z|�<AG�i�*-�:��Ŏ������abXT�!�	���j�ه�!���2�1�A���7��$A�2��;Bm�� =�b�_���S%H��^Y$ޢ/T��|�,k|��3a��`� ��V�{���b��S�1s)�nAe�
����K^%Y���p�����뉸G�4��~W�����kۍ��K�-H�O7�6=O���
�2���Y�!�U���9Ӟ��?��BOf��
�
<P�p��a"+�k��e�i��M����4�ȋ�
� �8:�ng,"H�Y��ǡr�d��r�=�?Xe�"��YX�����ـ��ǼJ����0D����*?B%���,z3[d.P}j������f�a �%`Q{+)�n�:�ʨ�%*�}���f��J�s��x�Wf1���~Sӂ�0yj���K7c�K��X��z�K�oCh<�J��D�I�V
�蒽Hԍ���)�P�(E�s�5�%�V�yb槫��f�f),�.�(�*�g�W; �1����R��Ȯgϒ;>��������b~���85(�k��SFe��0��擐'4�W���r�r�M��T�i�驻��}i�?=@l����w�nz����}�F�jJBB{Y�ݟJ�h��V���}?��V���9�ݕ7�Hh%8�B}e�u��vY t��%�klA���ڏ��p��R09��S2�~�)�B6u,řr�OFg��و�y7�;!@/�*q�ړ��/�{�\���.۠Pς��c���-��8-m�~��*l��7FΔ��^~T1�W��<�!����"dc��c�N�JO�:�1�>4�A�w=����L��O�s��9��Σ��Ɩ�ߦ��©V(��>|�q�fEl�nnF�+�HT��'���4��5��{M?S�4;[ǁ�� R Di�*���8�U�2�jE�XIU\Ɣ��Ԗțt?eغL"O{I�
f��Uo���%��Pg. ��R �L*~U;��<�%�����W�������RF��@1_�� �����9W�6�uCU@�oפN|�:e���U����z��)��Qg~_�p�+��H���1ϭ�iy]4�AIS��9�I�;�������k4���i��2%����㱓���	�]%�@�\�����7��Y���_h�ډGWR�x6�f.�!�əi���8'3��m {x��q��wO�31j�:
�,�0#�/�ED��/��I���(�4qb3`�ĲO������u3���)Q��ܗM�)�Vz�VK���<'�ݖ��O�q�����	Չ�	�'XWf�*ɝ�A�E
V�!���)���sB�`�=4ᇢ�W�P]�-tA�֜��TjUb[;�i'=Jf�Ǒ�M��O�Թ-�Y>�!2،���J��V�Ʋ��Yu�r� �v��!�sSo̓ձ���8�ݺ�'�Y��Z~�L�X�`#F�D����g���ˍ����iƾK�By�H@�����:�Xt�W��U=��W�4���ES��FxhJ4�!�>��dmj?��9���k��,d�����V�0��B7�y��bOb���I���~��;�(�H��B����e��\��u��qw҄5۰g~����m�u�2�QO�y:�?I(��߮#qC��1DƯ3I�a���Q���-��O
�X5���˹�1qu�ŝk�C�ka��D��KU�S�w�m���ݐtJ��N����Ͼd��ɏU Y�1״��ޖA�w+�9��߁�}^�C�P�\:�jE�G]3ʢ�ϑA���3�&�37�2$�w7x�H?�n5���p�=o��||�=yC2��3�wE|��ط@
�)]⫽#���!��7��ܚ�Q��a�h�\�Yc���_���K;���8��6\i�%���wxi�c6w�&�}j��g8n���	�`���J���pq�ij��[m08� `m�P}+��
PJr_,�MH"	_Q��HL@Y�Og5�`�iX�fA#�ݤu�Q��T�*J΃Q���҃_�F���ŤT6��[�7�@J��!�����Yd0�$�0I��JE�lHF=wr����S����4�+���0�^���dhrw�`��C�㍂>�DF�C�Ѫm/c��V��z>ߢ�F��%72ڢĮaPPN8+z+����4��J�m�6�B�d'�wy��<	��ƛ���e�u��
ZQ�3�@l��meRE��Y؟���Fy�?!I��y;�jE��I.@�{���r�v͈*��nUbX���I?�M��0��k�J��){�V|���n�Wi-���zJv`��{�a��u��~d�lCk��t�o��m�k!?q���Sҏ�F��y!�D��	��9����|�/Hb�b�[QX��>���[�?�P�׻_��=�hhY%2�q�0е#�K�����I�X���W�h��wX��v��h��Oכ��voR�����<���W����Ql��:�ÿ�3�ld�ɉ6���#�L
�q����xc�	�X2�����Ue�78U>�](�EP+P�ᛞ��'�2S$����2rp3˿+4	�Pc }7���i�=���l��04�VԺ\����>���nj$�k��d��e'�-a����bNT#e�X�L��;�k�Çr\Ffw��͢���l��$��X���4Ƌ�a53����=�h1����[U�ͨ�����g�&z5u	ذKo�e$��U��-��V}�Y�ulg�e��~0�w��_y���q��6�<4������+���.n�X���	؀�_C3�1��Yӽ��?�t�e�-��Wo��jrZVP��9��^����]�B����)0H��Hc&�O_�K�F�Bz3hq4��d ��Y�m2(%���l�
�irSmx�7Jlz��G�����_���q�~�aOs�j���:R<�)
�n�%Hz���xZ94�"N�������a%�-���.�'�^���_�W�������:�w��8�k�N��|�����X!��Q��!H�֍����	"��B6r���HY�OO:<�4D�e(����A�C�0�'����X��
0}b�&��z㶎�-�?���J9쓖�-�R���k�݄����ȃ�i��8�[��F�~�H=ޯ_��Ld��<�3�J�=�P�dT%O���(�˱r~��X��;��Y��̀�yn���c�im��0��9���j�-p���/��X�k�~&�Cv��V���=r�%ܷH(�(5C}mv3M���M��lV��|Ԯ��E[Q����;T6}���6Utz�Z�}
j��
�a�۟�/���c��D]�5Q��y�0n�_���YU�h��^��Y��8@"Ǖ�J�	�{Ջ�����}��U�ʉ��-&!|����3���r]sP)Kz��]#=v�R}�0��NQ;�ד/ym����Ku���������`z���A�ќ�,)O�UXu��6!�,|7L�w.��\,��F5�5ñ���[Z�e���+�H�ң�q��c�a~�Df��L���kuf���oD�Û�{�=*�Ќ-��ErA��\�&��aD���$��V���Ft�)t��HE�<bX\�����q�8+��3�(Pӳ!\�*��/1��.���M��xWB��-TQ��M��s7�5&x�L��5,|l8I�~������=�Ze�!	����O�N�J$Q]DMM����kHQ@��$%L��#���A| �ĵJ\�0�����\�Q�P�C���19Q��g�O(���G8��HO�C��/� ��당�JL����� ��%�*����KN�4�h������{q��,	q���.޾jr���)�a3�&�K|�-+�)��nܕ�}�&�-Z8虰� {�|Ջ�� �J��9ixD����A�`�GK�0�Mۆ=�U[����}�0��L򬾌3d�8[j�s��ȏ\�/�7�G��N&0K�౛|��s\`F"J��`���%bw+��$�=̢֣��9V,��!^%=���,H7�$�?d�kSH���p*\n�<"^<�M���qiNO�]L��	��?���@l��1��o�u�� '̦�����C'x��Q���l��8-@.��!��9K�4Sm͊�s��(I.NYs	�%�¿"8��5��c�����B|ŕ�j�p �Z�.�c�x#�E��ş�d�K�	o��`���v�<!댈����b�pF�H����|`/�\��Cָ9���1�/J'�Z�W/G��J��רoD�of�V��}��?<�P�Q�Ǜ���R�s�$U-����]��#���z�K^��Ǹ�_=�P�>�ۀ��z�Y$�\�q��O޸��5���6Ch�H���^�#�]�Y��c��7�>��W�W
����8GK�E �cT[����HtB��k�*k͊٦���;W����"t�U"GYԨ�wn������pI���p�7l���X����R=L�'�������m:E�$�7,�a��a�+�[��Ӏ��yd�Fl4:aD���'���e���H�w��-F)�S�z��z��|5���ۀ����P& ~0?�c6����%Q��t܋a���m�����7�lZW�{�1�(xkZD,�>���&a(�P������v���m;k�3z.�?��a��҆V�Xg��RF�����
���ԷC��Ԭ�U�xhE�7+<�m��cz�������s=]4DJW}��H�*���l����&� @���e"±��E���}P���<?�_[��|K���jJ^(Sf�(C$b,�Ύ����"@�=x�
4�3P���Ӽ��Q_�w�A9�w�[V��~�p�LE���~�ŎE��fa@��J�N�=��W�_�f�$gץX��jd�W�{�rJ��Q����	p
�c���%�Y�����b�i87M���.�m��}NS������:��{���I(��N�Xg�=��ٕ�M%��� �o:��nO�AK�>�{]L˖� �,�}P�d9\BU���6>��k@Bs�S'f�;)�{��:�O��B&`��1��	�����mc�]����y�����`��/:WOd5�UX':�e�4������%��;�"������7(��|LŮt!r��^
LU�ކ�E����"�(���xV._�b��ۥ4�cz��*�43����eSnz�R%���V��(�i�I��f�5>����CŐ�i頶x-"n�L֙��;���f�䎱�wV뱌h�ZP�%:1�H���ԥH�����Spތ]`#�!�t-ݙ8H�_��(�P�I!3{+5�{�5j�.ߎ_�B���I�� �U�%���[�kKmT\i(�������̈́�C��^JgwT#{�Lt�Eqd���ᘎy뺏�w�	x�=������\�dcp�Bq풪)����A��0��C��bC6�VX�$����b�ECJn��g��
vC�	Ĉ�ڵ5&���ü�\~hJQ��h����
=힔����B�� �5K���R�j���sKC� ��\�BH����$�UWD*����0�cC�&����	�A�=ɱ-\Q����Qx������ڻ�`TnL:w*���=�Ꮵp��tĘv��Nu/��9��AV�ms>�'9�~��K$��b�5���'YU�P!n�]8��`�7�j�]�B �������)��!F�yV�V��;˶�˰�Ð���tlD��l7��2ӫM �P��K�&๺�"����W��К�A$g'h;��0���!f$�9�9[ֵp�]�%��S����y��שGD��d���3�����)���̥�g�sm��a�7��٫�G?�u�{8[�iv=�Wc�
[����0�ȃ�8E~�~��Z]C��U��G�4v�=�Ћd[�;�D75��]D ��s'��-I�Jk��J=qQ�K;�Тȴv�3ËoE����7KL
&rG�u�0��EZH������h��d$,��4�Bwj�%�)�\��E�ܫ��"��أ]Xu�����߼�?��Z�7�WA���`�,�WqK��K�;^n�d�+�,��D5!���d EԈM���B
����c)�nTI3�r����.�l��ꣃl�:�(�J��A� Y�?^��x��l׭��*5\�h�G[�[�/�R5��cs�ef�J�FŔoH�5�	�,n^s�Ow��LKx nE�C���6ź�?�ܵ��п�C�J�#a-���M��(E�aρU'a��_,�^#}$7�労���z��D{���W�<pQF��x���PR��w0E�.}jO��;D��׷]D\�-�
ZR�A�;d�ibrH�����|�.�"q���%nAYL)�Ԛ-�	��{l��t׸���{��'�8A����?P��F4��`s��H��؅0�7�*�i:�^o{>YucI{�dQ`P����#tP
WI-m;p���a�Zpp�BߤĪd�6r.�W^��w���#db����RW?klT2��]��1Z�g��-�Z�*�s���:��7jH^;i�@z�:Ə"�{��ݜHu�R��-̰U�%
H!�X��E$M���ڍ��$=�c��QU{,$Cֻnp7(��b�ё��Ub��Gs
h%���{dO��q�O�.N��wV������m�5'%8���j8�24��ׂ݆�|v�ӝJ�J
qHK�IEC'���:�Y��V���hp#>䰥�tί0�����>2BL�_����W#�,m,���ԯ��7]/�1����� ���z��4�b��.S�ď�UJ�r^$#���j�wTZkOI@�Ae���]YFCV�k �5!�F�^����c��a�}Y�!�Uh�!f�����+�m��*�O�?�9:i�:�.�pt��7 Wذ��O�$� �y�T���pÞ�6�,�V��xD�z0� �^q��K&҉�L{�)OgO��Zs�K�ů�N/���e�Z}!3/��L�	��O �kRo�8ۓ�;f�>$�)Օ�0����vu�E.�g�2ѯ��!�f�r0A�_����m�<Q9l���ݐzX?n.��bӣ#��c>�w�1���l�Vt6%��hi�������¨%�=�"�8�9��	¿K�����:�
+���5��]n�oy����z�6R�H�3p�oQ��.�w�1W����lA"���k�P�矘��8K�)31��<�~6.�@����ZH�$՟�O԰tRk�Xƻ��=0{��X
�?�X$��b����(;�U9g�q��_��+����y/��C�q"��ؠŃ�����xqn��UU�� �a)a eD�2<}����K?˓,;�����l�2��2�zy,Pd�,4����6X��Ҭ�/����J���Q*kyˋ��ߠ���1IOS,��*ApD `ޙ[U7P����u� �bI��/gĀ��)WEυ�g;nP�#����q�fvD�
��?�e�u����֒bM�y�'�J���2��R	�Z�t��X5����lO��Β<���|͝^��/:���~�@��H����s�kz}j��}�BJV����8j���ä�a1j
d���e&�Մ�ͫ]�=�� N%d�V�؂m���8y�k��==�Y���٦QF�Ձ�дgԭ˹/DL� 
r�g41Qp݅2�S(�$�Ѩ��HG	�&��L,�ǁ����~�OWEz�p'�vN�K�����C~��l����KD��Pm	�~;��[�8��+�cdf&K��G��A{
���dwLsˣE�m���t������W���.�2��B>��8���&�������bR�W��{d��,y�:��1h�b�8k���)U������m���Hk&=-e!8��JD)_����9>p��X�j3�)��������w=[��70ϭѦ��ޚ�t�0i=C3����H�^;�bz��n�F�{��9�>.sLe�U�QQ3���<�kg��"U)�Z�[@���$���FӇ�6���&��R<.u,tH"�cVo��F	�V�ƞ�J�<��/ 1غVa_��i�0�!�g�َ~����"�yWQ��� kZA�w�6÷wV�-�Y��PjG�ڹsxq^!e����u����D����Vݷ&��.:a?PE)R��S�?�����e�G-G�ش6�勤ާ9��� �@�ߖ���u;;q�h�0m�R�͖��Ҽ�Y�R����" X��Œk��BA���+��^��\f�a����d3FE߷�B�������NG	�&?���~��r����Í�}v�kY�;���4�����{���ɫ���:���`P��IK&�P)��l�yZA���|�G�`=�ԷX�����#�����C̟!j6q)��z���N�>uD�L��6��)�U]n6�����-���l���t���Y�?Po�!�U�*7�\�V_���ɤa� h��l�R����du�:�mɾ���������>N2�t����׼�rߒ[�(������w2��{��+��H��*֒�D�=����ؤ�VN��=�S�� ��&�$p���Sf"�T��X �j�~�B�d%ma�?&�un��%���ZU�����	�>!Q�s����L	]H�X���?�h����קe�ʰDj"�:�ξJ��d1�r}(`7F�u��z�W���D��t��mb��(c�^β����k��d!x=D���L>�|��z1y	��]���Y��������؃{��D����
T<c4��/��Y�>��6��vQY����
��%��w�Wpv+���W̗���8Be�N��AJR�y���?��ױ�;'k#��xƦL�D�r8���;���Ay��S�Vd��=�5sc>����y����˧�9�~=����[�<��K���( ��iFE �}폯<yl�A_����=2����G�+����ā��������XA�����[ڰT����}i�W��"���8��X�VS9Zf,�n�ʠ�)�'���so<)'S�$����:�!FL(�������uߖ���s�p(������@�s�n�1m��Ӆɯ��B>?8�{� �ڹ�`�+d|��0&gkE��C���ߦ���E,Uܞ��(gP��&�tJ�r ��[F���:�S�g|Ϳ�