��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������-��
1����yr1FUb��q�ej�IϢE^U�nA��a��"��� �AMF'�k-���޷n;m�o�}Z?��$Ĕ��L�h������g�Y]�)�}�"��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�?2zֺ�i�UCv�~��t_.> �KX�d��@�����O�2H�%��
����)�j�6�Q�؇0��E��:��r�;xՐ�>��~U�Љ��ӎ/s{p�|2}�Æ����9���ELedI��5��!���+&A��N�����q���j��O�/	��l&2��g6��jk4�K�*�\�͵}�-�f�����)_Ӡ�?\0,���6;���YaM�ܿ���@'÷>�!�Ңr3��jw�n�9!�J!�W�
X�<9I]�a�,i|o�FzBHQ��]�GS�-ez��1p���H��b���ɍ̝[I�EIF�F���h���l�;���z�̲�02Y����jf��?7�E<5\��OO*������E�{8<aE^�UAf� �f0^���"ϧ�����\m�AK/qF�y���_�����%F\d��b�^���_Mޓa08mK�F���C����n�n��Y��Q��BY�}��r��h�N+� ��|~OG5u�CJ�'�O��w��	��E���e�׆J��[��4_��^(�x�N�7PC�<�8+s
��*�r�[09J��|L�,$o��h.�G�C=����Cl�����U�Q �9v�7 Ƹ��!R�{u�ٮoZ��%��{�ԓ�����O�t���y㻲�ȓ��y���W�mX�O��({#��H���Oİ�v }H���_��4��^�<e��=�h]/��y[�C�� oCt�n=:�'>0��]��?O��e�r	UT:�s�eY6?�6g�NɖЖ�*'�]X�=d�e�;���l�Q����z�_����[u��d��Y� ͪ��[����U��1�l�^�ǜ���˰�F�A�,t�h�zKtQ��b�����az�y��x�Ld���7�Wq�t��@�D�`�nc�;�8�k �oaWP0=Z>	���o�u�0M6�}f!�jb&�fؿI$�j�4����<��Bؙ��"$��T�;:�[��b2�9��*U�����`�H�Y�g��-��98ù��L��.a�Y;�i���Y��MT�b�^0�7CzC��#�Ϙ�%Dz��0Ό��:��#����D%Z~��B;!+��tQ[-\?�����k��-5���$�j��%����v_��s������3?�Z���WϘc�>K܈d5)3D%7p�奷[E:�ء��ӽ��-�"�3��4ş� c�B:<ʆ�g^�R|����77�AG���n���A�Ki��J��qM���X��o�Og"y�Y�vˮ��IS���WV����R�?-� C�_J��ru��n�`F]�O
/�jg��"���������,�-��8�,�w�^vtZ�f:Č�qM��v�m�T5t�՛ˊE�9��.î�v|�ʩ9ِ��b;
p\�>�\3�㳐N� �����(��0�Jl '�wam�&���8dĀ����rC��#m���қ`�"���DO�u� \\�CZuؕ�ZI|>��aNF���rݬ]�P\�̦���~�rb$>uG��x���m��p�!%�E�F���K�Xޅ���V�j%Q���$�6�`ֻ����c�a(�qF���;��gH�R�/���,�	*���>L�����iҢw��^9:��c�%�H�Ff�Dv�fs$�e#Y���^8��k /~�wb��b���F��m4�3P�3#Vu�y�
+��NHćXf��2��L�z�k�-���Y?a�hz2b]=�Z>!��-N)'5�H|QN�.�#�锈=�b�����r�8�i^46�M4���T'���ug�,�x���̜u �LX[K���^Q�P�uT�C|y��1�+'80.�������MS�/�_�Kbѷ��pb� ?C�繭�N��9�X���/40r%��x�WV�0�#�	�h_[�}�W�d��T��R��{��qy��.%���΋��a�n��6���8�cY����D��H(��;�? �36)%h�:��~
fs8΋�-�6��j�9��\�e��UK�u`�kq�u��\�T���L�����=筮E���)q�5a�MK͗���+)�,
�M�����Ł���q(�8�ú�jz�p�D�,`b�~`�1��P_QZ�1�5l��HEB���a�0s�ُwp�N��*�tG�����1M�ialA)*�&�8�Q�>L���cѬ�{�0m(&�|�V�1aX�=),"e�Vwm-��V6)&	s#	�߆���T�g�2���s������i��km��;���Y���Ϭ==� B�Co�#l!ۻ�i����o:+�?�V�"��Z��i �-�7���'f4-��x�b�H�У���/d��7X-� �&N������b���s�����xl�c�Dh�TTs,>O"h�Dzso��'-����O��dZ�7�D{zÑ./�n��°��7?�Cd�ަ�!�0�V|�\�Y�T�jwH�Moǎ�v��5��(����Bp�������l���D�пyI�/As�V�B�c.zFpv3ˆ������ O�z^�.���".tũsn�c�+��[uk=��p��(��}9|��2� ,�L�D�K�K!�ФL���)�����5����2�;�k�������>�<L,�Z�}X�J%ڇ6%a��f:�yY�t,rUY���� �J�@ϡ9�Wt+g@���I���I@~uOG��MB��4�������M΃����k��j%rr��&	��ŉ��+�6-q��z��k�0��hZ�$�90ʔ*Vt��Q4%�h��V��܏%G=��C��$��j�w��������g�k���_�瑈1��
8�EKƀ�:t�M.\*��@�aʼH�K�墼�J�\�,�d��O�$E$5��Tp�-.I�JW`A~d�<���+��u�/�U�e��
�^{5�V�-e�;�E�y.a����;]'�Hx�c'�}ٌ�O7*���$�����as��wm,]����ΩA�p�ZD*�z�Ǽou@���:T�"�u^��>������Q����-�DA��K�^c(�q�:���F{��Ƽ�2-��9�C<��鐚����b�3GwHI���P�[~Օm$W1G�۸�Wq���{H���fE�f<FQLT���P�"&� ����N��|'4�̔s���1�_<Mk��K$����k��6k����D���~�>���
�[9úIR�Wo�p=މ8k�`|�}�����2����p�:~��z؍Q���	�'\}#<�@"�����uoe��iB\Ug�vZ�8B�D�]�:-����iC��w���w���]�U����
W\E�i�� ]��ޢƗn��@..=�����{?_��G�{�/���|�Ru��b��Z&A��yM[/2���T>��Ha�������p��g� �L�y�I�6,���td��^��Wcރ�}����ݝ����}���nW(KZ�KB�6���V?l���Df�����M�?�ݻ*����q��R�
T6v�Kr�g�6P�_���?;j�>Ӏms�๣��������P���ԩ��}�*��[�FE=~U�']�)~M��fh�^�P�a��Μ�Ewuܱ�����Q5(�*��V!�<N��s���3����,�c�T��jk]5�q��(�/Jg�j+ҧ�	ĳ� ��:�s�n$�|�3CT�5���F%��U�K0�X�&�ř���f�P%Tr:�C�Ӯ_I.�f�mnF�����kN�|V7��c�8���<�������f��ߚj4c:qQ�^�c��z§���|�#S������%��[�,�T��vx������.Vr6�'V\Ѻ��J�j��͇�d%����׌.��O���<��P���6�M0�O��̹����:l�+\�J�}e�Ѐ<��W�9��PSn��H�9"�^2�4��#ǚ�G���-Է���6���A�O�%/A@�(������vލ�l�6ǐ���g����D%Ə�֙��U& S.���IG�w��'��FC9qWIF;=�������Y�!$�6���|.b�<.���^�K��@[b;�f.~b'�"���azĨ_x�[�5�4Ӟ�~��A��f�\�<�J�7SU�[�UA�t���4\p���C�-���0�T"C�9��`��{��eݣ�3�E����򄟔��O�[�ķ�pg�]g@~�q,PDz�[o4D~�߯�=�!MX0�Ҍ�!|�`MN_P�W�O}�-�q�:e�ӌ�.�#��g�WY�Dp�5_�R���Dڪ�l��#+x�Z]Y{d��y�*z�$E�.�24X:�����z|œZcf�� R���a�(�Fٶ|nu�C�*s%Z/iWT�3�
|n�ȵ WP���a�O��BO�n�Z���E�����?:��uPdw��8%�m*Gm!�Y���5�
�+�
6�Z=���NZ7�Z�ڈ	�[t ��o�5L��N�O%d��Q��=!{�b���`��BN��Z���sm"l:�͠��E�h� �6��A�h��P9�M:p��[ڒ���pY���w4��T��d�i鋄R���0��2+����T���air�^�<R�1��=o�._��)������K�	���"T��=��w���LC�V���v�����Q�0:F��A.���F�樬_�ZZL���cؾ��D�U�~v�؛�j�}h����` �G�����OZ1b�3�%;��p*�ǳ/�8��T���6R5b�f�o��n�us��!TVJ�܇��-5��\Z�&Ad�ʟ����j9�^^����R����ݛ}�=�
�6��?���˯\!����9c4�A�?@x
��5�0⛌ɘ�$�'>���<s˒< �%��ODC��-��/�w)Z	�<8�o��DWä�6~6D5�
藀����i�i����/x��<T�<yμ;a3��y!�4d'rQ��/�+�ŵ�������ΐ��G�?�J�Sw�(�.�9^�u�����4w_h���õ��D���lD���ãL�/�@�7n�V0A'� (��\Hǚ4_���W�(V����6�͘�ӷ�N�1d�-ƋO^i4nrmY~�ǲ�n:��4$�Ϣ������w�,p��'�4�]�:�%�D-Q<�N�u���$��m��~p��mlV�Iw艹�)A��(��XİJ3lX1i��c�Z����/�5?)~I+W��~�%�ɧ�.�h,�ً�=��a!�4C;JWƶd\��Q6�3��TL��E���Z���x۔`8&t�0���X�p\���)��.axj9 ��&��!)No�U��%/X�ޜ��=Ҽޑ�3"Y�v�5�p̅��}��)���"oz,W��Y�T+R�5u�Gϩb/$����*\#!0r�	ju_�l��A݅[/�:[
ݧ��#x�ky�N���P9��k"s'��ɝ�4}��߰���x�Z�"�v���6Fm�.hf�T�q�g�nV�Y����_��ZP�zz��y�B$4m/��	��P��$�[6,!r M
� ��Jh�SX�\=7�hz��Xheɣ�r�5�Ccj�Z�њ��-|uH�4%���g� F`�暳��Cy�P�V:�.�Z]�� 1�Kojo�\����1����:hip����[^�sut�TI�>�mh�(�lzf'E�Z|s�K�*�Ą
Q��@�6-��T��o�B�{@�~�6ǥ�!��ls���YB<E�C���&�]H#���9G�>, ��ZB7�vk��fgFw�_�1bXW��<�S�~�8]�4�|KK���F�=��}�җ�SW�c������<����Q��?��E��%��L�6��
��k��ŏ�D����>�1�.�K�܅?�7�:���[p}��T4k(v�2��ę���d�CU�l	-;2y����/_��4 ��8��m�6�'�ŷ���	9��C#xfCs��"��5NűZ#-����҄�����ӱd7
֓ی�m�:��ΐ(?���{"aFK��Z�sI��F��%w�֊f=��շ��#����ná��d�;����V�;�ږ�,p��C{�� =�~��Rt۫o��۴��B�9���S�)����]T��+힑%��al> ��݇��-h���	.��]�a��w��b��,�/�&��b�a=p<�6��x��]��n���@�2AT���|�C�#�oyjC��O|�)~Vr��l��)�eYk�Γ������h�oQ �5��&�9b2w[G�(���O��}�D��܏�V����;SyD�M�Ih-��[��R��86eB�!�<M�M&�=ŭ@�L��YA*��:��E�.Eԍ����'@%E�D6��a�h_��<��\I��c�(��hif��gmQj�'�B*7/�������u
��@r2Ƞ!��Qv�j�׾�;���	���,�?���o%����Z|?�i����#�Y�0���~ҳ����6T�&��}�:���Ȇ,s�&�#Ϸr���P~1�NG�8������ž�u�u�%H�̈́��`_��4-�{x�6�jZ���~/1��}0���pS����8��2����[�i���u�-U6���Ã��N���$f�w�U �*asE䑏R�r��|'"^����?�L����;\{#ށ�l3�T�y9?n�s])�7=:��Sj��o9ߜ�d�	�m�=������F�+�H�M<����h� SPߵe+e��Q�K���HNs�R����(�������!v=kt0�<j��L�3�yP����K��Bf*e��ٴ{2� ?��7����E������_u��/8b���|̅�ٌ�����pƱ����ڴb����&�3(�S�R��gm4Z��o�#H�T;���B��ұ��u��#V<߼����s&6�f�T������CG�����!A����Ŕ `l���&wm����́�:xT���|G�Dǰ�gS���}2��`��b��x'��Ӆb� ðU�9�������~���PR��{��m���5�ZX�%�#, ���kY4�����:�?�r��X*p�7D��W#e�&�P�.y-L�n��ZA"Hw�
M������3�O�]q&&%P`��"~�>���w1�X���5xy�� >�r�CR�6f�5w.���5��s�z�ϋ�!0~���dl��>��u�u�.�F�����^���Ӟ������X[�xW�����i�+�U��e��MRUq7�R� K��_ *o�W������M�tUL��'�WY��4g�L�8}�"F\��A�h*�v0P��ު	�S�=!�F�eq���8��f���<6��L]�CzJa~��	�N�����fsi��������3*���߹�L*";�H�;~�� 8�uS9?f��"�L�h���DM��=�z��ٍ��j�^L�[񜉱m7��xf�)hvpMq���}�Q��@bNe�*�z�d�J��B�%����|�)�g�:#�~~��{�Dg���{��˷s�M����uAu����p�O0��@�ue��CI�9܈����CrQ�t޲}�|,s��?>A��GUBʏ�Y��c��R4?�Vk{��|xR���vhS��I1'u����1щOT�C �<_2�=�2�8��>�~�?���`�w���X"�QC��H9ʒ��b���6�b�Ո���r`��W��?������ODZ [���Μ6	ް��JP�'mҽed�I#}�+j���Yi ��&$� ���4y�p�c����^m�g���reta<�BҎ�7jO�ZZ�WpG��y0{��Q~*�Qo���f��Qkұlz�yyTl��^Z:�`1iWj`o�\%����S!�lg�ѴsB#;N�f�=@eA�>�W�t�?�:A�#D3�`T���Qrf'T|l��nZ�z�F�D)����*�G(��	�B�����O��,D#�
�.�(�q,4�7�9��@�u�x�8	A��hH�^w��N]�1�J3�0ؾ'֟L���BUͥ���]/� �
����؜�P�*X��Gg4f��}L��<��O:�v�IC��ڪQ�y@(nL*�C�[i2ߋ���[�]�WS9��'�~f���Oe~�^�z��Z�n�xY�IM���4Z!+�!/(/:BS��9�i��-�!'�p��6D,�aGl�[�4D�\�:��w/��LmF/���W#;K�p�͇!�'$ݲ.j�.��e�+��{|��pPҺ�����|� dM��w&��B�,t�׆�.�w�����.��ʔ��َdtկ� � _���r�?>�3�:\��~�����}Z+�~Km������U�X������!�#F��b�m��r�V��k��A߂��}��z�4��/Āi�Zl"���A
���ofϪO %��w%�C!F�۞�r���X_���T}��Q�ޮM����cE�A~������s���!���^8��4V�IySD�Iy͞��.>\�&)*��]������8d���E��� \���z������;q$�-����g;v�o:R}x1�w�[N����&�D0�\�n�IJ!�K�)��-�~�zm���������ޱ�_�yؓK
<Q<�iD���J�7�T�I6i�<t�c8��Y��	��^�x�;BȖ��)&g����wir���S�D9�G&�I��]a({��ވ�b�J)�)��K��@�5���~b���d �E�C���m���(�Uxo�@ա�j��A&j��R�В3[VB	����a��!-wƺ4�x\��#��o�71�l�s��s�h��A�Dב��g�-�dT��N�q�� j�J����PK�.����0|NSOWZe�D����+��^�g��5@ƹТ"_�M�|�p�Đ�g�l���_ݠW����x<!V�"$xH���P��j����D`A]׉�[�͜�Ed�;H�O���oX��;h�a�.�M p5C [w�F�A��:���N�p$�bE�ǸȲSF�2�n��;K�ɀdӁJ]ik�N�|f�l��_/_�CA_c��?I����>#.2+:���̄ܐ�6y���P�ʻ$�Gu@*pyt���5�����LY����)�����-5�3U�Q���q�9m1�%S�Y=�R���;~֟(R�2�I.3T������{�Ժb&s	��H�	kt+�G�0]��9D�]�Q�N��E���,���+�+�~s��-� ��h�N�֓�!�``��I! �mKps$=��_C`o)����x�;����5��������������]�":��Y��Ḁ��2g���w�]� $1�3��sF�����*P���q'z�j���\�5	�FC�\���qP��$���a�ipU�R�Ӵ��"t�F3� $�c?����ί�"vZnV.C|}>JA;^�M��2g�н耡��������g_���y�	�r'ՋD��1�7�����''�*�l�Oo�*x�����3��T�2`����#����c��N�����EN
Rwp?)�� ��n�yI �VeTc)�	��D�|+`Ș(�c���O��_2T�)Zw��b]��abǐH:5=5[��"���iY��χ�ݲ!*\�-*������;��u����uk�S��:���Tk���C�;l.NH$:x���xԯ�m)��&�f-7L�L�B�U�q�	�?2��9?����$��=ǘ��1X.Ȋ�A�W�X�Qf\cD9)Y�l��Q?������"�;=>��­4w[��R"������K��_�1>�
�V��t��p�������I�Q�e]�M��Y>x�F>���hR�m�P��)�Jh�q&��6EԄ_˃��+�%^@�v��P_<�"6vѸ��Bo���0�o��B���G��aET`��<���Ȍ��0Diz��Hw�m#�+"z �#���� �����Y@;]|��/�T�E[1�MU�nx����惐f���n��ÇZ]�h�#�~���Q�CSo�3�����?���� ��8`�ބ�kæ>k"�r��x��.2+�����M1z0r���K���$AY8�pS(�-n���>���4�~\���]��.P6,׆3E�(=�g�V���:Di�\���_�F\/�i��)��@ ��0��,i�J�ǵ�ύ��r�U(f���yK��؏�k0�\;�RM_�\�!�����ش_���3�5J�7���}�A*�r+���uT�#
%ٴ��9Jί�iq�q�u�͏Wl3~a��V���d�k�R�����U���ɓ^P�R4���?�~C��	ҳ��� <�gy��'f��'a�V�&��\���)a�l
گ��ę����聼�B���NV�����nĝ��۔� �:q�ce$jJ��7�����V��V�`ɉ��#5#���0�_㕡�=�(�/`��ث�UO�x%By�Ԉ4v�>h��2F�#n��KW�� A�P��k�V
�l/Yb�`A�� �$u-�w ���Sy��yZ�(�$�@�sx�=~�n7ÈK���|[��c�4�:��r�%�6��e��?�ds�
k�ߗ��� �[ ��O4}�'�IҭD�9���� ����z��w�K�1��8� ;�jm��l�<�Ȁ�~���p)f�MpJ)�IcBQC�
�s�T��7����Fր#��sG3���;ʈ�{~*���K
ضqX͇��u����i�I�Ekox��3�&�眓F�R|�J�T�E/!@F،�+�l�ב�sz�K��h R��Q|���H��N`��t}�B��a�i=?��*�jڕ��<n�g]���7k&71��j'�j���g�3��0T�����HOU#��!(p
	��p`���l��|5822�(��%��c������\65�O[�a�'֗��:2ϡ���MNNK^�z�ě�*j��V��G�w<��o��L��p嗥�A�#I�N�I�.I:hɎ'8l�wԒD^Z�����1�Y�zv�'�S�.�\�3	ڤS{w��4�������[mY��!jln�π��Í����ie�
ב���_�]?3�"�\"y�Q�/��%�@����Ѩ$�T��o�o�ό��"�n��&w_�Q�Q����4L�e���}F)��\|���|Y����/*��;�dʟA #��*9~��8�d��<Lg��%寢�0��*�W�<��~mv�W��"�H��ֲ9{G��an7�}�d�%�f��]U �t�S�-�T����UZ�u�L����E���wAؕ�x� .B���-�C�,��Ȋ�����~	~9VV���0)�J�1�MLo� �1�Z��E�y�!�I�Y��G@���g�lbԔ|	�w����f����f�~��k/�xN��0�������t�;�U�5�$Q��0�X��A��(�{�_�Іh	�vk�vv���}��2�Z�2�׺�&�J%T��������h��XX��y���l��x��Y@臫3I�uh�8�c4-LTr&*��ĥ��J��c����fꉺ"ͺ�}J�ZvttL��Ø1��1��F�`�Γ)[�]p�*f�	D��Iܾ	n�ל1��6�B{]r5~�W�Hx�:�l!PQSV&mͬ��,�� ���[ZW���
#}u|�t�zhD�hӳ~;�|�W� ���1��ś��:��#9��N �ؚ�C?��8;~&N�G�{�������/�W&�` ��;��uؾ���#Oj���IVw)��F���&�a�"�b�	;
z�)��' xFT��J�y�f�8�x����a�2Ĉœ�tGqr���-��.������s�6B/�����H�|�I�4�T����ZR�"�� ��<V̚��>H�,Cv�^"� D_�{�LL�a��ݧ�O�txj��F�t5��ʢ����X[�'�]7S }��+��e 簠�B�3�7��/�|+� w(��#�a鱆��	@?�.��� �OD���n$�(+F2��'h=
��-B����?arp[/���*�ܛ.�%S��m#�B���:A��T}=g��l���o�=t+���/9N���x�ќ�I^wH��Kȥ~��yP���{b���+��G��0�[i�_�u�,�w�ȉ$�$����'�tr5Ae�~.�,
n
�;&<����<���ңǸ�t n�-�gjA��]&V�%�B!3���sD�J��S�V��/�!Ij��I����� R����M���E���T*����Qa�]w���ymSN ����,��?���~(�[x�춒@Uh'.X���e?�_8/ߔ�;��y_B#���)¿�F!��hz��Ӛƌ��)cԄg���I�[�o�%��@�[,���X!��@xLq��܆G:�k��C/!�r��l��j��%�@�&��������r�V��O�u9 ��ՠ(#��O<��9��uj���Y���`N�>a� �v��~w;����*h�����C��0���V�bu�J��m��c;�(�﹂��H�:���'vq�u����,>�ə�f���5���.��S(&�w�m��M� �`�&},��d�ݙ֋;�6��I]�p�y���_������\= 89�V������Qz�[c�[��v�u�z��(�ݦ��1w1���>Hhi/�Kl1�̕���r�u��_
{���\�Ɨ�VT��t$��d�[5?���Խ��0k[�/�9�Ku�<�kf�l����y#��T��vh`s��a~�e{��jy!<���^���u��;�\b�[�9�`�3�Dbb*7�mA��b�7).������N)���a<m�AS��\l���io��r�9bP��	ٲ���9��}݂E�i&JB�)zR�TVZ�~쇇<�p6���V"���WLtO�(=�]��-iں݃>�`IŐ��b��w��>�����9Wt�9&=ޤ@i> 5L};"��)�K�Aހ���
Y}�@��U�E,�>���^㈹�2���������A�m�o�8k8λ;�[�]�	����ɧ���NSѤc��kFX��5�]����+D+>���#? U�����1i�|ފ�n���1�4��h�����a+�D<�Q�o��͉�Q�dw�9��f�[��R����>���T}LF�!h�<�������� jzq�6��� ���Z�Qǣ�e^��cǢ��u ;����7^l\3���%9bx�o� �!����q`Թwjr�bU�Z�?g*)���,�W��,�Wz�Qjs�8>����3'����O'���(z��dr��.�X�#y��q�\Ҵj^6A|��<&��2��^��s��Of�kX��R9��M������)���o����A<�H���*�m�9����U�q�i�]ܵ�j�W~ѐjz~�w�^�e�iry�v&;��؉�.��,DИ�76�E���^�O��G�lP��f���n.�{d�o�=^B��e��Z֬[D�r2���Ǩ&qP�]@�SH�&�Z87(|���5O� R�(��j5Q2K�G���X7]"���I.ۡ�=���l��l�^C�^�茗�Kn2訯g�t`6��YT|s�$�	�.?G��g����v��ck{��>��#TF�gA_n��y�pݜiA�k���upx�N�A5�L��S����BSz�՚'O�����A���O�I��I:%$�����C�8���>�0�i|�T�_q�I�iԂX�7՘�	��8%�ן�oU�Dg8��:���^ҩ�;�V���K�o֏u'R�ؒk3��z�-;��Q�q`	�F�� �#/H"�t·a9��<.��1�4��^L`�/�C�5b�o�b�j1�8�D���s�J����ݙ&�@]��7�̙n�(OV��I�4�4,_ڊ�ԓZ�1GX�a+���W�P���pIғ��i����Q���3�A�昭��1tର)˲�5h|���vϟ<Ď����VA=w��_���������VS#W� �Q3��V�#��\�g�� =���޶i�c۾�j��;:0$�Nv�������ou�v]geF\|?���ƥ6Y?Q!%>�EN�9��(�d8�c?�u��Sj[�.�i�i���)A�'�L��^���$�r趶$�����*�1����-��K��D�5�e
-����g��e_�#<�)0?���'G��E�a��lRLE�u|�'���Q�Wc���]�>T�g����&�T��Pihi���p�f��"�� -4���,��Cg�����Ay:�i|H>����Ԁh�}}�*q��L�;�2f���[���L�WI�kXr�`wۭ~b|����F�;���M?g����x�q���9�/�����1��r+��2bo��]�O�:mnL�7�Q'k�=��+g���	q�T�ԏ56�	eߨ�a��è]�,'\rC-)�u�FݰnH
~<���Е;*��8�hTK�;gZ�&Rک=Ԋ�� �U�6��,A����M�$������/e"�rnmK��{+�K���6���d��*;ń[����퍕y�N}%4�W���n�8Qg�g��,TGC�F�~� 	�;�W��8D�R��WUk-ǖ*S�m'��ei�n����N�~D��8�Q��;i1K����ߝ�~u,SY-�ChK6��F���A�����/�Nr��2��`e�aw#&!�J90��;���Nw�D(��\�8#�T�2��S��%y�|��jEN�?��BP���r�֓���h�{�c,�)9���B䆰A�]\�uZ��0�|3��ٓ&{�Z�;����@���]�t�u��l)�)�f+�.������K� 3��Y��H0�uE]���o��ib4��7O� ��>~��H�ͩ�	]b������'��Z2��a��Ռ�b������wzK� LD����0�*c�v>���3g��:%�"������:��/w�H��S���ȏ��c>C��a����������I{y��]9�/�q�\���s�'� pj�'1���xt᎑h��4�K3%瞧��@Bн=h���HWɇ�1�u&/�~y��&-#�O��'%�{������t�y&"���Ä���Bt��Ճ��<A1��m!O���$��%��ͯ��%*~���!ڡ�!���V�,Fjn&�{��`�T P�L��4�����6J����0��5���՛�����ǈ/�St�L	��ɬg60l˺�
.,���5�?i�0��U�PK�~�;Mj|s���@�OS
�W!��%�H/���ޯ҂�A�;�y�~"��0�i�ؽ��_˘�^E\s���H�R��7��@��%d�ӟ���X�a_��d6�T� Z�������4z��L9��UX�Tq=�\��`�X�g��3�'�Vn�S���&��b��~Lb�븩����Q������E�DT�|jZ/������|�j���5�^�<?����%�'�i(V�3*�5�+C!��g�k�_b�����W~$_K*��yL�2�E��rH1C�,E��g�F��+'�c����s�Khf�eǿ�;���I/4�6]];r����ڰs��͠�J�Y�j8�$K�U��@J&�P�y1p���t���`��FM��0'�����|�+dY��:�Fg�a�ޏ�8CQ��ޜX!V�}�A�jH��B� ����o;���X0|���\5t��2��3y20
!mM��=($�~�����ҡ�!��=X��K�W�уC@�[��~4��1J��Ym�3��r�W�M�F�9@j9�X�{�V V]e�y&)?�Z��a�pe˙�O��O�$��+_�D����� ;)��,.K^_$c\s�(��A�Da ����ŮqZ����t���Ũd
�̷+���ɔ�-?�����ր�����X�*�����@n�2t=�w�-b|'�%��O7?��e�w8��*���CrRy����=�B;�B`b��}�Vz�$8��V-�AH�4�?ӄ��8~:rv�ѓ�cj��9�Q�tN8��o6�A�E����$|U�f�	�����$pm�X�\j��
�r���?"X\I%�	4�Jچ��K�R��la塝 ��D0$����Z�d?s0����-��1�L\+�d����(��N ]``P�8�������QK���$O?@G����rfϗ,��WY)L�IPH'~ :�*X0��������]��Y�!^��䔎�_[�~��˔_���b�g�P����������ŪKf��*Ds�4���5��Sk��M~����1"#�,�lr���p���-����8��3�˴�㈩(��6��@~����ν���a��b�n�Z������~U����k�埙*p��F���A���mgI�PU�m�F�ŷ�V�PF���r{H�T!�Z��s�@��}@���/Y��gv^�RgUv�\fj���5�-�P����#�tj�s^��˼��m��7R(k���D����bv�&+YO���Y�����ŀU� �_�J�D�Bb��I�����O����ǱK�UO��S��Sa�=���e���Bۇ�p�{`����)�
�-��K�in�ɾ�ed�ω��uo�`X���������!�\8�e
Q����AiA��rK��0��
�.��4X�K�G�f��:�OoD�OD���u���3;N�Yj���Ց�ۘ�aML�n4<�#�ɷ[������9�Mu)a���b$n.�jN��6*�����Z�������ou�!
�d�͑�~P2!��W�˄C:$��B�����+�Yz'|"JP�+K��L*�f_��k������D�L��l�N�hk�S���� ��jXL���b�ps�p��#��c���.����SL�b�7X�9m���B��u��97��oY��J��@���8��\�T�{�=M�0ÿ�V�wTt�:>�\V6@eҚpj�[9�HJ�U��S�*���?W�P�X���(��{�X�h�MZ����I���iS4.��s���g�r;L�,�Bb�3q�<:�?�4�Q�<���ޥ<��_�dIKzZ������5��/���`�v]r��| �@�G�:�ބ�N�n�F��0i.,��P9���W���}\�	��q:617V���o��ߨ[���� ���:�"Z驠J��FH��9a����HQ��3X[Z�w%���%P=T�!7L����i"�@}��;�<N��Q,��,ǒ<
�E�	��z�cUǧ%%$��Cp�G/ɬЅ�-��b��-�k2�R��"J��oͨ+i���J�%����2|{�w��ȡi|��p����-h��1�3-���,N�}@c�a�)�3ErfX����+X�L�,�N<�E/}�>��4F��LlT�¦��C����U?��V�����;�] ��O-gF��0��q�jd%>/S`��<��G�GN���~'o��6���V�۳����ųYd1�] �M��j3(d�3��~���/=���c[A)�MC���	S�^7��o�W�"JŶ�R����aFw���	�bޕ��	s�X������ia1���}}�H�@�X����%;Dd��p*�T=i���J���g�b�űJș�t.��3K���ɳ�?�ß�\
&MF.L������:�S��>���n��$ny�w�G�2D�]��U�����R��1D�D��+ubw%@�.�\��O� >�9���:>si����ı�i ��}�C�ۊ\��[�I	�n���z�˶]O;��%G|z�v�-0�-��O�\z�Kglnq��?��o`�)��&���Fz�U��ǰ�H�zE�ةؠx�V�`�ϨF8%��&���G�C�t %71�D�^:t�N��'o�T�v�rƜ[�N��EB﬍Ӝ3�Y�V���6��Ѭ��\����b� K��~��S:��E�	A��;�H�}�����љg��M���L���-�!�\�
��xm� c�<�����+8�p��6���Z"���v��(���J�zS8�p�0-! �A��g��u�0R%77�<���F
�Qsz�c�{��>�9tA�m甕ї��0PJy|�x������ߥ�Δă���X6ь5�_M�+4N��V���Z1�����/�Y~=��p,�{���i��n��w&�E��M�q��8�����m�P����U�"�#��ԍ�9O�*��:,c�ݺ޾�7:A�)�A=�8އ��V����=b��V�6D7�Y׊�4n�����'���L���<��
ʥ]��a	
�!/�h�'��LJמ��@�ء�dԱq���_�wf�XO	Z��W&_(b�� B�J�H�`i��Q�(b����'��Ϊ��?��� lju�+qE�.o����5�m=OH��[g��3�2���7 �w��L��YL�qͤ/�V>�1%~�������mKIRS@�ZKɯҽ��Z
YD۞�1}��X�ad��������5�x�^vFŖ�	ɵ�ڎ�g�9
��$�����4@���gt��GN8��uҁ�Ѧ��D��0a��T�]̯�Ӑg��-��j|k�=�"��pe)6ͧ��_bz 5����ɣ�5!"�HWc�	1��Q)��p���VtB	��Ӳ�������5
� ق�UnN�M�͜R��->ix�;�����x��IC74�O�5�Oσ��ƜDq�	�=nB�C��T�G�G
����x���,t���]��G���)9ؕL"�~�u�ҥ��7$I��Zi������羏�4�֟	*UkE�m-�Y��Vw��D^FǾ?z3��Rϲ�JQ�'�f|"O���t!�̄�`I�J@�4�����݈�\��Ý�iPG���a���9W�{f�����gWS��[g�������s�2k�ďV�:؟��r��*cMl���wT%���*�0����(�Dh������ C:�5�����^Bx�?;1D?.(�m%}�^���Ab����-���ө��ֹ��2SF�� c
�'�w�m�ZaƷt�sE�O�0�:�*/��:*���94�E���A�Q�w�$S9�����JVj<���n�V��l[(f���^_<�07l��c,�=��B:��d�m�Qڔ��B�����_˱|
��kv:�-d�P�^&�aa�U;f:�_�l�,?�]��m������Zg�^=���+R �G/����	9V��Z3%<ھ]t�Xx(q�ȳH��5�#479=\,�Q��]���8++IT�{܀$��C�^B�'�����*��~͑/�?�=JJ��d�j�A͍#d<ħJ�6F^�U��Lp�2}�Ё�;�Ϸ2�Lf� ��CГ�d��F���~Yc8��7�nl�O��7Mu �5a��o/ɵh��z,�Ae��q6I�A-lN9Ҋ��	n�_�V�� �8z������c���"�F]��*0����$VaL�}ԟa\�`��($w�E���a��RO>�˯C־'�ߺ��,?9�(\2�l��W�{�]��g֢��wYua���m�ڟ��,{HV������W.��=}_��R��8H��zTtE�kJv����@\m�I8>�>�Fh�X�E}��հ*%n_ŝ�7��o�b&@X!��K�&,?M)8s+��3?_��Vx�6n)d'S�.an��3
���?m�M
�AՉ	X����WݜCV�Rn�d�T�7t��\;Y��K�kv&���(����w"f�ޡ��E�