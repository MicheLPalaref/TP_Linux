��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������-��
1����yr1FUb��q�ej�IϢE^U�nA��a��"��� �AMF'�k-���޷n;m�o�}Z?��$Ĕ��L�h������g�Y]�)�}�"��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�?2zֺ�i�UCv�~��t_.> �KX����Q�!�N���k�
]�[�a���5�~��ѥ~�_!-�Ǵu�k0��s��@�b�L��Ih�.@4��I�~�l�*K��o��6Y{��� �U��A���:N��-2�� �ʦ@��u㋝�#���(E��(�c�J��=ZfF��e�R	!��;����%L�R<}��m�X�H���ڱ6��ߨDEfoţ��LJ&��E�b��[�cڎ�̔�TgZkY��gFۈB�/��L����i�F���_~�O��X�v{�8�̥�A@.�+0m#$;C.
�w�N�9��h̙	Dm!�8���Ǵ�NYY�WX� [y�d��ҽ��Є�s
J����C�4����{�z��������x�.��6�ŧ�9�@hP|�~k����~4�o�$��q�0f�%�vie,�@U̖O��B�DT���K�yf����R�^i��:�Y,\��Q���~�[C��Q�P����G�������Y�\�C�~�}�s���ԅ�<9�$��w��U~qn�9��Ɛ����w���L�*v�	<���4�F��p&����W�b��~�����M{} 6�O� kJ\�y����L3�YC��D����k~�]�Ŏ��8N�-��0 ,LKk�� aG�QWئ��ى5����yv��U}Mg)j>�(	o������)Sd\��
�z�/z.Ro��?Uch];�gR7w�;�ӑ�������f-fF�����{S���Y�aE�1W�	�m2��,_���J*@Ν�e8cS ĥ��������r�0v��>�'b��+쥒uO(�v���􁱏�ƛ"j;��|��M���b����&NJ�� �(v���u{#����ǩ48UD_��@V��2�z� ")爴��kxuJ��䚞�ͻ���6s͞�si���0�]���Kq5��n� ��SW�h9���
ĝ(�X8���HR��M�����)� � �q�H��[��U)66�9C9���kq
�`�ѣ08�'�)O��Pmj�n����*���ӯ`���c��I����#�~�c��9*��s2.����~l��$/�A�Dp�ċ(������D���ZO�gsB���ٶqQ�9&�צ�J��\Q��<����h��=��zW��_��cZ�9�}�Ӝ	��0�&ĳ��~~�������9�$��')+�"�ynŪ��SU�,w-p԰g�*�V��
�l����Nf:�o��$/صj5��gӑ�¶9JX����gI�ο��Cuj0�8Y"K�6P���6�O����m��B�@�*f�|m�fI�F5!���)�>�q�u��M
��i1����Jz�vg�ϕ���3F'��Vψv3�m�Bw��y�m@ݍ�/�N��Z� &�ϜR�3�*����$a�d��8
�/d:p�D���SX0yw������8���(粆T�h�: �WEp�ۏg�äW�:yB�lR��s�O�P�\�C��S�~��zM��'��?l8�V�_��	�b'_��)�y!R�s��>&.#�|�L䷧5x�ė�+�-�J��%)�s! ��N@C�A��}R��F�~B�'�AsR�O�0?i���5���2��$'Ȝn����Ņ]��' %��U����7M"{�<s����ڸ��CF�����5�:�'�0������ɬ�����6�US�7�܀��
��7�.�7���",,�N��ݐ���(�ֱLG#�4�&s��b��A�h�T�0���23W�aa�QC4G_YF豨������U�v�(�4dݯFC�<�+�Ge.c��A������c�7��}2@F�"k[ޏP5Z��K��'%�hZGޕ�;��Xf;\�����j��)��[V�]P��n+���Q�%�ٷ���o.*��P��Z�ϳ}N1�fe����	�n >U!�9�MӲ��ӆ�u�Tx�md�}X�A�8 E�2�6�1-:2f�^��s>��?$�0:��ԯ�<�@M~(Z.����"oX�|D�PU3�PK���2�Գ=l&>�$$�"�i=b��!���x7��?:��3e�c��j�w4��or,�r��z��6m��  #��{bY��c��sa��=�- �`GJ�Ȣu?����:�a��|��,�\.-���
Q����5!�y�0�[�k�������斃���#6v �+����0��9s�s��;B��{�Ԓn��	�9D�ۢ*�!@�шH���ĕ'~n�<�G���dk{r��Ѣ[�Ѥ6zl��
ǐp5�7���uH ���+i\F�p�ŭ�����AY%ZC�F�Ͼ��`��T%;Y_�$g��bn�r�EGz;\�zB�� /1Zz��ܛAӛ���Yk���&�@���C�G&�9�?��*�C��iW/y�+�D���=�P!��;��Ō���Y�k��t��Ӄ�����l&���&|�|TJ��#��teh5aq!���5�Ƿ���� �D*���4�7���/�6�b�h���t~��9��(�
�Cۮ���ӽ�գ� �3ρqo?Iց��H�2!a5T��N�nZ��1z'���@}������G����O*�{]Z��#,O��&nc��-�mmR
F�/O�Rxa�()����g�9*�"�y�.�,�URz�՟���?V����J���7�C�n#�{*)NF����>��o`��ڬ/9�!�j䳦#��2!!��B3�Gm����^�~EI�����5f'�J�9�����j}S`B�l<�h\kE�ˤj����
�r'���_����e�:�~[tӮȅ�?:(���0��Y�8��n;4�F2�0M�HϪ�A��'.�m�(�'.����j�k^f�{{��K�h=Q��s�7	"d�Z+uK����J�ZwY}�.������A\�k�_�������9$����vH��~_�Z�= �?-����a&L#3P�fTsg��2ߺ��<���5�ğ��(��h���DWm��k� ��dD��I>�!���𜺘�3l�����%����c.Z��Ta4�����'b[�Vt��/s�Q	b��Ϭt���1����5Ilz�!O�����Ap�2� �Z��4�³ew8-�RI�˂���՗�-�Ȍ1R˴U�s�k�;7���CU�!�Z���)3g6�HH��|CϝA����>�J���F��f����*wE'~���^d�vD�u����I/B�KЩ ��x�P2��ҋpK�|bٲy?<���wC0����Q5�9i��z�V"���yn<�7U§I��?��^���B�AŚL%��~���]�M'F���;��B�ϙŸm��=�<�.���=jؚGt�ܯ8�)i�pj_���ŵ��Y|�b�!��@�O��h����nQ������Ķ1�Z��N�	?�{�"}>�!�����=԰��n�ܞ�Ō��5�|ɍ;v�ȳ�Wd^�����0YԠ��8��|�/`6�T!<��V煼DkuJ�rM<��P| ���B>LDr���7P�6����)�h��>��dQe1f)Nk�_���?rbƐx�.�=߰g��T��R�z%0����
�hd�12Q�ۿ+��2��K�"�g8e*�*?71
J]�Z��G�CN�+��8�X�|�D`7��uCKm��{A�\�Ȯ	�I����Ӡ��&���W�
8�����t��O��/�H�t�5���U�"p�_jh�J��_���OZN�A�$|����ۻ3��DO�:&��8G�e�a��1l嶥�NG{� .� �ٖ�p1�&��Oyk�����뢠ѠpҞ*�}��*��a������^g|���
 �ȩ�6�x�7�&��
��6�I1� ��,HB�:�4���cDh4(���9�#�a8��ad���e�߱��ԗ=:��	�����L�DV��K��-���BGi�'�9$�� TԷh��DY��ɒ�1qs77>q q��г����W�eo��j�P#�y�b���:q��g� �.D�oqXl�&��r�](��L� ,�E���ph�ْ��9L��$��!�����U+�@$U�Q���o�?��g�@����9�j�����0��e_��a��tiR��Ӿs��-ǈmˏZ��-�p�ZG�%�G�i��B�d5P���P���@S�Z���$_����q"�Uv-oЊ�ԌS�� ��(�ͨ�p#w�{�Jn�����j��kcM��?-I��h�SV��~	���'�!�U�v_�'۶���B�U˶���qɅKh�3��dPO�-�70g����\%��
t�X�uP�W�y���� �D��� �B��2��[���S��2{��od�kI�h��O=��9V��[�ރ��,}N<(�Γ���v�¥ 6�L;7=��\O�X��U�c�� �_�J�O���V������+�al���4�f%{� |Պ;W������)�����	&�3f���E.gjX��q6�E�v���ۮ!i�Au�%�&@d���S!��69Y�����n�����-�w��&���57�Y��L�P�V�4у�s�VI+�	Ӱ2�1 �i���i���T�d�/K�ͻ�Sfbg�Ӱ�K��|`s�q�`O�eZSD��ij� ��^����U�=e��Q�R�. )���G8��I�C4:	7��.ӈ�G:����2H5k�u��~�$��P]ѫTq�T�*�7�W$�Q���nG��(+25 �M>�@�ǑƐ��>'l?����O�\�?�?F�t]�&�e��ܗ���yn�Ȍ�4�H�l�9!0�B�ޖY�C��h�}�x8�މu2/��O@n�%��m���"�GHy���e��'vD��c]��$��*'�MR4SE�8~�򠃳J�#�j-�X�K6̋.���Aצ�������\�-P5��ԏ��ؙ����6fs���F��9+\ua�(a�p����~��";�n�\oN�#���S�����8T�N9CQjGX����6:z[��Y��@^�;��(�D�S���Y�u�~ ��C���?+���Eӓ��|�ï� �0�ުJ*�5!i�y�n�����a�+�M����`� 9c}�'���4�_�s�F�Y�'Uf��V��N2}dk_L�7e�$���ʜ(+�"�~�['��l�VD���rN�FIT�M%���lc���Z��R��6����cjѓ���%��'����nƃ������&�}S����K���T�C�&&�tx�)1yeS������W��Hg	�m	�`Iy��
`�P!W���|!��e���P �P�%�'���"�D}����WE=�q�n,�ӟ�o�å�$�bygv�%�q-��2w�Xt�)�&J����D]�̓�m)>���tFY����f�q/�JJ$�8VZxg�)׳���s�dg�u�뵰p���Zi06S]�'�<��P��p��V�\ȴ��E
׾���"��&�&.p�=[���TO��9��>��q�qI/�����&i�㌉�ݺ�p�z�����y�:��8�f�d�z��<D	TO�|�L\S=�>���6ާ��:�?�?�E�T�GH�I����)���?�2����������3a�sw/��])�EǼ1�$�݌U��|z6�)6�2�ZyW2wI��G��f��9��,KL����Fp�V5�~���PC�F�������:�g����8�ڞ���7v�>�D�jBe�����R��N�g)�V	�߸��p!����c�eE=eP�� �0;J�0�Zy_;��e
jQa�Gُv�!�4u�|g^0PQ���[@\�V�G��W