// soc_system.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,                          //               alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,                         //                                          .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,                        //                                          .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid,                    //                                          .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,                       //                                          .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,                       //                                          .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,                            //                                          .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,                            //                                          .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,                            //                                          .vid_v
		output wire        camera_pwdn_n_external_connection_export,                     //         camera_pwdn_n_external_connection.export
		input  wire        clk_clk,                                                      //                                       clk.clk
		input  wire        hps_0_f2h_cold_reset_req_reset_n,                             //                  hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,                            //                 hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_dma_req0_dma_req,                                   //                        hps_0_f2h_dma_req0.dma_req
		input  wire        hps_0_f2h_dma_req0_dma_single,                                //                                          .dma_single
		output wire        hps_0_f2h_dma_req0_dma_ack,                                   //                                          .dma_ack
		input  wire        hps_0_f2h_dma_req1_dma_req,                                   //                        hps_0_f2h_dma_req1.dma_req
		input  wire        hps_0_f2h_dma_req1_dma_single,                                //                                          .dma_single
		output wire        hps_0_f2h_dma_req1_dma_ack,                                   //                                          .dma_ack
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,                         //                   hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,                             //                  hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,                                      //                           hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,                        //                              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,                          //                                          .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,                          //                                          .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,                          //                                          .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,                          //                                          .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,                          //                                          .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,                          //                                          .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,                           //                                          .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,                        //                                          .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,                        //                                          .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,                        //                                          .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,                          //                                          .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,                          //                                          .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,                          //                                          .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,                            //                                          .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,                            //                                          .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,                            //                                          .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,                            //                                          .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,                            //                                          .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,                            //                                          .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,                            //                                          .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,                             //                                          .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,                             //                                          .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,                            //                                          .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,                             //                                          .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,                             //                                          .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,                             //                                          .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,                             //                                          .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,                             //                                          .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,                             //                                          .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,                             //                                          .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,                             //                                          .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,                             //                                          .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,                             //                                          .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,                            //                                          .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,                            //                                          .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,                            //                                          .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,                            //                                          .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim0_inst_CLK,                           //                                          .hps_io_spim0_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim0_inst_MOSI,                          //                                          .hps_io_spim0_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim0_inst_MISO,                          //                                          .hps_io_spim0_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim0_inst_SS0,                           //                                          .hps_io_spim0_inst_SS0
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,                           //                                          .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,                          //                                          .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,                          //                                          .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,                           //                                          .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,                            //                                          .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,                            //                                          .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,                            //                                          .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,                            //                                          .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,                            //                                          .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,                            //                                          .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,                         //                                          .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,                         //                                          .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO37,                         //                                          .hps_io_gpio_inst_GPIO37
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,                         //                                          .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO41,                         //                                          .hps_io_gpio_inst_GPIO41
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO44,                         //                                          .hps_io_gpio_inst_GPIO44
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,                         //                                          .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,                         //                                          .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,                         //                                          .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,                         //                                          .hps_io_gpio_inst_GPIO61
		inout  wire        i2c_opencores_camera_export_scl_pad_io,                       //               i2c_opencores_camera_export.scl_pad_io
		inout  wire        i2c_opencores_camera_export_sda_pad_io,                       //                                          .sda_pad_io
		inout  wire        i2c_opencores_light_export_scl_pad_io,                        //                i2c_opencores_light_export.scl_pad_io
		inout  wire        i2c_opencores_light_export_sda_pad_io,                        //                                          .sda_pad_io
		inout  wire        i2c_opencores_mipi_export_scl_pad_io,                         //                 i2c_opencores_mipi_export.scl_pad_io
		inout  wire        i2c_opencores_mipi_export_sda_pad_io,                         //                                          .sda_pad_io
		input  wire        ir_rx_conduit_end_export,                                     //                         ir_rx_conduit_end.export
		input  wire [3:0]  key_external_connection_export,                               //                   key_external_connection.export
		output wire [9:0]  ledr_external_connection_export,                              //                  ledr_external_connection.export
		input  wire        light_int_external_connection_export,                         //             light_int_external_connection.export
		output wire [14:0] memory_mem_a,                                                 //                                    memory.mem_a
		output wire [2:0]  memory_mem_ba,                                                //                                          .mem_ba
		output wire        memory_mem_ck,                                                //                                          .mem_ck
		output wire        memory_mem_ck_n,                                              //                                          .mem_ck_n
		output wire        memory_mem_cke,                                               //                                          .mem_cke
		output wire        memory_mem_cs_n,                                              //                                          .mem_cs_n
		output wire        memory_mem_ras_n,                                             //                                          .mem_ras_n
		output wire        memory_mem_cas_n,                                             //                                          .mem_cas_n
		output wire        memory_mem_we_n,                                              //                                          .mem_we_n
		output wire        memory_mem_reset_n,                                           //                                          .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                                //                                          .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                               //                                          .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                             //                                          .mem_dqs_n
		output wire        memory_mem_odt,                                               //                                          .mem_odt
		output wire [3:0]  memory_mem_dm,                                                //                                          .mem_dm
		input  wire        memory_oct_rzqin,                                             //                                          .oct_rzqin
		output wire        mipi_reset_n_external_connection_export,                      //          mipi_reset_n_external_connection.export
		input  wire        mpu_int_external_connection_export,                           //               mpu_int_external_connection.export
		input  wire        reset_reset_n,                                                //                                     reset.reset_n
		output wire [47:0] seg7_conduit_end_writedata,                                   //                          seg7_conduit_end.writedata
		input  wire        spi_external_MISO,                                            //                              spi_external.MISO
		output wire        spi_external_MOSI,                                            //                                          .MOSI
		output wire        spi_external_SCLK,                                            //                                          .SCLK
		output wire        spi_external_SS_n,                                            //                                          .SS_n
		input  wire        spi_mpu_external_MISO,                                        //                          spi_mpu_external.MISO
		output wire        spi_mpu_external_MOSI,                                        //                                          .MOSI
		output wire        spi_mpu_external_SCLK,                                        //                                          .SCLK
		output wire        spi_mpu_external_SS_n,                                        //                                          .SS_n
		input  wire [9:0]  sw_external_connection_export,                                //                    sw_external_connection.export
		output wire        terasic_alsa_chip_conduit_end_xck,                            //             terasic_alsa_chip_conduit_end.xck
		inout  wire        terasic_alsa_chip_conduit_end_adclrck,                        //                                          .adclrck
		input  wire        terasic_alsa_chip_conduit_end_adcdat,                         //                                          .adcdat
		inout  wire        terasic_alsa_chip_conduit_end_bclk,                           //                                          .bclk
		output wire        terasic_alsa_chip_conduit_end_dacdat,                         //                                          .dacdat
		inout  wire        terasic_alsa_chip_conduit_end_daclrck,                        //                                          .daclrck
		input  wire        terasic_alsa_clock_sink_44_clk,                               //                terasic_alsa_clock_sink_44.clk
		input  wire        terasic_alsa_clock_sink_48_clk,                               //                terasic_alsa_clock_sink_48.clk
		input  wire        terasic_alsa_dma_conduit_end_capture_dma_ack,                 //              terasic_alsa_dma_conduit_end.capture_dma_ack
		output wire        terasic_alsa_dma_conduit_end_capture_dma_req,                 //                                          .capture_dma_req
		input  wire        terasic_alsa_dma_conduit_end_playback_dma_ack,                //                                          .playback_dma_ack
		output wire        terasic_alsa_dma_conduit_end_playback_dma_req,                //                                          .playback_dma_req
		inout  wire        ts_i2c_export_scl_pad_io,                                     //                             ts_i2c_export.scl_pad_io
		inout  wire        ts_i2c_export_sda_pad_io,                                     //                                          .sda_pad_io
		input  wire        ts_interrupt_external_connection_export,                      //          ts_interrupt_external_connection.export
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_clk,            // tv_decoder_alt_vip_cl_cvi_0_clocked_video.vid_clk
		input  wire [7:0]  tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_data,           //                                          .vid_data
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_de,             //                                          .vid_de
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_datavalid,      //                                          .vid_datavalid
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_locked,         //                                          .vid_locked
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_f,              //                                          .vid_f
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_v_sync,         //                                          .vid_v_sync
		input  wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_h_sync,         //                                          .vid_h_sync
		input  wire [7:0]  tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_color_encoding, //                                          .vid_color_encoding
		input  wire [7:0]  tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_bit_width,      //                                          .vid_bit_width
		output wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_sof,                //                                          .sof
		output wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_sof_locked,         //                                          .sof_locked
		output wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_refclk_div,         //                                          .refclk_div
		output wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_clipping,           //                                          .clipping
		output wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_padding,            //                                          .padding
		output wire        tv_decoder_alt_vip_cl_cvi_0_clocked_video_overflow,           //                                          .overflow
		input  wire [11:0] tv_decoder_camera_conduit_end_camera_d,                       //             tv_decoder_camera_conduit_end.camera_d
		input  wire        tv_decoder_camera_conduit_end_camera_fval,                    //                                          .camera_fval
		input  wire        tv_decoder_camera_conduit_end_camera_lval,                    //                                          .camera_lval
		input  wire        tv_decoder_camera_conduit_end_camera_pixclk,                  //                                          .camera_pixclk
		output wire [12:0] tv_decoder_sdram_wire_addr,                                   //                     tv_decoder_sdram_wire.addr
		output wire [1:0]  tv_decoder_sdram_wire_ba,                                     //                                          .ba
		output wire        tv_decoder_sdram_wire_cas_n,                                  //                                          .cas_n
		output wire        tv_decoder_sdram_wire_cke,                                    //                                          .cke
		output wire        tv_decoder_sdram_wire_cs_n,                                   //                                          .cs_n
		inout  wire [15:0] tv_decoder_sdram_wire_dq,                                     //                                          .dq
		output wire [1:0]  tv_decoder_sdram_wire_dqm,                                    //                                          .dqm
		output wire        tv_decoder_sdram_wire_ras_n,                                  //                                          .ras_n
		output wire        tv_decoder_sdram_wire_we_n,                                   //                                          .we_n
		input  wire        vga_stream_clk                                                //                                vga_stream.clk
	);

	wire          tv_decoder_alt_vip_cl_vfb_0_dout_valid;                              // tv_decoder:alt_vip_cl_vfb_0_dout_valid -> alt_vip_cl_mixer_0:din1_valid
	wire   [23:0] tv_decoder_alt_vip_cl_vfb_0_dout_data;                               // tv_decoder:alt_vip_cl_vfb_0_dout_data -> alt_vip_cl_mixer_0:din1_data
	wire          tv_decoder_alt_vip_cl_vfb_0_dout_ready;                              // alt_vip_cl_mixer_0:din1_ready -> tv_decoder:alt_vip_cl_vfb_0_dout_ready
	wire          tv_decoder_alt_vip_cl_vfb_0_dout_startofpacket;                      // tv_decoder:alt_vip_cl_vfb_0_dout_startofpacket -> alt_vip_cl_mixer_0:din1_startofpacket
	wire          tv_decoder_alt_vip_cl_vfb_0_dout_endofpacket;                        // tv_decoder:alt_vip_cl_vfb_0_dout_endofpacket -> alt_vip_cl_mixer_0:din1_endofpacket
	wire          alt_vip_vfr_vga_avalon_streaming_source_valid;                       // alt_vip_vfr_vga:dout_valid -> alt_vip_cl_cps_0:din_0_valid
	wire   [31:0] alt_vip_vfr_vga_avalon_streaming_source_data;                        // alt_vip_vfr_vga:dout_data -> alt_vip_cl_cps_0:din_0_data
	wire          alt_vip_vfr_vga_avalon_streaming_source_ready;                       // alt_vip_cl_cps_0:din_0_ready -> alt_vip_vfr_vga:dout_ready
	wire          alt_vip_vfr_vga_avalon_streaming_source_startofpacket;               // alt_vip_vfr_vga:dout_startofpacket -> alt_vip_cl_cps_0:din_0_startofpacket
	wire          alt_vip_vfr_vga_avalon_streaming_source_endofpacket;                 // alt_vip_vfr_vga:dout_endofpacket -> alt_vip_cl_cps_0:din_0_endofpacket
	wire          alt_vip_cl_mixer_0_dout_valid;                                       // alt_vip_cl_mixer_0:dout_valid -> alt_vip_itc_0:is_valid
	wire   [23:0] alt_vip_cl_mixer_0_dout_data;                                        // alt_vip_cl_mixer_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_cl_mixer_0_dout_ready;                                       // alt_vip_itc_0:is_ready -> alt_vip_cl_mixer_0:dout_ready
	wire          alt_vip_cl_mixer_0_dout_startofpacket;                               // alt_vip_cl_mixer_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_cl_mixer_0_dout_endofpacket;                                 // alt_vip_cl_mixer_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          alt_vip_cl_cps_0_dout_0_valid;                                       // alt_vip_cl_cps_0:dout_0_valid -> alt_vip_cl_mixer_0:din0_valid
	wire   [23:0] alt_vip_cl_cps_0_dout_0_data;                                        // alt_vip_cl_cps_0:dout_0_data -> alt_vip_cl_mixer_0:din0_data
	wire          alt_vip_cl_cps_0_dout_0_ready;                                       // alt_vip_cl_mixer_0:din0_ready -> alt_vip_cl_cps_0:dout_0_ready
	wire          alt_vip_cl_cps_0_dout_0_startofpacket;                               // alt_vip_cl_cps_0:dout_0_startofpacket -> alt_vip_cl_mixer_0:din0_startofpacket
	wire          alt_vip_cl_cps_0_dout_0_endofpacket;                                 // alt_vip_cl_cps_0:dout_0_endofpacket -> alt_vip_cl_mixer_0:din0_endofpacket
	wire  [127:0] alt_vip_vfr_vga_avalon_master_readdata;                              // mm_interconnect_0:alt_vip_vfr_vga_avalon_master_readdata -> alt_vip_vfr_vga:master_readdata
	wire          alt_vip_vfr_vga_avalon_master_waitrequest;                           // mm_interconnect_0:alt_vip_vfr_vga_avalon_master_waitrequest -> alt_vip_vfr_vga:master_waitrequest
	wire   [31:0] alt_vip_vfr_vga_avalon_master_address;                               // alt_vip_vfr_vga:master_address -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_address
	wire          alt_vip_vfr_vga_avalon_master_read;                                  // alt_vip_vfr_vga:master_read -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_read
	wire          alt_vip_vfr_vga_avalon_master_readdatavalid;                         // mm_interconnect_0:alt_vip_vfr_vga_avalon_master_readdatavalid -> alt_vip_vfr_vga:master_readdatavalid
	wire    [5:0] alt_vip_vfr_vga_avalon_master_burstcount;                            // alt_vip_vfr_vga:master_burstcount -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_burstcount
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;                        // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;                         // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;                         // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wready;                        // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;                           // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rready;                        // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;                         // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;                           // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;                        // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;                        // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;                        // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;                        // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;                         // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;                          // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;                        // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;                        // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;                        // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;                         // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arready;                       // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;                         // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awready;                       // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;                        // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bready;                        // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rlast;                         // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wlast;                         // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;                         // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;                          // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;                           // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;                        // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;                        // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;                        // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;                        // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire   [31:0] nios2_gen2_data_master_readdata;                                     // mm_interconnect_1:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire          nios2_gen2_data_master_waitrequest;                                  // mm_interconnect_1:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire          nios2_gen2_data_master_debugaccess;                                  // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_data_master_debugaccess
	wire   [18:0] nios2_gen2_data_master_address;                                      // nios2_gen2:d_address -> mm_interconnect_1:nios2_gen2_data_master_address
	wire    [3:0] nios2_gen2_data_master_byteenable;                                   // nios2_gen2:d_byteenable -> mm_interconnect_1:nios2_gen2_data_master_byteenable
	wire          nios2_gen2_data_master_read;                                         // nios2_gen2:d_read -> mm_interconnect_1:nios2_gen2_data_master_read
	wire          nios2_gen2_data_master_readdatavalid;                                // mm_interconnect_1:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire          nios2_gen2_data_master_write;                                        // nios2_gen2:d_write -> mm_interconnect_1:nios2_gen2_data_master_write
	wire   [31:0] nios2_gen2_data_master_writedata;                                    // nios2_gen2:d_writedata -> mm_interconnect_1:nios2_gen2_data_master_writedata
	wire          mm_bridge_0_m0_waitrequest;                                          // mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [31:0] mm_bridge_0_m0_readdata;                                             // mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                          // mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	wire   [18:0] mm_bridge_0_m0_address;                                              // mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	wire          mm_bridge_0_m0_read;                                                 // mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	wire    [3:0] mm_bridge_0_m0_byteenable;                                           // mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                                        // mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [31:0] mm_bridge_0_m0_writedata;                                            // mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                                // mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	wire    [0:0] mm_bridge_0_m0_burstcount;                                           // mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	wire   [31:0] nios2_gen2_instruction_master_readdata;                              // mm_interconnect_1:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire          nios2_gen2_instruction_master_waitrequest;                           // mm_interconnect_1:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire   [17:0] nios2_gen2_instruction_master_address;                               // nios2_gen2:i_address -> mm_interconnect_1:nios2_gen2_instruction_master_address
	wire          nios2_gen2_instruction_master_read;                                  // nios2_gen2:i_read -> mm_interconnect_1:nios2_gen2_instruction_master_read
	wire          nios2_gen2_instruction_master_readdatavalid;                         // mm_interconnect_1:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_readdata;      // tv_decoder:alt_vip_cl_cvi_0_control_readdata -> mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_readdata
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_waitrequest;   // tv_decoder:alt_vip_cl_cvi_0_control_waitrequest -> mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_waitrequest
	wire    [4:0] mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_address;       // mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_address -> tv_decoder:alt_vip_cl_cvi_0_control_address
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_read;          // mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_read -> tv_decoder:alt_vip_cl_cvi_0_control_read
	wire    [3:0] mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_byteenable;    // mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_byteenable -> tv_decoder:alt_vip_cl_cvi_0_control_byteenable
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_write;         // mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_write -> tv_decoder:alt_vip_cl_cvi_0_control_write
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_writedata;     // mm_interconnect_1:tv_decoder_alt_vip_cl_cvi_0_control_writedata -> tv_decoder:alt_vip_cl_cvi_0_control_writedata
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_readdata;      // tv_decoder:alt_vip_cl_scl_0_control_readdata -> mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_readdata
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_waitrequest;   // tv_decoder:alt_vip_cl_scl_0_control_waitrequest -> mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_waitrequest
	wire    [6:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_address;       // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_address -> tv_decoder:alt_vip_cl_scl_0_control_address
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_read;          // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_read -> tv_decoder:alt_vip_cl_scl_0_control_read
	wire    [3:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_byteenable;    // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_byteenable -> tv_decoder:alt_vip_cl_scl_0_control_byteenable
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_readdatavalid; // tv_decoder:alt_vip_cl_scl_0_control_readdatavalid -> mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_readdatavalid
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_write;         // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_write -> tv_decoder:alt_vip_cl_scl_0_control_write
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_writedata;     // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_0_control_writedata -> tv_decoder:alt_vip_cl_scl_0_control_writedata
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_readdata;      // tv_decoder:alt_vip_cl_scl_1_control_readdata -> mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_readdata
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_waitrequest;   // tv_decoder:alt_vip_cl_scl_1_control_waitrequest -> mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_waitrequest
	wire    [6:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_address;       // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_address -> tv_decoder:alt_vip_cl_scl_1_control_address
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_read;          // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_read -> tv_decoder:alt_vip_cl_scl_1_control_read
	wire    [3:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_byteenable;    // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_byteenable -> tv_decoder:alt_vip_cl_scl_1_control_byteenable
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_readdatavalid; // tv_decoder:alt_vip_cl_scl_1_control_readdatavalid -> mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_readdatavalid
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_write;         // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_write -> tv_decoder:alt_vip_cl_scl_1_control_write
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_writedata;     // mm_interconnect_1:tv_decoder_alt_vip_cl_scl_1_control_writedata -> tv_decoder:alt_vip_cl_scl_1_control_writedata
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_readdata;      // tv_decoder:alt_vip_cl_swi_0_control_readdata -> mm_interconnect_1:tv_decoder_alt_vip_cl_swi_0_control_readdata
	wire    [4:0] mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_address;       // mm_interconnect_1:tv_decoder_alt_vip_cl_swi_0_control_address -> tv_decoder:alt_vip_cl_swi_0_control_address
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_read;          // mm_interconnect_1:tv_decoder_alt_vip_cl_swi_0_control_read -> tv_decoder:alt_vip_cl_swi_0_control_read
	wire          mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_write;         // mm_interconnect_1:tv_decoder_alt_vip_cl_swi_0_control_write -> tv_decoder:alt_vip_cl_swi_0_control_write
	wire   [31:0] mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_writedata;     // mm_interconnect_1:tv_decoder_alt_vip_cl_swi_0_control_writedata -> tv_decoder:alt_vip_cl_swi_0_control_writedata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;              // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;           // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;               // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                 // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;             // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire          mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_chipselect;      // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_chipselect -> i2c_opencores_mipi:wb_stb_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_readdata;        // i2c_opencores_mipi:wb_dat_o -> mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_readdata
	wire          mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_waitrequest;     // i2c_opencores_mipi:wb_ack_o -> mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_address;         // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_address -> i2c_opencores_mipi:wb_adr_i
	wire          mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_write;           // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_write -> i2c_opencores_mipi:wb_we_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_writedata;       // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_writedata -> i2c_opencores_mipi:wb_dat_i
	wire          mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_chipselect;    // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_chipselect -> i2c_opencores_camera:wb_stb_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_readdata;      // i2c_opencores_camera:wb_dat_o -> mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_readdata
	wire          mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_waitrequest;   // i2c_opencores_camera:wb_ack_o -> mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_address;       // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_address -> i2c_opencores_camera:wb_adr_i
	wire          mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_write;         // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_write -> i2c_opencores_camera:wb_we_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_writedata;     // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_writedata -> i2c_opencores_camera:wb_dat_i
	wire   [31:0] mm_interconnect_1_alt_vip_cl_mixer_0_control_readdata;               // alt_vip_cl_mixer_0:control_readdata -> mm_interconnect_1:alt_vip_cl_mixer_0_control_readdata
	wire          mm_interconnect_1_alt_vip_cl_mixer_0_control_waitrequest;            // alt_vip_cl_mixer_0:control_waitrequest -> mm_interconnect_1:alt_vip_cl_mixer_0_control_waitrequest
	wire    [6:0] mm_interconnect_1_alt_vip_cl_mixer_0_control_address;                // mm_interconnect_1:alt_vip_cl_mixer_0_control_address -> alt_vip_cl_mixer_0:control_address
	wire          mm_interconnect_1_alt_vip_cl_mixer_0_control_read;                   // mm_interconnect_1:alt_vip_cl_mixer_0_control_read -> alt_vip_cl_mixer_0:control_read
	wire    [3:0] mm_interconnect_1_alt_vip_cl_mixer_0_control_byteenable;             // mm_interconnect_1:alt_vip_cl_mixer_0_control_byteenable -> alt_vip_cl_mixer_0:control_byteenable
	wire          mm_interconnect_1_alt_vip_cl_mixer_0_control_readdatavalid;          // alt_vip_cl_mixer_0:control_readdatavalid -> mm_interconnect_1:alt_vip_cl_mixer_0_control_readdatavalid
	wire          mm_interconnect_1_alt_vip_cl_mixer_0_control_write;                  // mm_interconnect_1:alt_vip_cl_mixer_0_control_write -> alt_vip_cl_mixer_0:control_write
	wire   [31:0] mm_interconnect_1_alt_vip_cl_mixer_0_control_writedata;              // mm_interconnect_1:alt_vip_cl_mixer_0_control_writedata -> alt_vip_cl_mixer_0:control_writedata
	wire   [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;                 // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;                  // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_1_nios2_gen2_debug_mem_slave_readdata;               // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_debug_mem_slave_readdata
	wire          mm_interconnect_1_nios2_gen2_debug_mem_slave_waitrequest;            // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_debug_mem_slave_waitrequest
	wire          mm_interconnect_1_nios2_gen2_debug_mem_slave_debugaccess;            // mm_interconnect_1:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_1_nios2_gen2_debug_mem_slave_address;                // mm_interconnect_1:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire          mm_interconnect_1_nios2_gen2_debug_mem_slave_read;                   // mm_interconnect_1:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire    [3:0] mm_interconnect_1_nios2_gen2_debug_mem_slave_byteenable;             // mm_interconnect_1:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire          mm_interconnect_1_nios2_gen2_debug_mem_slave_write;                  // mm_interconnect_1:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire   [31:0] mm_interconnect_1_nios2_gen2_debug_mem_slave_writedata;              // mm_interconnect_1:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire          mm_interconnect_1_onchip_memory2_s1_chipselect;                      // mm_interconnect_1:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire   [63:0] mm_interconnect_1_onchip_memory2_s1_readdata;                        // onchip_memory2:readdata -> mm_interconnect_1:onchip_memory2_s1_readdata
	wire   [12:0] mm_interconnect_1_onchip_memory2_s1_address;                         // mm_interconnect_1:onchip_memory2_s1_address -> onchip_memory2:address
	wire    [7:0] mm_interconnect_1_onchip_memory2_s1_byteenable;                      // mm_interconnect_1:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire          mm_interconnect_1_onchip_memory2_s1_write;                           // mm_interconnect_1:onchip_memory2_s1_write -> onchip_memory2:write
	wire   [63:0] mm_interconnect_1_onchip_memory2_s1_writedata;                       // mm_interconnect_1:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire          mm_interconnect_1_onchip_memory2_s1_clken;                           // mm_interconnect_1:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire          mm_interconnect_1_timer_s1_chipselect;                               // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire   [15:0] mm_interconnect_1_timer_s1_readdata;                                 // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire    [2:0] mm_interconnect_1_timer_s1_address;                                  // mm_interconnect_1:timer_s1_address -> timer:address
	wire          mm_interconnect_1_timer_s1_write;                                    // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire   [15:0] mm_interconnect_1_timer_s1_writedata;                                // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire          mm_interconnect_1_ledr_s1_chipselect;                                // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire   [31:0] mm_interconnect_1_ledr_s1_readdata;                                  // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire    [1:0] mm_interconnect_1_ledr_s1_address;                                   // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire          mm_interconnect_1_ledr_s1_write;                                     // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire   [31:0] mm_interconnect_1_ledr_s1_writedata;                                 // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire          mm_interconnect_1_camera_pwdn_n_s1_chipselect;                       // mm_interconnect_1:camera_pwdn_n_s1_chipselect -> camera_pwdn_n:chipselect
	wire   [31:0] mm_interconnect_1_camera_pwdn_n_s1_readdata;                         // camera_pwdn_n:readdata -> mm_interconnect_1:camera_pwdn_n_s1_readdata
	wire    [1:0] mm_interconnect_1_camera_pwdn_n_s1_address;                          // mm_interconnect_1:camera_pwdn_n_s1_address -> camera_pwdn_n:address
	wire          mm_interconnect_1_camera_pwdn_n_s1_write;                            // mm_interconnect_1:camera_pwdn_n_s1_write -> camera_pwdn_n:write_n
	wire   [31:0] mm_interconnect_1_camera_pwdn_n_s1_writedata;                        // mm_interconnect_1:camera_pwdn_n_s1_writedata -> camera_pwdn_n:writedata
	wire          mm_interconnect_1_mipi_reset_n_s1_chipselect;                        // mm_interconnect_1:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire   [31:0] mm_interconnect_1_mipi_reset_n_s1_readdata;                          // mipi_reset_n:readdata -> mm_interconnect_1:mipi_reset_n_s1_readdata
	wire    [1:0] mm_interconnect_1_mipi_reset_n_s1_address;                           // mm_interconnect_1:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire          mm_interconnect_1_mipi_reset_n_s1_write;                             // mm_interconnect_1:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire   [31:0] mm_interconnect_1_mipi_reset_n_s1_writedata;                         // mm_interconnect_1:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire    [4:0] mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_paddr;              // mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_paddr -> TERASIC_ALSA:clkctrl_paddr
	wire          mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pready;             // TERASIC_ALSA:clkctrl_pready -> mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_pready
	wire   [31:0] mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_prdata;             // TERASIC_ALSA:clkctrl_prdata -> mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_prdata
	wire   [31:0] mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pwdata;             // mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_pwdata -> TERASIC_ALSA:clkctrl_pwdata
	wire          mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_penable;            // mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_penable -> TERASIC_ALSA:clkctrl_penable
	wire          mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_psel;               // mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_psel -> TERASIC_ALSA:clkctrl_psel
	wire          mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pwrite;             // mm_interconnect_1:TERASIC_ALSA_apb_slave_clkctrl_pwrite -> TERASIC_ALSA:clkctrl_pwrite
	wire    [4:0] mm_interconnect_1_terasic_alsa_apb_slave_output_paddr;               // mm_interconnect_1:TERASIC_ALSA_apb_slave_output_paddr -> TERASIC_ALSA:output_paddr
	wire          mm_interconnect_1_terasic_alsa_apb_slave_output_pready;              // TERASIC_ALSA:output_pready -> mm_interconnect_1:TERASIC_ALSA_apb_slave_output_pready
	wire   [31:0] mm_interconnect_1_terasic_alsa_apb_slave_output_prdata;              // TERASIC_ALSA:output_prdata -> mm_interconnect_1:TERASIC_ALSA_apb_slave_output_prdata
	wire   [31:0] mm_interconnect_1_terasic_alsa_apb_slave_output_pwdata;              // mm_interconnect_1:TERASIC_ALSA_apb_slave_output_pwdata -> TERASIC_ALSA:output_pwdata
	wire          mm_interconnect_1_terasic_alsa_apb_slave_output_penable;             // mm_interconnect_1:TERASIC_ALSA_apb_slave_output_penable -> TERASIC_ALSA:output_penable
	wire          mm_interconnect_1_terasic_alsa_apb_slave_output_psel;                // mm_interconnect_1:TERASIC_ALSA_apb_slave_output_psel -> TERASIC_ALSA:output_psel
	wire          mm_interconnect_1_terasic_alsa_apb_slave_output_pwrite;              // mm_interconnect_1:TERASIC_ALSA_apb_slave_output_pwrite -> TERASIC_ALSA:output_pwrite
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata;             // alt_vip_vfr_vga:slave_readdata -> mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_readdata
	wire    [4:0] mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address;              // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_address -> alt_vip_vfr_vga:slave_address
	wire          mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read;                 // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_read -> alt_vip_vfr_vga:slave_read
	wire          mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write;                // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_write -> alt_vip_vfr_vga:slave_write
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata;            // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_writedata -> alt_vip_vfr_vga:slave_writedata
	wire          mm_interconnect_1_ir_rx_avalon_slave_chipselect;                     // mm_interconnect_1:ir_rx_avalon_slave_chipselect -> ir_rx:s_cs_n
	wire   [31:0] mm_interconnect_1_ir_rx_avalon_slave_readdata;                       // ir_rx:s_readdata -> mm_interconnect_1:ir_rx_avalon_slave_readdata
	wire    [0:0] mm_interconnect_1_ir_rx_avalon_slave_address;                        // mm_interconnect_1:ir_rx_avalon_slave_address -> ir_rx:s_address
	wire          mm_interconnect_1_ir_rx_avalon_slave_read;                           // mm_interconnect_1:ir_rx_avalon_slave_read -> ir_rx:s_read
	wire          mm_interconnect_1_ir_rx_avalon_slave_write;                          // mm_interconnect_1:ir_rx_avalon_slave_write -> ir_rx:s_write
	wire   [31:0] mm_interconnect_1_ir_rx_avalon_slave_writedata;                      // mm_interconnect_1:ir_rx_avalon_slave_writedata -> ir_rx:s_writedata
	wire          mm_interconnect_1_ts_i2c_avalon_slave_0_chipselect;                  // mm_interconnect_1:ts_i2c_avalon_slave_0_chipselect -> ts_i2c:wb_stb_i
	wire    [7:0] mm_interconnect_1_ts_i2c_avalon_slave_0_readdata;                    // ts_i2c:wb_dat_o -> mm_interconnect_1:ts_i2c_avalon_slave_0_readdata
	wire          mm_interconnect_1_ts_i2c_avalon_slave_0_waitrequest;                 // ts_i2c:wb_ack_o -> mm_interconnect_1:ts_i2c_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_1_ts_i2c_avalon_slave_0_address;                     // mm_interconnect_1:ts_i2c_avalon_slave_0_address -> ts_i2c:wb_adr_i
	wire          mm_interconnect_1_ts_i2c_avalon_slave_0_write;                       // mm_interconnect_1:ts_i2c_avalon_slave_0_write -> ts_i2c:wb_we_i
	wire    [7:0] mm_interconnect_1_ts_i2c_avalon_slave_0_writedata;                   // mm_interconnect_1:ts_i2c_avalon_slave_0_writedata -> ts_i2c:wb_dat_i
	wire          mm_interconnect_1_i2c_opencores_light_avalon_slave_0_chipselect;     // mm_interconnect_1:i2c_opencores_light_avalon_slave_0_chipselect -> i2c_opencores_light:wb_stb_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_light_avalon_slave_0_readdata;       // i2c_opencores_light:wb_dat_o -> mm_interconnect_1:i2c_opencores_light_avalon_slave_0_readdata
	wire          mm_interconnect_1_i2c_opencores_light_avalon_slave_0_waitrequest;    // i2c_opencores_light:wb_ack_o -> mm_interconnect_1:i2c_opencores_light_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_1_i2c_opencores_light_avalon_slave_0_address;        // mm_interconnect_1:i2c_opencores_light_avalon_slave_0_address -> i2c_opencores_light:wb_adr_i
	wire          mm_interconnect_1_i2c_opencores_light_avalon_slave_0_write;          // mm_interconnect_1:i2c_opencores_light_avalon_slave_0_write -> i2c_opencores_light:wb_we_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_light_avalon_slave_0_writedata;      // mm_interconnect_1:i2c_opencores_light_avalon_slave_0_writedata -> i2c_opencores_light:wb_dat_i
	wire          mm_interconnect_1_key_s1_chipselect;                                 // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire   [31:0] mm_interconnect_1_key_s1_readdata;                                   // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire    [1:0] mm_interconnect_1_key_s1_address;                                    // mm_interconnect_1:key_s1_address -> key:address
	wire          mm_interconnect_1_key_s1_write;                                      // mm_interconnect_1:key_s1_write -> key:write_n
	wire   [31:0] mm_interconnect_1_key_s1_writedata;                                  // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire          mm_interconnect_1_sw_s1_chipselect;                                  // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire   [31:0] mm_interconnect_1_sw_s1_readdata;                                    // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire    [1:0] mm_interconnect_1_sw_s1_address;                                     // mm_interconnect_1:sw_s1_address -> sw:address
	wire          mm_interconnect_1_sw_s1_write;                                       // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire   [31:0] mm_interconnect_1_sw_s1_writedata;                                   // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire          mm_interconnect_1_ts_interrupt_s1_chipselect;                        // mm_interconnect_1:ts_interrupt_s1_chipselect -> ts_interrupt:chipselect
	wire   [31:0] mm_interconnect_1_ts_interrupt_s1_readdata;                          // ts_interrupt:readdata -> mm_interconnect_1:ts_interrupt_s1_readdata
	wire    [1:0] mm_interconnect_1_ts_interrupt_s1_address;                           // mm_interconnect_1:ts_interrupt_s1_address -> ts_interrupt:address
	wire          mm_interconnect_1_ts_interrupt_s1_write;                             // mm_interconnect_1:ts_interrupt_s1_write -> ts_interrupt:write_n
	wire   [31:0] mm_interconnect_1_ts_interrupt_s1_writedata;                         // mm_interconnect_1:ts_interrupt_s1_writedata -> ts_interrupt:writedata
	wire          mm_interconnect_1_mpu_int_s1_chipselect;                             // mm_interconnect_1:mpu_int_s1_chipselect -> mpu_int:chipselect
	wire   [31:0] mm_interconnect_1_mpu_int_s1_readdata;                               // mpu_int:readdata -> mm_interconnect_1:mpu_int_s1_readdata
	wire    [1:0] mm_interconnect_1_mpu_int_s1_address;                                // mm_interconnect_1:mpu_int_s1_address -> mpu_int:address
	wire          mm_interconnect_1_mpu_int_s1_write;                                  // mm_interconnect_1:mpu_int_s1_write -> mpu_int:write_n
	wire   [31:0] mm_interconnect_1_mpu_int_s1_writedata;                              // mm_interconnect_1:mpu_int_s1_writedata -> mpu_int:writedata
	wire          mm_interconnect_1_light_int_s1_chipselect;                           // mm_interconnect_1:light_int_s1_chipselect -> light_int:chipselect
	wire   [31:0] mm_interconnect_1_light_int_s1_readdata;                             // light_int:readdata -> mm_interconnect_1:light_int_s1_readdata
	wire    [1:0] mm_interconnect_1_light_int_s1_address;                              // mm_interconnect_1:light_int_s1_address -> light_int:address
	wire          mm_interconnect_1_light_int_s1_write;                                // mm_interconnect_1:light_int_s1_write -> light_int:write_n
	wire   [31:0] mm_interconnect_1_light_int_s1_writedata;                            // mm_interconnect_1:light_int_s1_writedata -> light_int:writedata
	wire   [31:0] mm_interconnect_1_seg7_slave_readdata;                               // seg7:s_readdata -> mm_interconnect_1:seg7_slave_readdata
	wire    [2:0] mm_interconnect_1_seg7_slave_address;                                // mm_interconnect_1:seg7_slave_address -> seg7:s_address
	wire          mm_interconnect_1_seg7_slave_read;                                   // mm_interconnect_1:seg7_slave_read -> seg7:s_read
	wire          mm_interconnect_1_seg7_slave_write;                                  // mm_interconnect_1:seg7_slave_write -> seg7:s_write
	wire   [31:0] mm_interconnect_1_seg7_slave_writedata;                              // mm_interconnect_1:seg7_slave_writedata -> seg7:s_writedata
	wire          mm_interconnect_1_spi_spi_control_port_chipselect;                   // mm_interconnect_1:spi_spi_control_port_chipselect -> spi:spi_select
	wire   [15:0] mm_interconnect_1_spi_spi_control_port_readdata;                     // spi:data_to_cpu -> mm_interconnect_1:spi_spi_control_port_readdata
	wire    [2:0] mm_interconnect_1_spi_spi_control_port_address;                      // mm_interconnect_1:spi_spi_control_port_address -> spi:mem_addr
	wire          mm_interconnect_1_spi_spi_control_port_read;                         // mm_interconnect_1:spi_spi_control_port_read -> spi:read_n
	wire          mm_interconnect_1_spi_spi_control_port_write;                        // mm_interconnect_1:spi_spi_control_port_write -> spi:write_n
	wire   [15:0] mm_interconnect_1_spi_spi_control_port_writedata;                    // mm_interconnect_1:spi_spi_control_port_writedata -> spi:data_from_cpu
	wire          mm_interconnect_1_spi_mpu_spi_control_port_chipselect;               // mm_interconnect_1:spi_mpu_spi_control_port_chipselect -> spi_mpu:spi_select
	wire   [15:0] mm_interconnect_1_spi_mpu_spi_control_port_readdata;                 // spi_mpu:data_to_cpu -> mm_interconnect_1:spi_mpu_spi_control_port_readdata
	wire    [2:0] mm_interconnect_1_spi_mpu_spi_control_port_address;                  // mm_interconnect_1:spi_mpu_spi_control_port_address -> spi_mpu:mem_addr
	wire          mm_interconnect_1_spi_mpu_spi_control_port_read;                     // mm_interconnect_1:spi_mpu_spi_control_port_read -> spi_mpu:read_n
	wire          mm_interconnect_1_spi_mpu_spi_control_port_write;                    // mm_interconnect_1:spi_mpu_spi_control_port_write -> spi_mpu:write_n
	wire   [15:0] mm_interconnect_1_spi_mpu_spi_control_port_writedata;                // mm_interconnect_1:spi_mpu_spi_control_port_writedata -> spi_mpu:data_from_cpu
	wire          mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_chipselect; // mm_interconnect_1:tv_decoder_stream_capture_avalon_slave_chipselect -> tv_decoder:stream_capture_avalon_slave_chipselect_n
	wire   [31:0] mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_readdata;   // tv_decoder:stream_capture_avalon_slave_readdata -> mm_interconnect_1:tv_decoder_stream_capture_avalon_slave_readdata
	wire    [2:0] mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_address;    // mm_interconnect_1:tv_decoder_stream_capture_avalon_slave_address -> tv_decoder:stream_capture_avalon_slave_address
	wire          mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_read;       // mm_interconnect_1:tv_decoder_stream_capture_avalon_slave_read -> tv_decoder:stream_capture_avalon_slave_read
	wire          mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_write;      // mm_interconnect_1:tv_decoder_stream_capture_avalon_slave_write -> tv_decoder:stream_capture_avalon_slave_write
	wire   [31:0] mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_writedata;  // mm_interconnect_1:tv_decoder_stream_capture_avalon_slave_writedata -> tv_decoder:stream_capture_avalon_slave_writedata
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                     // hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                       // hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                       // hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                         // mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                      // hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                       // hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                         // hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                     // hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                      // hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                      // hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                      // hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                      // hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                       // hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                     // hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                     // hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                        // hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                      // hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                      // hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                      // hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                       // mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                     // mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                       // mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                     // mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                     // hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                      // hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                      // hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                       // mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                       // hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                       // mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                        // hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                         // mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                      // hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                     // hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_2_mm_bridge_0_s0_readdata;                           // mm_bridge_0:s0_readdata -> mm_interconnect_2:mm_bridge_0_s0_readdata
	wire          mm_interconnect_2_mm_bridge_0_s0_waitrequest;                        // mm_bridge_0:s0_waitrequest -> mm_interconnect_2:mm_bridge_0_s0_waitrequest
	wire          mm_interconnect_2_mm_bridge_0_s0_debugaccess;                        // mm_interconnect_2:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire   [18:0] mm_interconnect_2_mm_bridge_0_s0_address;                            // mm_interconnect_2:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire          mm_interconnect_2_mm_bridge_0_s0_read;                               // mm_interconnect_2:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire    [3:0] mm_interconnect_2_mm_bridge_0_s0_byteenable;                         // mm_interconnect_2:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire          mm_interconnect_2_mm_bridge_0_s0_readdatavalid;                      // mm_bridge_0:s0_readdatavalid -> mm_interconnect_2:mm_bridge_0_s0_readdatavalid
	wire          mm_interconnect_2_mm_bridge_0_s0_write;                              // mm_interconnect_2:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire   [31:0] mm_interconnect_2_mm_bridge_0_s0_writedata;                          // mm_interconnect_2:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire    [0:0] mm_interconnect_2_mm_bridge_0_s0_burstcount;                         // mm_interconnect_2:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire          tv_decoder_stream_capture_avalon_master_chipselect;                  // tv_decoder:stream_capture_avalon_master_chipselect_n -> mm_interconnect_3:tv_decoder_stream_capture_avalon_master_chipselect
	wire          tv_decoder_stream_capture_avalon_master_waitrequest;                 // mm_interconnect_3:tv_decoder_stream_capture_avalon_master_waitrequest -> tv_decoder:stream_capture_avalon_master_waitrequest_n
	wire   [31:0] tv_decoder_stream_capture_avalon_master_address;                     // tv_decoder:stream_capture_avalon_master_address -> mm_interconnect_3:tv_decoder_stream_capture_avalon_master_address
	wire          tv_decoder_stream_capture_avalon_master_write;                       // tv_decoder:stream_capture_avalon_master_write -> mm_interconnect_3:tv_decoder_stream_capture_avalon_master_write
	wire   [31:0] tv_decoder_stream_capture_avalon_master_writedata;                   // tv_decoder:stream_capture_avalon_master_writedata -> mm_interconnect_3:tv_decoder_stream_capture_avalon_master_writedata
	wire   [31:0] mm_interconnect_3_hps_0_f2h_sdram0_data_readdata;                    // hps_0:f2h_sdram0_READDATA -> mm_interconnect_3:hps_0_f2h_sdram0_data_readdata
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_waitrequest;                 // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_3:hps_0_f2h_sdram0_data_waitrequest
	wire   [29:0] mm_interconnect_3_hps_0_f2h_sdram0_data_address;                     // mm_interconnect_3:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_read;                        // mm_interconnect_3:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	wire    [3:0] mm_interconnect_3_hps_0_f2h_sdram0_data_byteenable;                  // mm_interconnect_3:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_readdatavalid;               // hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_3:hps_0_f2h_sdram0_data_readdatavalid
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_write;                       // mm_interconnect_3:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire   [31:0] mm_interconnect_3_hps_0_f2h_sdram0_data_writedata;                   // mm_interconnect_3:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_3_hps_0_f2h_sdram0_data_burstcount;                  // mm_interconnect_3:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire          irq_mapper_receiver0_irq;                                            // ts_i2c:wb_inta_o -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                            // i2c_opencores_camera:wb_inta_o -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                            // i2c_opencores_mipi:wb_inta_o -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                            // i2c_opencores_light:wb_inta_o -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                            // ts_interrupt:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                            // mpu_int:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                            // light_int:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                            // key:irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                            // sw:irq -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver9_irq;                                            // spi:irq -> irq_mapper:receiver9_irq
	wire          irq_mapper_receiver10_irq;                                           // spi_mpu:irq -> irq_mapper:receiver10_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                                  // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                  // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          irq_mapper_002_receiver0_irq;                                        // timer:irq -> irq_mapper_002:receiver0_irq
	wire          irq_mapper_002_receiver1_irq;                                        // jtag_uart:av_irq -> irq_mapper_002:receiver1_irq
	wire   [31:0] nios2_gen2_irq_irq;                                                  // irq_mapper_002:sender_irq -> nios2_gen2:irq
	wire          rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [TERASIC_ALSA:reset_n, alt_vip_vfr_vga:master_reset, camera_pwdn_n:reset_n, i2c_opencores_camera:wb_rst_i, i2c_opencores_light:wb_rst_i, i2c_opencores_mipi:wb_rst_i, ir_rx:reset_n, jtag_uart:rst_n, key:reset_n, ledr:reset_n, light_int:reset_n, mipi_reset_n:reset_n, mm_bridge_0:reset, mm_interconnect_0:alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mm_bridge_0_reset_reset_bridge_in_reset_reset, mpu_int:reset_n, onchip_memory2:reset, rst_translator:in_reset, seg7:s_reset, spi:reset_n, spi_mpu:reset_n, sw:reset_n, sysid_qsys:reset_n, timer:reset_n, ts_i2c:wb_rst_i, ts_interrupt:reset_n]
	wire          rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [alt_vip_cl_cps_0:main_reset, alt_vip_cl_mixer_0:main_reset_reset, alt_vip_itc_0:rst, alt_vip_vfr_vga:reset, mm_interconnect_1:alt_vip_cl_mixer_0_main_reset_reset_bridge_in_reset_reset, mm_interconnect_1:tv_decoder_clk_50_reset_reset_bridge_in_reset_reset, mm_interconnect_3:tv_decoder_clk_50_reset_reset_bridge_in_reset_reset, mm_interconnect_3:tv_decoder_stream_capture_avalon_master_translator_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                                  // rst_controller_002:reset_out -> [irq_mapper_002:reset, mm_interconnect_1:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n]
	wire          rst_controller_002_reset_out_reset_req;                              // rst_controller_002:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire          nios2_gen2_debug_reset_request_reset;                                // nios2_gen2:debug_reset_request -> rst_controller_002:reset_in0
	wire          rst_controller_003_reset_out_reset;                                  // rst_controller_003:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_004_reset_out_reset;                                  // rst_controller_004:reset_out -> mm_interconnect_3:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset

	TERASIC_ALSA terasic_alsa (
		.clk              (clk_clk),                                                  //             clock.clk
		.reset_n          (~rst_controller_reset_out_reset),                          //             reset.reset_n
		.AUD_XCK          (terasic_alsa_chip_conduit_end_xck),                        //  chip_conduit_end.xck
		.AUD_ADCLRCK      (terasic_alsa_chip_conduit_end_adclrck),                    //                  .adclrck
		.AUD_ADCDAT       (terasic_alsa_chip_conduit_end_adcdat),                     //                  .adcdat
		.AUD_BCLK         (terasic_alsa_chip_conduit_end_bclk),                       //                  .bclk
		.AUD_DACDAT       (terasic_alsa_chip_conduit_end_dacdat),                     //                  .dacdat
		.AUD_DACLRCK      (terasic_alsa_chip_conduit_end_daclrck),                    //                  .daclrck
		.output_paddr     (mm_interconnect_1_terasic_alsa_apb_slave_output_paddr),    //  apb_slave_output.paddr
		.output_penable   (mm_interconnect_1_terasic_alsa_apb_slave_output_penable),  //                  .penable
		.output_prdata    (mm_interconnect_1_terasic_alsa_apb_slave_output_prdata),   //                  .prdata
		.output_pready    (mm_interconnect_1_terasic_alsa_apb_slave_output_pready),   //                  .pready
		.output_psel      (mm_interconnect_1_terasic_alsa_apb_slave_output_psel),     //                  .psel
		.output_pwdata    (mm_interconnect_1_terasic_alsa_apb_slave_output_pwdata),   //                  .pwdata
		.output_pwrite    (mm_interconnect_1_terasic_alsa_apb_slave_output_pwrite),   //                  .pwrite
		.clkctrl_paddr    (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_paddr),   // apb_slave_clkctrl.paddr
		.clkctrl_penable  (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_penable), //                  .penable
		.clkctrl_prdata   (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_prdata),  //                  .prdata
		.clkctrl_pready   (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pready),  //                  .pready
		.clkctrl_psel     (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_psel),    //                  .psel
		.clkctrl_pwdata   (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pwdata),  //                  .pwdata
		.clkctrl_pwrite   (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pwrite),  //                  .pwrite
		.capture_dma_ack  (terasic_alsa_dma_conduit_end_capture_dma_ack),             //   dma_conduit_end.capture_dma_ack
		.capture_dma_req  (terasic_alsa_dma_conduit_end_capture_dma_req),             //                  .capture_dma_req
		.playback_dma_ack (terasic_alsa_dma_conduit_end_playback_dma_ack),            //                  .playback_dma_ack
		.playback_dma_req (terasic_alsa_dma_conduit_end_playback_dma_req),            //                  .playback_dma_req
		.clk_44           (terasic_alsa_clock_sink_44_clk),                           //     clock_sink_44.clk
		.clk_48           (terasic_alsa_clock_sink_48_clk)                            //     clock_sink_48.clk
	);

	soc_system_alt_vip_cl_cps_0 #(
		.BITS_PER_SYMBOL     (8),
		.USER_PACKET_SUPPORT ("PASSTHROUGH")
	) alt_vip_cl_cps_0 (
		.main_clock           (vga_stream_clk),                                        // main_clock.clk
		.main_reset           (rst_controller_001_reset_out_reset),                    // main_reset.reset
		.din_0_data           (alt_vip_vfr_vga_avalon_streaming_source_data),          //      din_0.data
		.din_0_valid          (alt_vip_vfr_vga_avalon_streaming_source_valid),         //           .valid
		.din_0_startofpacket  (alt_vip_vfr_vga_avalon_streaming_source_startofpacket), //           .startofpacket
		.din_0_endofpacket    (alt_vip_vfr_vga_avalon_streaming_source_endofpacket),   //           .endofpacket
		.din_0_ready          (alt_vip_vfr_vga_avalon_streaming_source_ready),         //           .ready
		.dout_0_data          (alt_vip_cl_cps_0_dout_0_data),                          //     dout_0.data
		.dout_0_valid         (alt_vip_cl_cps_0_dout_0_valid),                         //           .valid
		.dout_0_startofpacket (alt_vip_cl_cps_0_dout_0_startofpacket),                 //           .startofpacket
		.dout_0_endofpacket   (alt_vip_cl_cps_0_dout_0_endofpacket),                   //           .endofpacket
		.dout_0_ready         (alt_vip_cl_cps_0_dout_0_ready)                          //           .ready
	);

	soc_system_alt_vip_cl_mixer_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_WIDTH                    (800),
		.MAX_HEIGHT                   (480),
		.IS_422                       (1),
		.USER_PACKET_SUPPORT          ("PASSTHROUGH"),
		.USER_PACKET_FIFO_DEPTH       (0)
	) alt_vip_cl_mixer_0 (
		.main_clock_clk        (vga_stream_clk),                                             // main_clock.clk
		.main_reset_reset      (rst_controller_001_reset_out_reset),                         // main_reset.reset
		.din0_data             (alt_vip_cl_cps_0_dout_0_data),                               //       din0.data
		.din0_valid            (alt_vip_cl_cps_0_dout_0_valid),                              //           .valid
		.din0_startofpacket    (alt_vip_cl_cps_0_dout_0_startofpacket),                      //           .startofpacket
		.din0_endofpacket      (alt_vip_cl_cps_0_dout_0_endofpacket),                        //           .endofpacket
		.din0_ready            (alt_vip_cl_cps_0_dout_0_ready),                              //           .ready
		.din1_data             (tv_decoder_alt_vip_cl_vfb_0_dout_data),                      //       din1.data
		.din1_valid            (tv_decoder_alt_vip_cl_vfb_0_dout_valid),                     //           .valid
		.din1_startofpacket    (tv_decoder_alt_vip_cl_vfb_0_dout_startofpacket),             //           .startofpacket
		.din1_endofpacket      (tv_decoder_alt_vip_cl_vfb_0_dout_endofpacket),               //           .endofpacket
		.din1_ready            (tv_decoder_alt_vip_cl_vfb_0_dout_ready),                     //           .ready
		.dout_data             (alt_vip_cl_mixer_0_dout_data),                               //       dout.data
		.dout_valid            (alt_vip_cl_mixer_0_dout_valid),                              //           .valid
		.dout_startofpacket    (alt_vip_cl_mixer_0_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (alt_vip_cl_mixer_0_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (alt_vip_cl_mixer_0_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_1_alt_vip_cl_mixer_0_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_1_alt_vip_cl_mixer_0_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_1_alt_vip_cl_mixer_0_control_write),         //           .write
		.control_writedata     (mm_interconnect_1_alt_vip_cl_mixer_0_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_1_alt_vip_cl_mixer_0_control_read),          //           .read
		.control_readdata      (mm_interconnect_1_alt_vip_cl_mixer_0_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_1_alt_vip_cl_mixer_0_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_1_alt_vip_cl_mixer_0_control_waitrequest)    //           .waitrequest
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (800),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (8000),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (7999),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (30),
		.H_FRONT_PORCH                 (210),
		.H_BACK_PORCH                  (16),
		.V_SYNC_LENGTH                 (13),
		.V_FRONT_PORCH                 (22),
		.V_BACK_PORCH                  (10),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (vga_stream_clk),                            //       is_clk_rst.clk
		.rst           (rst_controller_001_reset_out_reset),        // is_clk_rst_reset.reset
		.is_data       (alt_vip_cl_mixer_0_dout_data),              //              din.data
		.is_valid      (alt_vip_cl_mixer_0_dout_valid),             //                 .valid
		.is_ready      (alt_vip_cl_mixer_0_dout_ready),             //                 .ready
		.is_sop        (alt_vip_cl_mixer_0_dout_startofpacket),     //                 .startofpacket
		.is_eop        (alt_vip_cl_mixer_0_dout_endofpacket),       //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (4),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (800),
		.MAX_IMAGE_HEIGHT               (480),
		.MEM_PORT_WIDTH                 (128),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_vga (
		.clock                (vga_stream_clk),                                           //             clock_reset.clk
		.reset                (rst_controller_001_reset_out_reset),                       //       clock_reset_reset.reset
		.master_clock         (clk_clk),                                                  //            clock_master.clk
		.master_reset         (rst_controller_reset_out_reset),                           //      clock_master_reset.reset
		.slave_address        (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                         //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_vga_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_vga_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_vga_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_vga_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_vga_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_vga_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_vga_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_vga_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_vga_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_vga_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_vga_avalon_master_waitrequest)                 //                        .waitrequest
	);

	soc_system_camera_pwdn_n camera_pwdn_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_1_camera_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_camera_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_camera_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_camera_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_camera_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (camera_pwdn_n_external_connection_export)       // external_connection.export
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),                      //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),                     // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),                      //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),                  //   f2h_stm_hw_events.stm_hwevents
		.f2h_dma_req0_req         (hps_0_f2h_dma_req0_dma_req),                            //        f2h_dma_req0.dma_req
		.f2h_dma_req0_single      (hps_0_f2h_dma_req0_dma_single),                         //                    .dma_single
		.f2h_dma_req0_ack         (hps_0_f2h_dma_req0_dma_ack),                            //                    .dma_ack
		.f2h_dma_req1_req         (hps_0_f2h_dma_req1_dma_req),                            //        f2h_dma_req1.dma_req
		.f2h_dma_req1_single      (hps_0_f2h_dma_req1_dma_single),                         //                    .dma_single
		.f2h_dma_req1_ack         (hps_0_f2h_dma_req1_dma_ack),                            //                    .dma_ack
		.mem_a                    (memory_mem_a),                                          //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                         //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                         //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                       //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                        //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                       //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                      //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                      //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                       //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                    //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                         //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                        //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                      //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                        //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                         //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                      //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),                 //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),                   //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),                   //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),                   //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),                   //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),                   //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),                   //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),                    //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),                 //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),                 //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),                 //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),                   //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),                   //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),                   //                    .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),                     //                    .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),                     //                    .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),                     //                    .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),                     //                    .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),                     //                    .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),                     //                    .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),                     //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                      //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                      //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),                     //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                      //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                      //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                      //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                      //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                      //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                      //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                      //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                      //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                      //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                      //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),                     //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),                     //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),                     //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),                     //                    .hps_io_usb1_inst_NXT
		.hps_io_spim0_inst_CLK    (hps_0_hps_io_hps_io_spim0_inst_CLK),                    //                    .hps_io_spim0_inst_CLK
		.hps_io_spim0_inst_MOSI   (hps_0_hps_io_hps_io_spim0_inst_MOSI),                   //                    .hps_io_spim0_inst_MOSI
		.hps_io_spim0_inst_MISO   (hps_0_hps_io_hps_io_spim0_inst_MISO),                   //                    .hps_io_spim0_inst_MISO
		.hps_io_spim0_inst_SS0    (hps_0_hps_io_hps_io_spim0_inst_SS0),                    //                    .hps_io_spim0_inst_SS0
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),                    //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),                   //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),                   //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),                    //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),                     //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),                     //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),                     //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),                     //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),                     //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),                     //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                  //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                  //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO37  (hps_0_hps_io_hps_io_gpio_inst_GPIO37),                  //                    .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                  //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_0_hps_io_hps_io_gpio_inst_GPIO41),                  //                    .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO44  (hps_0_hps_io_hps_io_gpio_inst_GPIO44),                  //                    .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),                  //                    .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                  //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                  //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                  //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                               //           h2f_reset.reset_n
		.f2h_sdram0_clk           (vga_stream_clk),                                        //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_3_hps_0_f2h_sdram0_data_address),       //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_3_hps_0_f2h_sdram0_data_burstcount),    //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_3_hps_0_f2h_sdram0_data_waitrequest),   //                    .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_3_hps_0_f2h_sdram0_data_readdata),      //                    .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_3_hps_0_f2h_sdram0_data_readdatavalid), //                    .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_3_hps_0_f2h_sdram0_data_read),          //                    .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_3_hps_0_f2h_sdram0_data_writedata),     //                    .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_3_hps_0_f2h_sdram0_data_byteenable),    //                    .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_3_hps_0_f2h_sdram0_data_write),         //                    .write
		.h2f_axi_clk              (clk_clk),                                               //       h2f_axi_clock.clk
		.h2f_AWID                 (),                                                      //      h2f_axi_master.awid
		.h2f_AWADDR               (),                                                      //                    .awaddr
		.h2f_AWLEN                (),                                                      //                    .awlen
		.h2f_AWSIZE               (),                                                      //                    .awsize
		.h2f_AWBURST              (),                                                      //                    .awburst
		.h2f_AWLOCK               (),                                                      //                    .awlock
		.h2f_AWCACHE              (),                                                      //                    .awcache
		.h2f_AWPROT               (),                                                      //                    .awprot
		.h2f_AWVALID              (),                                                      //                    .awvalid
		.h2f_AWREADY              (),                                                      //                    .awready
		.h2f_WID                  (),                                                      //                    .wid
		.h2f_WDATA                (),                                                      //                    .wdata
		.h2f_WSTRB                (),                                                      //                    .wstrb
		.h2f_WLAST                (),                                                      //                    .wlast
		.h2f_WVALID               (),                                                      //                    .wvalid
		.h2f_WREADY               (),                                                      //                    .wready
		.h2f_BID                  (),                                                      //                    .bid
		.h2f_BRESP                (),                                                      //                    .bresp
		.h2f_BVALID               (),                                                      //                    .bvalid
		.h2f_BREADY               (),                                                      //                    .bready
		.h2f_ARID                 (),                                                      //                    .arid
		.h2f_ARADDR               (),                                                      //                    .araddr
		.h2f_ARLEN                (),                                                      //                    .arlen
		.h2f_ARSIZE               (),                                                      //                    .arsize
		.h2f_ARBURST              (),                                                      //                    .arburst
		.h2f_ARLOCK               (),                                                      //                    .arlock
		.h2f_ARCACHE              (),                                                      //                    .arcache
		.h2f_ARPROT               (),                                                      //                    .arprot
		.h2f_ARVALID              (),                                                      //                    .arvalid
		.h2f_ARREADY              (),                                                      //                    .arready
		.h2f_RID                  (),                                                      //                    .rid
		.h2f_RDATA                (),                                                      //                    .rdata
		.h2f_RRESP                (),                                                      //                    .rresp
		.h2f_RLAST                (),                                                      //                    .rlast
		.h2f_RVALID               (),                                                      //                    .rvalid
		.h2f_RREADY               (),                                                      //                    .rready
		.f2h_axi_clk              (clk_clk),                                               //       f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_hps_0_f2h_axi_slave_awid),            //       f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),          //                    .awaddr
		.f2h_AWLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),           //                    .awlen
		.f2h_AWSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),          //                    .awsize
		.f2h_AWBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_awburst),         //                    .awburst
		.f2h_AWLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),          //                    .awlock
		.f2h_AWCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_awcache),         //                    .awcache
		.f2h_AWPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),          //                    .awprot
		.f2h_AWVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid),         //                    .awvalid
		.f2h_AWREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_awready),         //                    .awready
		.f2h_AWUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),          //                    .awuser
		.f2h_WID                  (mm_interconnect_0_hps_0_f2h_axi_slave_wid),             //                    .wid
		.f2h_WDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),           //                    .wdata
		.f2h_WSTRB                (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),           //                    .wstrb
		.f2h_WLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),           //                    .wlast
		.f2h_WVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),          //                    .wvalid
		.f2h_WREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_wready),          //                    .wready
		.f2h_BID                  (mm_interconnect_0_hps_0_f2h_axi_slave_bid),             //                    .bid
		.f2h_BRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),           //                    .bresp
		.f2h_BVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),          //                    .bvalid
		.f2h_BREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_bready),          //                    .bready
		.f2h_ARID                 (mm_interconnect_0_hps_0_f2h_axi_slave_arid),            //                    .arid
		.f2h_ARADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),          //                    .araddr
		.f2h_ARLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),           //                    .arlen
		.f2h_ARSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),          //                    .arsize
		.f2h_ARBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_arburst),         //                    .arburst
		.f2h_ARLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),          //                    .arlock
		.f2h_ARCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_arcache),         //                    .arcache
		.f2h_ARPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),          //                    .arprot
		.f2h_ARVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid),         //                    .arvalid
		.f2h_ARREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_arready),         //                    .arready
		.f2h_ARUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),          //                    .aruser
		.f2h_RID                  (mm_interconnect_0_hps_0_f2h_axi_slave_rid),             //                    .rid
		.f2h_RDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),           //                    .rdata
		.f2h_RRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),           //                    .rresp
		.f2h_RLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),           //                    .rlast
		.f2h_RVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),          //                    .rvalid
		.f2h_RREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_rready),          //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                                               //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                          //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                        //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                         //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                        //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                       //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                        //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                       //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                        //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                       //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                       //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                           //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                         //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                         //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                         //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                        //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                        //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                           //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                         //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                        //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                        //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                          //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                        //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                         //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                        //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                       //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                        //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                       //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                        //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                       //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                       //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                           //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                         //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                         //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                         //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                        //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                        //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                                    //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                                     //            f2h_irq1.irq
	);

	i2c_opencores i2c_opencores_camera (
		.wb_clk_i   (clk_clk),                                                           //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                    //      clock_reset.reset
		.scl_pad_io (i2c_opencores_camera_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_camera_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver1_irq)                                           // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_light (
		.wb_clk_i   (clk_clk),                                                          //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                   //      clock_reset.reset
		.scl_pad_io (i2c_opencores_light_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_light_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver3_irq)                                          // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_mipi (
		.wb_clk_i   (clk_clk),                                                         //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                  //      clock_reset.reset
		.scl_pad_io (i2c_opencores_mipi_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_mipi_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver2_irq)                                         // interrupt_sender.irq
	);

	TERASIC_IR_RX_FIFO ir_rx (
		.s_read      (mm_interconnect_1_ir_rx_avalon_slave_read),        //     avalon_slave.read
		.s_cs_n      (~mm_interconnect_1_ir_rx_avalon_slave_chipselect), //                 .chipselect_n
		.s_readdata  (mm_interconnect_1_ir_rx_avalon_slave_readdata),    //                 .readdata
		.s_write     (mm_interconnect_1_ir_rx_avalon_slave_write),       //                 .write
		.s_writedata (mm_interconnect_1_ir_rx_avalon_slave_writedata),   //                 .writedata
		.s_address   (mm_interconnect_1_ir_rx_avalon_slave_address),     //                 .address
		.clk         (clk_clk),                                          //       clock_sink.clk
		.reset_n     (~rst_controller_reset_out_reset),                  // clock_sink_reset.reset_n
		.ir          (ir_rx_conduit_end_export),                         //      conduit_end.export
		.irq         ()                                                  // interrupt_sender.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                               //               irq.irq
	);

	soc_system_key key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver7_irq)             //                 irq.irq
	);

	soc_system_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	soc_system_light_int light_int (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_light_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_light_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_light_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_light_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_light_int_s1_readdata),   //                    .readdata
		.in_port    (light_int_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                   //                 irq.irq
	);

	soc_system_camera_pwdn_n mipi_reset_n (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (19),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_2_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_2_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_2_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_2_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_2_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_2_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_2_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_2_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_2_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_2_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	soc_system_light_int mpu_int (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_mpu_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_mpu_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_mpu_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_mpu_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_mpu_int_s1_readdata),   //                    .readdata
		.in_port    (mpu_int_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                 //                 irq.irq
	);

	soc_system_nios2_gen2 nios2_gen2 (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	soc_system_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	TERASIC_SEG7 #(
		.SEG7_NUM       (6),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.SEG7        (seg7_conduit_end_writedata),             // conduit_end.writedata
		.s_clk       (clk_clk),                                //  clock_sink.clk
		.s_reset     (rst_controller_reset_out_reset),         //  reset_sink.reset
		.s_address   (mm_interconnect_1_seg7_slave_address),   //       slave.address
		.s_read      (mm_interconnect_1_seg7_slave_read),      //            .read
		.s_readdata  (mm_interconnect_1_seg7_slave_readdata),  //            .readdata
		.s_write     (mm_interconnect_1_seg7_slave_write),     //            .write
		.s_writedata (mm_interconnect_1_seg7_slave_writedata)  //            .writedata
	);

	soc_system_spi spi (
		.clk           (clk_clk),                                           //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver9_irq),                          //              irq.irq
		.MISO          (spi_external_MISO),                                 //         external.export
		.MOSI          (spi_external_MOSI),                                 //                 .export
		.SCLK          (spi_external_SCLK),                                 //                 .export
		.SS_n          (spi_external_SS_n)                                  //                 .export
	);

	soc_system_spi_mpu spi_mpu (
		.clk           (clk_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_spi_mpu_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_spi_mpu_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_spi_mpu_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_spi_mpu_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_spi_mpu_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_spi_mpu_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver10_irq),                             //              irq.irq
		.MISO          (spi_mpu_external_MISO),                                 //         external.export
		.MOSI          (spi_mpu_external_MOSI),                                 //                 .export
		.SCLK          (spi_mpu_external_SCLK),                                 //                 .export
		.SS_n          (spi_mpu_external_SS_n)                                  //                 .export
	);

	soc_system_sw sw (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver8_irq)            //                 irq.irq
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)           //   irq.irq
	);

	i2c_opencores ts_i2c (
		.wb_clk_i   (clk_clk),                                             //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                      //      clock_reset.reset
		.scl_pad_io (ts_i2c_export_scl_pad_io),                            //           export.export
		.sda_pad_io (ts_i2c_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_1_ts_i2c_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_ts_i2c_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_ts_i2c_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_ts_i2c_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_ts_i2c_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_ts_i2c_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                             // interrupt_sender.irq
	);

	soc_system_ts_interrupt ts_interrupt (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_ts_interrupt_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ts_interrupt_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ts_interrupt_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ts_interrupt_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ts_interrupt_s1_readdata),   //                    .readdata
		.in_port    (ts_interrupt_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                      //                 irq.irq
	);

	soc_system_tv_decoder tv_decoder (
		.alt_vip_cl_cvi_0_clocked_video_vid_clk            (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_clk),                    // alt_vip_cl_cvi_0_clocked_video.vid_clk
		.alt_vip_cl_cvi_0_clocked_video_vid_data           (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_data),                   //                               .vid_data
		.alt_vip_cl_cvi_0_clocked_video_vid_de             (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_de),                     //                               .vid_de
		.alt_vip_cl_cvi_0_clocked_video_vid_datavalid      (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_datavalid),              //                               .vid_datavalid
		.alt_vip_cl_cvi_0_clocked_video_vid_locked         (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_locked),                 //                               .vid_locked
		.alt_vip_cl_cvi_0_clocked_video_vid_f              (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_f),                      //                               .vid_f
		.alt_vip_cl_cvi_0_clocked_video_vid_v_sync         (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_v_sync),                 //                               .vid_v_sync
		.alt_vip_cl_cvi_0_clocked_video_vid_h_sync         (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_h_sync),                 //                               .vid_h_sync
		.alt_vip_cl_cvi_0_clocked_video_vid_color_encoding (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_color_encoding),         //                               .vid_color_encoding
		.alt_vip_cl_cvi_0_clocked_video_vid_bit_width      (tv_decoder_alt_vip_cl_cvi_0_clocked_video_vid_bit_width),              //                               .vid_bit_width
		.alt_vip_cl_cvi_0_clocked_video_sof                (tv_decoder_alt_vip_cl_cvi_0_clocked_video_sof),                        //                               .sof
		.alt_vip_cl_cvi_0_clocked_video_sof_locked         (tv_decoder_alt_vip_cl_cvi_0_clocked_video_sof_locked),                 //                               .sof_locked
		.alt_vip_cl_cvi_0_clocked_video_refclk_div         (tv_decoder_alt_vip_cl_cvi_0_clocked_video_refclk_div),                 //                               .refclk_div
		.alt_vip_cl_cvi_0_clocked_video_clipping           (tv_decoder_alt_vip_cl_cvi_0_clocked_video_clipping),                   //                               .clipping
		.alt_vip_cl_cvi_0_clocked_video_padding            (tv_decoder_alt_vip_cl_cvi_0_clocked_video_padding),                    //                               .padding
		.alt_vip_cl_cvi_0_clocked_video_overflow           (tv_decoder_alt_vip_cl_cvi_0_clocked_video_overflow),                   //                               .overflow
		.alt_vip_cl_cvi_0_control_address                  (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_address),        //       alt_vip_cl_cvi_0_control.address
		.alt_vip_cl_cvi_0_control_read                     (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_read),           //                               .read
		.alt_vip_cl_cvi_0_control_readdata                 (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_readdata),       //                               .readdata
		.alt_vip_cl_cvi_0_control_write                    (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_write),          //                               .write
		.alt_vip_cl_cvi_0_control_writedata                (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_writedata),      //                               .writedata
		.alt_vip_cl_cvi_0_control_byteenable               (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_byteenable),     //                               .byteenable
		.alt_vip_cl_cvi_0_control_waitrequest              (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_waitrequest),    //                               .waitrequest
		.alt_vip_cl_scl_0_control_address                  (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_address),        //       alt_vip_cl_scl_0_control.address
		.alt_vip_cl_scl_0_control_byteenable               (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_byteenable),     //                               .byteenable
		.alt_vip_cl_scl_0_control_write                    (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_write),          //                               .write
		.alt_vip_cl_scl_0_control_writedata                (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_writedata),      //                               .writedata
		.alt_vip_cl_scl_0_control_read                     (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_read),           //                               .read
		.alt_vip_cl_scl_0_control_readdata                 (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_readdata),       //                               .readdata
		.alt_vip_cl_scl_0_control_readdatavalid            (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_readdatavalid),  //                               .readdatavalid
		.alt_vip_cl_scl_0_control_waitrequest              (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_waitrequest),    //                               .waitrequest
		.alt_vip_cl_scl_1_control_address                  (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_address),        //       alt_vip_cl_scl_1_control.address
		.alt_vip_cl_scl_1_control_byteenable               (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_byteenable),     //                               .byteenable
		.alt_vip_cl_scl_1_control_write                    (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_write),          //                               .write
		.alt_vip_cl_scl_1_control_writedata                (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_writedata),      //                               .writedata
		.alt_vip_cl_scl_1_control_read                     (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_read),           //                               .read
		.alt_vip_cl_scl_1_control_readdata                 (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_readdata),       //                               .readdata
		.alt_vip_cl_scl_1_control_readdatavalid            (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_readdatavalid),  //                               .readdatavalid
		.alt_vip_cl_scl_1_control_waitrequest              (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_waitrequest),    //                               .waitrequest
		.alt_vip_cl_swi_0_control_read                     (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_read),           //       alt_vip_cl_swi_0_control.read
		.alt_vip_cl_swi_0_control_write                    (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_write),          //                               .write
		.alt_vip_cl_swi_0_control_address                  (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_address),        //                               .address
		.alt_vip_cl_swi_0_control_writedata                (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_writedata),      //                               .writedata
		.alt_vip_cl_swi_0_control_readdata                 (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_readdata),       //                               .readdata
		.alt_vip_cl_vfb_0_dout_data                        (tv_decoder_alt_vip_cl_vfb_0_dout_data),                                //          alt_vip_cl_vfb_0_dout.data
		.alt_vip_cl_vfb_0_dout_valid                       (tv_decoder_alt_vip_cl_vfb_0_dout_valid),                               //                               .valid
		.alt_vip_cl_vfb_0_dout_startofpacket               (tv_decoder_alt_vip_cl_vfb_0_dout_startofpacket),                       //                               .startofpacket
		.alt_vip_cl_vfb_0_dout_endofpacket                 (tv_decoder_alt_vip_cl_vfb_0_dout_endofpacket),                         //                               .endofpacket
		.alt_vip_cl_vfb_0_dout_ready                       (tv_decoder_alt_vip_cl_vfb_0_dout_ready),                               //                               .ready
		.camera_conduit_end_camera_d                       (tv_decoder_camera_conduit_end_camera_d),                               //             camera_conduit_end.camera_d
		.camera_conduit_end_camera_fval                    (tv_decoder_camera_conduit_end_camera_fval),                            //                               .camera_fval
		.camera_conduit_end_camera_lval                    (tv_decoder_camera_conduit_end_camera_lval),                            //                               .camera_lval
		.camera_conduit_end_camera_pixclk                  (tv_decoder_camera_conduit_end_camera_pixclk),                          //                               .camera_pixclk
		.clk_50_clk                                        (clk_clk),                                                              //                         clk_50.clk
		.clk_50_reset_reset_n                              (reset_reset_n),                                                        //                   clk_50_reset.reset_n
		.clk_vip_clk                                       (vga_stream_clk),                                                       //                        clk_vip.clk
		.zs_addr_from_the_sdram                            (tv_decoder_sdram_wire_addr),                                           //                     sdram_wire.addr
		.zs_ba_from_the_sdram                              (tv_decoder_sdram_wire_ba),                                             //                               .ba
		.zs_cas_n_from_the_sdram                           (tv_decoder_sdram_wire_cas_n),                                          //                               .cas_n
		.zs_cke_from_the_sdram                             (tv_decoder_sdram_wire_cke),                                            //                               .cke
		.zs_cs_n_from_the_sdram                            (tv_decoder_sdram_wire_cs_n),                                           //                               .cs_n
		.zs_dq_to_and_from_the_sdram                       (tv_decoder_sdram_wire_dq),                                             //                               .dq
		.zs_dqm_from_the_sdram                             (tv_decoder_sdram_wire_dqm),                                            //                               .dqm
		.zs_ras_n_from_the_sdram                           (tv_decoder_sdram_wire_ras_n),                                          //                               .ras_n
		.zs_we_n_from_the_sdram                            (tv_decoder_sdram_wire_we_n),                                           //                               .we_n
		.stream_capture_avalon_master_chipselect_n         (tv_decoder_stream_capture_avalon_master_chipselect),                   //   stream_capture_avalon_master.chipselect_n
		.stream_capture_avalon_master_address              (tv_decoder_stream_capture_avalon_master_address),                      //                               .address
		.stream_capture_avalon_master_write                (tv_decoder_stream_capture_avalon_master_write),                        //                               .write
		.stream_capture_avalon_master_writedata            (tv_decoder_stream_capture_avalon_master_writedata),                    //                               .writedata
		.stream_capture_avalon_master_waitrequest_n        (~tv_decoder_stream_capture_avalon_master_waitrequest),                 //                               .waitrequest_n
		.stream_capture_avalon_slave_read                  (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_read),        //    stream_capture_avalon_slave.read
		.stream_capture_avalon_slave_readdata              (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_readdata),    //                               .readdata
		.stream_capture_avalon_slave_write                 (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_write),       //                               .write
		.stream_capture_avalon_slave_writedata             (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_writedata),   //                               .writedata
		.stream_capture_avalon_slave_chipselect_n          (~mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_chipselect), //                               .chipselect_n
		.stream_capture_avalon_slave_address               (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_address)      //                               .address
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.clk_50_clk_clk                                                   (clk_clk),                                       //                                                 clk_50_clk.clk
		.alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                //   alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.alt_vip_vfr_vga_avalon_master_address                            (alt_vip_vfr_vga_avalon_master_address),         //                              alt_vip_vfr_vga_avalon_master.address
		.alt_vip_vfr_vga_avalon_master_waitrequest                        (alt_vip_vfr_vga_avalon_master_waitrequest),     //                                                           .waitrequest
		.alt_vip_vfr_vga_avalon_master_burstcount                         (alt_vip_vfr_vga_avalon_master_burstcount),      //                                                           .burstcount
		.alt_vip_vfr_vga_avalon_master_read                               (alt_vip_vfr_vga_avalon_master_read),            //                                                           .read
		.alt_vip_vfr_vga_avalon_master_readdata                           (alt_vip_vfr_vga_avalon_master_readdata),        //                                                           .readdata
		.alt_vip_vfr_vga_avalon_master_readdatavalid                      (alt_vip_vfr_vga_avalon_master_readdatavalid)    //                                                           .readdatavalid
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.TERASIC_ALSA_apb_slave_clkctrl_paddr                      (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_paddr),              //                      TERASIC_ALSA_apb_slave_clkctrl.paddr
		.TERASIC_ALSA_apb_slave_clkctrl_psel                       (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_psel),               //                                                    .psel
		.TERASIC_ALSA_apb_slave_clkctrl_penable                    (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_penable),            //                                                    .penable
		.TERASIC_ALSA_apb_slave_clkctrl_pwrite                     (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pwrite),             //                                                    .pwrite
		.TERASIC_ALSA_apb_slave_clkctrl_pwdata                     (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pwdata),             //                                                    .pwdata
		.TERASIC_ALSA_apb_slave_clkctrl_prdata                     (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_prdata),             //                                                    .prdata
		.TERASIC_ALSA_apb_slave_clkctrl_pready                     (mm_interconnect_1_terasic_alsa_apb_slave_clkctrl_pready),             //                                                    .pready
		.TERASIC_ALSA_apb_slave_output_paddr                       (mm_interconnect_1_terasic_alsa_apb_slave_output_paddr),               //                       TERASIC_ALSA_apb_slave_output.paddr
		.TERASIC_ALSA_apb_slave_output_psel                        (mm_interconnect_1_terasic_alsa_apb_slave_output_psel),                //                                                    .psel
		.TERASIC_ALSA_apb_slave_output_penable                     (mm_interconnect_1_terasic_alsa_apb_slave_output_penable),             //                                                    .penable
		.TERASIC_ALSA_apb_slave_output_pwrite                      (mm_interconnect_1_terasic_alsa_apb_slave_output_pwrite),              //                                                    .pwrite
		.TERASIC_ALSA_apb_slave_output_pwdata                      (mm_interconnect_1_terasic_alsa_apb_slave_output_pwdata),              //                                                    .pwdata
		.TERASIC_ALSA_apb_slave_output_prdata                      (mm_interconnect_1_terasic_alsa_apb_slave_output_prdata),              //                                                    .prdata
		.TERASIC_ALSA_apb_slave_output_pready                      (mm_interconnect_1_terasic_alsa_apb_slave_output_pready),              //                                                    .pready
		.clk_50_clk_clk                                            (clk_clk),                                                             //                                          clk_50_clk.clk
		.vga_stream_out_clk_clk                                    (vga_stream_clk),                                                      //                                  vga_stream_out_clk.clk
		.alt_vip_cl_mixer_0_main_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                  // alt_vip_cl_mixer_0_main_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                      //             mm_bridge_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset              (rst_controller_002_reset_out_reset),                                  //              nios2_gen2_reset_reset_bridge_in_reset.reset
		.tv_decoder_clk_50_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                                  //       tv_decoder_clk_50_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                                    (mm_bridge_0_m0_address),                                              //                                      mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                                (mm_bridge_0_m0_waitrequest),                                          //                                                    .waitrequest
		.mm_bridge_0_m0_burstcount                                 (mm_bridge_0_m0_burstcount),                                           //                                                    .burstcount
		.mm_bridge_0_m0_byteenable                                 (mm_bridge_0_m0_byteenable),                                           //                                                    .byteenable
		.mm_bridge_0_m0_read                                       (mm_bridge_0_m0_read),                                                 //                                                    .read
		.mm_bridge_0_m0_readdata                                   (mm_bridge_0_m0_readdata),                                             //                                                    .readdata
		.mm_bridge_0_m0_readdatavalid                              (mm_bridge_0_m0_readdatavalid),                                        //                                                    .readdatavalid
		.mm_bridge_0_m0_write                                      (mm_bridge_0_m0_write),                                                //                                                    .write
		.mm_bridge_0_m0_writedata                                  (mm_bridge_0_m0_writedata),                                            //                                                    .writedata
		.mm_bridge_0_m0_debugaccess                                (mm_bridge_0_m0_debugaccess),                                          //                                                    .debugaccess
		.nios2_gen2_data_master_address                            (nios2_gen2_data_master_address),                                      //                              nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                        (nios2_gen2_data_master_waitrequest),                                  //                                                    .waitrequest
		.nios2_gen2_data_master_byteenable                         (nios2_gen2_data_master_byteenable),                                   //                                                    .byteenable
		.nios2_gen2_data_master_read                               (nios2_gen2_data_master_read),                                         //                                                    .read
		.nios2_gen2_data_master_readdata                           (nios2_gen2_data_master_readdata),                                     //                                                    .readdata
		.nios2_gen2_data_master_readdatavalid                      (nios2_gen2_data_master_readdatavalid),                                //                                                    .readdatavalid
		.nios2_gen2_data_master_write                              (nios2_gen2_data_master_write),                                        //                                                    .write
		.nios2_gen2_data_master_writedata                          (nios2_gen2_data_master_writedata),                                    //                                                    .writedata
		.nios2_gen2_data_master_debugaccess                        (nios2_gen2_data_master_debugaccess),                                  //                                                    .debugaccess
		.nios2_gen2_instruction_master_address                     (nios2_gen2_instruction_master_address),                               //                       nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                 (nios2_gen2_instruction_master_waitrequest),                           //                                                    .waitrequest
		.nios2_gen2_instruction_master_read                        (nios2_gen2_instruction_master_read),                                  //                                                    .read
		.nios2_gen2_instruction_master_readdata                    (nios2_gen2_instruction_master_readdata),                              //                                                    .readdata
		.nios2_gen2_instruction_master_readdatavalid               (nios2_gen2_instruction_master_readdatavalid),                         //                                                    .readdatavalid
		.alt_vip_cl_mixer_0_control_address                        (mm_interconnect_1_alt_vip_cl_mixer_0_control_address),                //                          alt_vip_cl_mixer_0_control.address
		.alt_vip_cl_mixer_0_control_write                          (mm_interconnect_1_alt_vip_cl_mixer_0_control_write),                  //                                                    .write
		.alt_vip_cl_mixer_0_control_read                           (mm_interconnect_1_alt_vip_cl_mixer_0_control_read),                   //                                                    .read
		.alt_vip_cl_mixer_0_control_readdata                       (mm_interconnect_1_alt_vip_cl_mixer_0_control_readdata),               //                                                    .readdata
		.alt_vip_cl_mixer_0_control_writedata                      (mm_interconnect_1_alt_vip_cl_mixer_0_control_writedata),              //                                                    .writedata
		.alt_vip_cl_mixer_0_control_byteenable                     (mm_interconnect_1_alt_vip_cl_mixer_0_control_byteenable),             //                                                    .byteenable
		.alt_vip_cl_mixer_0_control_readdatavalid                  (mm_interconnect_1_alt_vip_cl_mixer_0_control_readdatavalid),          //                                                    .readdatavalid
		.alt_vip_cl_mixer_0_control_waitrequest                    (mm_interconnect_1_alt_vip_cl_mixer_0_control_waitrequest),            //                                                    .waitrequest
		.alt_vip_vfr_vga_avalon_slave_address                      (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address),              //                        alt_vip_vfr_vga_avalon_slave.address
		.alt_vip_vfr_vga_avalon_slave_write                        (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write),                //                                                    .write
		.alt_vip_vfr_vga_avalon_slave_read                         (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read),                 //                                                    .read
		.alt_vip_vfr_vga_avalon_slave_readdata                     (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata),             //                                                    .readdata
		.alt_vip_vfr_vga_avalon_slave_writedata                    (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata),            //                                                    .writedata
		.camera_pwdn_n_s1_address                                  (mm_interconnect_1_camera_pwdn_n_s1_address),                          //                                    camera_pwdn_n_s1.address
		.camera_pwdn_n_s1_write                                    (mm_interconnect_1_camera_pwdn_n_s1_write),                            //                                                    .write
		.camera_pwdn_n_s1_readdata                                 (mm_interconnect_1_camera_pwdn_n_s1_readdata),                         //                                                    .readdata
		.camera_pwdn_n_s1_writedata                                (mm_interconnect_1_camera_pwdn_n_s1_writedata),                        //                                                    .writedata
		.camera_pwdn_n_s1_chipselect                               (mm_interconnect_1_camera_pwdn_n_s1_chipselect),                       //                                                    .chipselect
		.i2c_opencores_camera_avalon_slave_0_address               (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_address),       //                 i2c_opencores_camera_avalon_slave_0.address
		.i2c_opencores_camera_avalon_slave_0_write                 (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_write),         //                                                    .write
		.i2c_opencores_camera_avalon_slave_0_readdata              (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_readdata),      //                                                    .readdata
		.i2c_opencores_camera_avalon_slave_0_writedata             (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_writedata),     //                                                    .writedata
		.i2c_opencores_camera_avalon_slave_0_waitrequest           (~mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_waitrequest),  //                                                    .waitrequest
		.i2c_opencores_camera_avalon_slave_0_chipselect            (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_chipselect),    //                                                    .chipselect
		.i2c_opencores_light_avalon_slave_0_address                (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_address),        //                  i2c_opencores_light_avalon_slave_0.address
		.i2c_opencores_light_avalon_slave_0_write                  (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_write),          //                                                    .write
		.i2c_opencores_light_avalon_slave_0_readdata               (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_readdata),       //                                                    .readdata
		.i2c_opencores_light_avalon_slave_0_writedata              (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_writedata),      //                                                    .writedata
		.i2c_opencores_light_avalon_slave_0_waitrequest            (~mm_interconnect_1_i2c_opencores_light_avalon_slave_0_waitrequest),   //                                                    .waitrequest
		.i2c_opencores_light_avalon_slave_0_chipselect             (mm_interconnect_1_i2c_opencores_light_avalon_slave_0_chipselect),     //                                                    .chipselect
		.i2c_opencores_mipi_avalon_slave_0_address                 (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_address),         //                   i2c_opencores_mipi_avalon_slave_0.address
		.i2c_opencores_mipi_avalon_slave_0_write                   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_write),           //                                                    .write
		.i2c_opencores_mipi_avalon_slave_0_readdata                (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_readdata),        //                                                    .readdata
		.i2c_opencores_mipi_avalon_slave_0_writedata               (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_writedata),       //                                                    .writedata
		.i2c_opencores_mipi_avalon_slave_0_waitrequest             (~mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_waitrequest),    //                                                    .waitrequest
		.i2c_opencores_mipi_avalon_slave_0_chipselect              (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_chipselect),      //                                                    .chipselect
		.ir_rx_avalon_slave_address                                (mm_interconnect_1_ir_rx_avalon_slave_address),                        //                                  ir_rx_avalon_slave.address
		.ir_rx_avalon_slave_write                                  (mm_interconnect_1_ir_rx_avalon_slave_write),                          //                                                    .write
		.ir_rx_avalon_slave_read                                   (mm_interconnect_1_ir_rx_avalon_slave_read),                           //                                                    .read
		.ir_rx_avalon_slave_readdata                               (mm_interconnect_1_ir_rx_avalon_slave_readdata),                       //                                                    .readdata
		.ir_rx_avalon_slave_writedata                              (mm_interconnect_1_ir_rx_avalon_slave_writedata),                      //                                                    .writedata
		.ir_rx_avalon_slave_chipselect                             (mm_interconnect_1_ir_rx_avalon_slave_chipselect),                     //                                                    .chipselect
		.jtag_uart_avalon_jtag_slave_address                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),               //                         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),                 //                                                    .write
		.jtag_uart_avalon_jtag_slave_read                          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),                  //                                                    .read
		.jtag_uart_avalon_jtag_slave_readdata                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),              //                                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),             //                                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),           //                                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),            //                                                    .chipselect
		.key_s1_address                                            (mm_interconnect_1_key_s1_address),                                    //                                              key_s1.address
		.key_s1_write                                              (mm_interconnect_1_key_s1_write),                                      //                                                    .write
		.key_s1_readdata                                           (mm_interconnect_1_key_s1_readdata),                                   //                                                    .readdata
		.key_s1_writedata                                          (mm_interconnect_1_key_s1_writedata),                                  //                                                    .writedata
		.key_s1_chipselect                                         (mm_interconnect_1_key_s1_chipselect),                                 //                                                    .chipselect
		.ledr_s1_address                                           (mm_interconnect_1_ledr_s1_address),                                   //                                             ledr_s1.address
		.ledr_s1_write                                             (mm_interconnect_1_ledr_s1_write),                                     //                                                    .write
		.ledr_s1_readdata                                          (mm_interconnect_1_ledr_s1_readdata),                                  //                                                    .readdata
		.ledr_s1_writedata                                         (mm_interconnect_1_ledr_s1_writedata),                                 //                                                    .writedata
		.ledr_s1_chipselect                                        (mm_interconnect_1_ledr_s1_chipselect),                                //                                                    .chipselect
		.light_int_s1_address                                      (mm_interconnect_1_light_int_s1_address),                              //                                        light_int_s1.address
		.light_int_s1_write                                        (mm_interconnect_1_light_int_s1_write),                                //                                                    .write
		.light_int_s1_readdata                                     (mm_interconnect_1_light_int_s1_readdata),                             //                                                    .readdata
		.light_int_s1_writedata                                    (mm_interconnect_1_light_int_s1_writedata),                            //                                                    .writedata
		.light_int_s1_chipselect                                   (mm_interconnect_1_light_int_s1_chipselect),                           //                                                    .chipselect
		.mipi_reset_n_s1_address                                   (mm_interconnect_1_mipi_reset_n_s1_address),                           //                                     mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                                     (mm_interconnect_1_mipi_reset_n_s1_write),                             //                                                    .write
		.mipi_reset_n_s1_readdata                                  (mm_interconnect_1_mipi_reset_n_s1_readdata),                          //                                                    .readdata
		.mipi_reset_n_s1_writedata                                 (mm_interconnect_1_mipi_reset_n_s1_writedata),                         //                                                    .writedata
		.mipi_reset_n_s1_chipselect                                (mm_interconnect_1_mipi_reset_n_s1_chipselect),                        //                                                    .chipselect
		.mpu_int_s1_address                                        (mm_interconnect_1_mpu_int_s1_address),                                //                                          mpu_int_s1.address
		.mpu_int_s1_write                                          (mm_interconnect_1_mpu_int_s1_write),                                  //                                                    .write
		.mpu_int_s1_readdata                                       (mm_interconnect_1_mpu_int_s1_readdata),                               //                                                    .readdata
		.mpu_int_s1_writedata                                      (mm_interconnect_1_mpu_int_s1_writedata),                              //                                                    .writedata
		.mpu_int_s1_chipselect                                     (mm_interconnect_1_mpu_int_s1_chipselect),                             //                                                    .chipselect
		.nios2_gen2_debug_mem_slave_address                        (mm_interconnect_1_nios2_gen2_debug_mem_slave_address),                //                          nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                          (mm_interconnect_1_nios2_gen2_debug_mem_slave_write),                  //                                                    .write
		.nios2_gen2_debug_mem_slave_read                           (mm_interconnect_1_nios2_gen2_debug_mem_slave_read),                   //                                                    .read
		.nios2_gen2_debug_mem_slave_readdata                       (mm_interconnect_1_nios2_gen2_debug_mem_slave_readdata),               //                                                    .readdata
		.nios2_gen2_debug_mem_slave_writedata                      (mm_interconnect_1_nios2_gen2_debug_mem_slave_writedata),              //                                                    .writedata
		.nios2_gen2_debug_mem_slave_byteenable                     (mm_interconnect_1_nios2_gen2_debug_mem_slave_byteenable),             //                                                    .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                    (mm_interconnect_1_nios2_gen2_debug_mem_slave_waitrequest),            //                                                    .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                    (mm_interconnect_1_nios2_gen2_debug_mem_slave_debugaccess),            //                                                    .debugaccess
		.onchip_memory2_s1_address                                 (mm_interconnect_1_onchip_memory2_s1_address),                         //                                   onchip_memory2_s1.address
		.onchip_memory2_s1_write                                   (mm_interconnect_1_onchip_memory2_s1_write),                           //                                                    .write
		.onchip_memory2_s1_readdata                                (mm_interconnect_1_onchip_memory2_s1_readdata),                        //                                                    .readdata
		.onchip_memory2_s1_writedata                               (mm_interconnect_1_onchip_memory2_s1_writedata),                       //                                                    .writedata
		.onchip_memory2_s1_byteenable                              (mm_interconnect_1_onchip_memory2_s1_byteenable),                      //                                                    .byteenable
		.onchip_memory2_s1_chipselect                              (mm_interconnect_1_onchip_memory2_s1_chipselect),                      //                                                    .chipselect
		.onchip_memory2_s1_clken                                   (mm_interconnect_1_onchip_memory2_s1_clken),                           //                                                    .clken
		.seg7_slave_address                                        (mm_interconnect_1_seg7_slave_address),                                //                                          seg7_slave.address
		.seg7_slave_write                                          (mm_interconnect_1_seg7_slave_write),                                  //                                                    .write
		.seg7_slave_read                                           (mm_interconnect_1_seg7_slave_read),                                   //                                                    .read
		.seg7_slave_readdata                                       (mm_interconnect_1_seg7_slave_readdata),                               //                                                    .readdata
		.seg7_slave_writedata                                      (mm_interconnect_1_seg7_slave_writedata),                              //                                                    .writedata
		.spi_spi_control_port_address                              (mm_interconnect_1_spi_spi_control_port_address),                      //                                spi_spi_control_port.address
		.spi_spi_control_port_write                                (mm_interconnect_1_spi_spi_control_port_write),                        //                                                    .write
		.spi_spi_control_port_read                                 (mm_interconnect_1_spi_spi_control_port_read),                         //                                                    .read
		.spi_spi_control_port_readdata                             (mm_interconnect_1_spi_spi_control_port_readdata),                     //                                                    .readdata
		.spi_spi_control_port_writedata                            (mm_interconnect_1_spi_spi_control_port_writedata),                    //                                                    .writedata
		.spi_spi_control_port_chipselect                           (mm_interconnect_1_spi_spi_control_port_chipselect),                   //                                                    .chipselect
		.spi_mpu_spi_control_port_address                          (mm_interconnect_1_spi_mpu_spi_control_port_address),                  //                            spi_mpu_spi_control_port.address
		.spi_mpu_spi_control_port_write                            (mm_interconnect_1_spi_mpu_spi_control_port_write),                    //                                                    .write
		.spi_mpu_spi_control_port_read                             (mm_interconnect_1_spi_mpu_spi_control_port_read),                     //                                                    .read
		.spi_mpu_spi_control_port_readdata                         (mm_interconnect_1_spi_mpu_spi_control_port_readdata),                 //                                                    .readdata
		.spi_mpu_spi_control_port_writedata                        (mm_interconnect_1_spi_mpu_spi_control_port_writedata),                //                                                    .writedata
		.spi_mpu_spi_control_port_chipselect                       (mm_interconnect_1_spi_mpu_spi_control_port_chipselect),               //                                                    .chipselect
		.sw_s1_address                                             (mm_interconnect_1_sw_s1_address),                                     //                                               sw_s1.address
		.sw_s1_write                                               (mm_interconnect_1_sw_s1_write),                                       //                                                    .write
		.sw_s1_readdata                                            (mm_interconnect_1_sw_s1_readdata),                                    //                                                    .readdata
		.sw_s1_writedata                                           (mm_interconnect_1_sw_s1_writedata),                                   //                                                    .writedata
		.sw_s1_chipselect                                          (mm_interconnect_1_sw_s1_chipselect),                                  //                                                    .chipselect
		.sysid_qsys_control_slave_address                          (mm_interconnect_1_sysid_qsys_control_slave_address),                  //                            sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                         (mm_interconnect_1_sysid_qsys_control_slave_readdata),                 //                                                    .readdata
		.timer_s1_address                                          (mm_interconnect_1_timer_s1_address),                                  //                                            timer_s1.address
		.timer_s1_write                                            (mm_interconnect_1_timer_s1_write),                                    //                                                    .write
		.timer_s1_readdata                                         (mm_interconnect_1_timer_s1_readdata),                                 //                                                    .readdata
		.timer_s1_writedata                                        (mm_interconnect_1_timer_s1_writedata),                                //                                                    .writedata
		.timer_s1_chipselect                                       (mm_interconnect_1_timer_s1_chipselect),                               //                                                    .chipselect
		.ts_i2c_avalon_slave_0_address                             (mm_interconnect_1_ts_i2c_avalon_slave_0_address),                     //                               ts_i2c_avalon_slave_0.address
		.ts_i2c_avalon_slave_0_write                               (mm_interconnect_1_ts_i2c_avalon_slave_0_write),                       //                                                    .write
		.ts_i2c_avalon_slave_0_readdata                            (mm_interconnect_1_ts_i2c_avalon_slave_0_readdata),                    //                                                    .readdata
		.ts_i2c_avalon_slave_0_writedata                           (mm_interconnect_1_ts_i2c_avalon_slave_0_writedata),                   //                                                    .writedata
		.ts_i2c_avalon_slave_0_waitrequest                         (~mm_interconnect_1_ts_i2c_avalon_slave_0_waitrequest),                //                                                    .waitrequest
		.ts_i2c_avalon_slave_0_chipselect                          (mm_interconnect_1_ts_i2c_avalon_slave_0_chipselect),                  //                                                    .chipselect
		.ts_interrupt_s1_address                                   (mm_interconnect_1_ts_interrupt_s1_address),                           //                                     ts_interrupt_s1.address
		.ts_interrupt_s1_write                                     (mm_interconnect_1_ts_interrupt_s1_write),                             //                                                    .write
		.ts_interrupt_s1_readdata                                  (mm_interconnect_1_ts_interrupt_s1_readdata),                          //                                                    .readdata
		.ts_interrupt_s1_writedata                                 (mm_interconnect_1_ts_interrupt_s1_writedata),                         //                                                    .writedata
		.ts_interrupt_s1_chipselect                                (mm_interconnect_1_ts_interrupt_s1_chipselect),                        //                                                    .chipselect
		.tv_decoder_alt_vip_cl_cvi_0_control_address               (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_address),       //                 tv_decoder_alt_vip_cl_cvi_0_control.address
		.tv_decoder_alt_vip_cl_cvi_0_control_write                 (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_write),         //                                                    .write
		.tv_decoder_alt_vip_cl_cvi_0_control_read                  (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_read),          //                                                    .read
		.tv_decoder_alt_vip_cl_cvi_0_control_readdata              (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_readdata),      //                                                    .readdata
		.tv_decoder_alt_vip_cl_cvi_0_control_writedata             (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_writedata),     //                                                    .writedata
		.tv_decoder_alt_vip_cl_cvi_0_control_byteenable            (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_byteenable),    //                                                    .byteenable
		.tv_decoder_alt_vip_cl_cvi_0_control_waitrequest           (mm_interconnect_1_tv_decoder_alt_vip_cl_cvi_0_control_waitrequest),   //                                                    .waitrequest
		.tv_decoder_alt_vip_cl_scl_0_control_address               (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_address),       //                 tv_decoder_alt_vip_cl_scl_0_control.address
		.tv_decoder_alt_vip_cl_scl_0_control_write                 (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_write),         //                                                    .write
		.tv_decoder_alt_vip_cl_scl_0_control_read                  (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_read),          //                                                    .read
		.tv_decoder_alt_vip_cl_scl_0_control_readdata              (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_readdata),      //                                                    .readdata
		.tv_decoder_alt_vip_cl_scl_0_control_writedata             (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_writedata),     //                                                    .writedata
		.tv_decoder_alt_vip_cl_scl_0_control_byteenable            (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_byteenable),    //                                                    .byteenable
		.tv_decoder_alt_vip_cl_scl_0_control_readdatavalid         (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_readdatavalid), //                                                    .readdatavalid
		.tv_decoder_alt_vip_cl_scl_0_control_waitrequest           (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_0_control_waitrequest),   //                                                    .waitrequest
		.tv_decoder_alt_vip_cl_scl_1_control_address               (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_address),       //                 tv_decoder_alt_vip_cl_scl_1_control.address
		.tv_decoder_alt_vip_cl_scl_1_control_write                 (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_write),         //                                                    .write
		.tv_decoder_alt_vip_cl_scl_1_control_read                  (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_read),          //                                                    .read
		.tv_decoder_alt_vip_cl_scl_1_control_readdata              (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_readdata),      //                                                    .readdata
		.tv_decoder_alt_vip_cl_scl_1_control_writedata             (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_writedata),     //                                                    .writedata
		.tv_decoder_alt_vip_cl_scl_1_control_byteenable            (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_byteenable),    //                                                    .byteenable
		.tv_decoder_alt_vip_cl_scl_1_control_readdatavalid         (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_readdatavalid), //                                                    .readdatavalid
		.tv_decoder_alt_vip_cl_scl_1_control_waitrequest           (mm_interconnect_1_tv_decoder_alt_vip_cl_scl_1_control_waitrequest),   //                                                    .waitrequest
		.tv_decoder_alt_vip_cl_swi_0_control_address               (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_address),       //                 tv_decoder_alt_vip_cl_swi_0_control.address
		.tv_decoder_alt_vip_cl_swi_0_control_write                 (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_write),         //                                                    .write
		.tv_decoder_alt_vip_cl_swi_0_control_read                  (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_read),          //                                                    .read
		.tv_decoder_alt_vip_cl_swi_0_control_readdata              (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_readdata),      //                                                    .readdata
		.tv_decoder_alt_vip_cl_swi_0_control_writedata             (mm_interconnect_1_tv_decoder_alt_vip_cl_swi_0_control_writedata),     //                                                    .writedata
		.tv_decoder_stream_capture_avalon_slave_address            (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_address),    //              tv_decoder_stream_capture_avalon_slave.address
		.tv_decoder_stream_capture_avalon_slave_write              (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_write),      //                                                    .write
		.tv_decoder_stream_capture_avalon_slave_read               (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_read),       //                                                    .read
		.tv_decoder_stream_capture_avalon_slave_readdata           (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_readdata),   //                                                    .readdata
		.tv_decoder_stream_capture_avalon_slave_writedata          (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_writedata),  //                                                    .writedata
		.tv_decoder_stream_capture_avalon_slave_chipselect         (mm_interconnect_1_tv_decoder_stream_capture_avalon_slave_chipselect)  //                                                    .chipselect
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                   //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                 //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                  //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                 //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                 //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                 //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                    //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                  //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                  //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                  //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                 //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                 //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                    //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                  //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                 //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                 //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                   //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                 //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                  //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                 //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                 //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                 //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                    //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                  //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                  //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                  //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                 //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                 //                                                              .rready
		.clk_50_clk_clk                                                      (clk_clk),                                        //                                                    clk_50_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),             // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                 //                       mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                                              (mm_interconnect_2_mm_bridge_0_s0_address),       //                                                mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                                (mm_interconnect_2_mm_bridge_0_s0_write),         //                                                              .write
		.mm_bridge_0_s0_read                                                 (mm_interconnect_2_mm_bridge_0_s0_read),          //                                                              .read
		.mm_bridge_0_s0_readdata                                             (mm_interconnect_2_mm_bridge_0_s0_readdata),      //                                                              .readdata
		.mm_bridge_0_s0_writedata                                            (mm_interconnect_2_mm_bridge_0_s0_writedata),     //                                                              .writedata
		.mm_bridge_0_s0_burstcount                                           (mm_interconnect_2_mm_bridge_0_s0_burstcount),    //                                                              .burstcount
		.mm_bridge_0_s0_byteenable                                           (mm_interconnect_2_mm_bridge_0_s0_byteenable),    //                                                              .byteenable
		.mm_bridge_0_s0_readdatavalid                                        (mm_interconnect_2_mm_bridge_0_s0_readdatavalid), //                                                              .readdatavalid
		.mm_bridge_0_s0_waitrequest                                          (mm_interconnect_2_mm_bridge_0_s0_waitrequest),   //                                                              .waitrequest
		.mm_bridge_0_s0_debugaccess                                          (mm_interconnect_2_mm_bridge_0_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.vga_stream_out_clk_clk                                                               (vga_stream_clk),                                        //                                                             vga_stream_out_clk.clk
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset                   (rst_controller_004_reset_out_reset),                    //                   hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.tv_decoder_clk_50_reset_reset_bridge_in_reset_reset                                  (rst_controller_001_reset_out_reset),                    //                                  tv_decoder_clk_50_reset_reset_bridge_in_reset.reset
		.tv_decoder_stream_capture_avalon_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // tv_decoder_stream_capture_avalon_master_translator_reset_reset_bridge_in_reset.reset
		.tv_decoder_stream_capture_avalon_master_address                                      (tv_decoder_stream_capture_avalon_master_address),       //                                        tv_decoder_stream_capture_avalon_master.address
		.tv_decoder_stream_capture_avalon_master_waitrequest                                  (tv_decoder_stream_capture_avalon_master_waitrequest),   //                                                                               .waitrequest
		.tv_decoder_stream_capture_avalon_master_chipselect                                   (~tv_decoder_stream_capture_avalon_master_chipselect),   //                                                                               .chipselect
		.tv_decoder_stream_capture_avalon_master_write                                        (tv_decoder_stream_capture_avalon_master_write),         //                                                                               .write
		.tv_decoder_stream_capture_avalon_master_writedata                                    (tv_decoder_stream_capture_avalon_master_writedata),     //                                                                               .writedata
		.hps_0_f2h_sdram0_data_address                                                        (mm_interconnect_3_hps_0_f2h_sdram0_data_address),       //                                                          hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                                          (mm_interconnect_3_hps_0_f2h_sdram0_data_write),         //                                                                               .write
		.hps_0_f2h_sdram0_data_read                                                           (mm_interconnect_3_hps_0_f2h_sdram0_data_read),          //                                                                               .read
		.hps_0_f2h_sdram0_data_readdata                                                       (mm_interconnect_3_hps_0_f2h_sdram0_data_readdata),      //                                                                               .readdata
		.hps_0_f2h_sdram0_data_writedata                                                      (mm_interconnect_3_hps_0_f2h_sdram0_data_writedata),     //                                                                               .writedata
		.hps_0_f2h_sdram0_data_burstcount                                                     (mm_interconnect_3_hps_0_f2h_sdram0_data_burstcount),    //                                                                               .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                                     (mm_interconnect_3_hps_0_f2h_sdram0_data_byteenable),    //                                                                               .byteenable
		.hps_0_f2h_sdram0_data_readdatavalid                                                  (mm_interconnect_3_hps_0_f2h_sdram0_data_readdatavalid), //                                                                               .readdatavalid
		.hps_0_f2h_sdram0_data_waitrequest                                                    (mm_interconnect_3_hps_0_f2h_sdram0_data_waitrequest)    //                                                                               .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk            (),                          //        clk.clk
		.reset          (),                          //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),  //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),  //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),  //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),  //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),  //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),  //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),  //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),  //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),  //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),  //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq), // receiver10.irq
		.sender_irq     (hps_0_f2h_irq0_irq)         //     sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_irq_mapper_002 irq_mapper_002 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (vga_stream_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (nios2_gen2_debug_reset_request_reset),   // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (vga_stream_clk),                     //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
