��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�x}��j��S�b_�)F�1�(d'Â,L.��ꙺ��e�˭'�{���)�Ilf\�@,�y��Z�n�X�D�P��c�����=���]Od�w��yD.΃��o�N�o?ղ�*nek��XԾ��(�H4��ov
�_�U�t�
��΄kdaq�%1�
K=�?E���P14P)L��Cro��$g�׎k�����-��o�����N�=�s�c��Y�ų�wK��F��M	���'6�`!�k(�:�niGo3���y/zfd��C������8h"�߭�&0�X�(w@%Y��~!ʍ؇�������}�����|�"��HS��]�i����#�yH v��$�W6j��9L�'q�h�U�淰�W>�gn��%��\�j��1���ɭs'[ l}_��ʳ�/Xr��@7���?�|Y�Q��*3UE&0v輤�cY��w�q��}�'�
�Rf����0����W�q�<�=5�S�����2��ZV�N��8sO�"�G/F�T�WĆ���yW��D�L=3h��g�q�U9�9��)QSCW�Qf�Q��K��S~Jӥs_����f�� ��6@�Q��"��,L�	�	˸ʆ1G�Af�N#�e���r�'�,�pc��$ټ�6�|���yą�D�ie\�mo�AH�x���4%!�LK�7�A#��(-��G�l��ۂV��G���+v��ʜS�ڑ5]�U]�\�`�m� �A�>V�5���m�|��,��υ#����;��z��!=��嬻��U�UOH�iJ���tcð�))��X��ɭ<�����(�fT��Nx3\���o]O�Lo�C�JzW)���G\@qKo�����Z�D�/�����T[��u=f_���7�X�tԠϨ�]��O4��r��징^���΂U���<C��c��_=&�P���Wȋ���X�Ć,�"�u�龞G���$�U@/	
�W����C�..d�D��V���Ɇ�tY��L�=ň�(8I#4C��,�.�E�0���i��+=~� �~��f%�s�(�E�$�q��Z����B-6P�|�~-��=$���pp�G��?��H��v��oW�d���F[��_az����i8�z�F~��8Ѷ:A�W�M~���}�F9X�w�R�j��|T�;�C>;>�/����;Dm��׵ԪTkҘ6ᝳ���RQO@���mj�W=�=�ֹyd�� �	����tXcUA�۩��d�"eT�ܧ�:�@���S��6ʀ-�Ō[y������Ac��w�n�4`x�7���Cs)���j��@v:�	oK����(�f�+��JqըrRǋ5̓��
$��5|�m*4�HTڮ�݌���eٟ~I�����WĶ�į�����f���M���O�w>Ԇ3�+W,�N����9��[ z���ib���#,I<��R�|�7�do��)�q�UVI�B�ݰvJ���;���,g�k�u�[=�CP{��n_i�L]�Eߒ]�*{���N��o�`��N�&_��?�Hg��� ��^o@��2�^��4#�_�
�#�����9Вђ@�b��Zq�	����P�}@Z�`���n�c�s����m���}�#���Q�t����l4�4e2���l�,�>��@��\�lʹhW��f�V����lw���2V>?K��2�g�"���rI�@�3$��o�9�� �}ˉ�+dJl[��w'I��+�R�d�Q�G�k
�<�YѺ�/5�(Y]I���,: $D��W�O��ử��K��*�?�x䲼��b��?(G�����s���=e�n΋�����)AX��*E�H}�i*R�h��>��aj�&����T�_��u�5�v��_�" ؋3'�^��HLr	I��Cr��aыXq����TTԤ�V�jǸn�tE/��ps�N6��9�vo9��r��K�,��.�
���;i�L�Q�[�V�9gi`��Ɨ؍ ���xs@��Kur֍�ioY*�*�N�O{��C�ʟ]�^���>��Y6 Y��GK|H�����:@�B�2�I9h���I������>s=6��ٸ&3I�j: r�O֙"U�灢���\�(��+N� �r�����ׅ�#3�}\X�*EQ�r�_�d~6�o$&�i�m��k�l�����M\ 1��MV^���-��ы� [kVG�󅘈�yݓ�-,!X���&��%���Ϣ�yB/��`49��[.S�r#��W�P��)�N5���(��k�e�i� �ڼ�V&��:�>����n�8����{l���3&��@��ڛj��+���m�;6�h���{T��g��frq���C�i��e����;��^l�طMB�^�!������p�R�{���U���o���W ��˷��#�p����^	��/,h�˽7�p�� H�I6tr��a��ަ�M%!c[ȷ��-��Թ�<�@~�E�3���y�73�"�Ͽp`�=Fr�JW���W�h!f�o=OU7B��b[Q�����>F7�كv�-�����ԨE
�P���y��6A~�S=�vܟ��G�w�R4�g��Gވ�5�1P_�f"̊|��N����5 6Ȯ�%x�Kl#,����A?(��6w�e.K���Di��U�5��wP/���T�/�����O�t�3�D��Hȏ���F'į{�%h��LU���[/�%/�S�|`�~��4qD�N!�%�W������,�+f�_�g�)��p�Z���f���Wa�-&k���[ɛ��jǷ! P�_��5��1L.��[J�p��\!p:�j��-��]� ��V�|I�~�]�ҝ�P��s����ڈ�p��b��>1�gS�@	��i+��t��؟U�ggN��.������
�Vy,A=\�����I��Y���=ű
�����	+б��.�G�PCI����j���Zv%���J(�ÿ�慤PL{�5K���f�%w�c�$�~]H;"sm��B;�i��.������6"r+-�	����.�x(���8��ބtF��F"��?к�)�����~e�Y�"E�k@�o̮��K�j9���4k�s0�T`�PA���M��ş)]�'����Lf%�ڎ��$4�H�c�?��+	�!|�2�p�1��$�#�a���s���V�f]%E���П�9�=������'��s$Y]�"�N��_ �E�-F��˫�����e���6T�n���\��"����`kN�ZA�*����c|F17yW*Sj���������Ti��N���7I��T
i���@_�>۪�v��&�5����2WU�Q�g���΀��F�-�r�yPe��Qׂ�T����1ܤ4NO�2��n�-â=�s��\kXO��b��7 c��<��f�(U���w@s|�!��%�T\fH\�e�=�s���2Tk7�HT=e�/�&�L��.��W����kwCA����vbrd��_s!��5k�c3�*e�Ҫ�A����x��i���)q����^U?�VT>��ө�#��,�$�� o�֟~��2р�S�����~��5��ۀ4J���}���z:��قs��S!�{�1nQӋ,����,��Э���SC��~�7�2 6�	[RQ��U"���ym��xc��t֬��Ө$#��m+���^�#3��A	��-SlK�\��������{bȷ<(��I��n+�f���>�=B���H����huq�x/:v~xR��%n���L}�dпl�M��r��K<؏�!H�Zǈ�����ƭ�n��nzv�Hk׸�'�a90�(H���(�<�ә�%m��/� BG�H�zR2VbM_��Ȏ�6��ߪ��!�>�A�����H�C�c�Shb�5�7`��)պ0�@�Cd���Ǒf XG��j�V'����$�hnQ�>��őzD+�J6PV3�墍��	�#ȧ�.��C���oH���uq�Fj�US�
G�v^w����6�"|��b �
�P��7m��WS�/����+L_1 �*��(+�����D�
�ʅqQ���Y�朮�D�H\oW�����'ᏡYŧ&�`�9Q�-c9n��*����>����!߆.���(�d��H)� #e�c&x�b�x$��<6�$�e�\^���E}�(�O��Ѱ��;��]�R�
#c~X�G^�{d�<#���}��C-��D.[�sB
^��0u�Q��6ݩ�SA��
����f�c�h��j�e����'��*K�Z�I�:���p�FV�5.i=X��K1���ҟ^��"�@�f�9/�o�b�!�A!F1$�]�pĊH��-���hK�!�+��Ô��4̐��	OmB�W�l�gok��j^�B�5x,H߾o����`���֊���Rʀb۪�lP�rҶ;X�ۅ��Ú@ͻ�G�!�Ĩ�2�T%b�x��v����a��O=ﺵ ��X�~tXS��V�C��!���楜v�����Ų�9ӘC���M������p�q���--�J���Q5�����d�㠫�6Ђo�89��A���ǈ�8ِ��A2X��tQ2�&�(1�,�bt���L@6�,צ��Ѫ�VЧ�wt>���S� ����-�e�y>�eDr���j�G��۳ �^��"�w�-�d��#;�-��W'd��.��^SY�/Q�uWW��|��p):і�?� }�0=�lq���D��{�&Sw��ĥ���v�����!���_��P��ı��ػx�Y%6����c>�D"K&*��T��[�aW�*�� ���=ӯ49�`90Y�:"�t����tLv��n݊���)�Jb։(�Idy��V���g<�T��������6�cPz�>��WC3_	n�"�1[<)9V٧(B�+��-�8O�#��οF�8�=�'��ϣ��g��c`B��r;?g��i��
�~��h5K ���c���짼�LuK��Q��#JV������(�f*�H�I�?���t��ҋ19)KCb���h[k��G o|A�����է 4V#�5IQ|%ک0\A뗟'6��&J'�R׃'�mQ�4DŃO�ߞC�� �O+KrB�F�`�\S�e	׶�Zt�r7�G�#6�ꭟ��	��u�5��΍��t�/���W������"�u�iII[����9?�������UN׺C��\��n[ϓ,�ST����'܂�Ά�;�L�R죻Ο}����\�G�ۗ��=pg�8p�׭�A(m=�,�w���M?3Z����y���V�mk�=�	S���}@��o/�(E�[x6��L�c��-v�b�>#<�����w��V�+��E���=�(������s<�M`%��q@�Ktc�V��ѺA��Bo:M(r�*f�6��D�Q5"�(%_�ŕut�U�~R�mE��Ȋ��hy��"�U�ֻ�h	N)t,��$��W�U�&c�z�.��vNRf������n�˓a���Y�{3��z�[�̣�,�dqއ��3�݌�A��d�\�8���#�a�Lf^����s�9	A1dMMkl�z�w��jN�'H���^;�y�v���$�ڶԄ��@<ֵY��cb&�4���������LEI���;X!<wEj���^'ɸ��t�wR�����r&ѿ0bR�R6�ƻ<�^��k$�r�C�G����	���G%����>=
�Ǒ���Wo��C���G#���+@���������|���Zg�5[5;�������h��P�)*�����dKl!ˤ��T8{����)gzE�fx:��i�s�ĺ��v#��i�V�:�չ�A��6Lg~L����w��ɰ{edۗN�}4�wIc��3\�pZ$��?xq�6��n$�#�	��"\=�R�INˁ[y��"v��KY�	2%K3��J�f)o����%��3�<�Z�Z��� e�@�XQ��_�Ӆ�\t���-~�����i�Q�� q�s���u&�VN��}i"�D�X��ʁ���nK���J�\�&�O��gU�t�^r�8Jxjr���3�8�����-[�DS�f����):�����x�.�s��B��s�����D2*a'�}sm��-x���<N��t%�D:FcE|��t���bf�n�k�r�O���J�5J�6Fy;a�bn�*+���ɒ]P=6Hխ�'�C$�@�W�3��sm���HX�Va�(� �,��E��.��|s�;��Nk^@cC���bw�C��7�B��*��3g0-Hz�*$��`�-yLpz)ęl�WR�Fe��R���ΗoL���R���A�~�Z}������@k��ۥ�7�(H� ����M�şi]��%�|9&P�Y��?:��+�2��|����i���.����v�Vu\���~
{��)���o?`������I�H��D�v*������I���e��Q:�y�xraW�F�B���Z�Io���Bg�	 ��o���aT4��x$O?���鏈�`i�b�f(%{��|~�-�h#�-A�L��B���W�M�|��Timj���!����p�4�Ȍ%jfsy�%���d 2�*�]��9C��E4Q�++�e���j��9��є�:<J؝�R���Բ�G���ᠹ踅=W������W8E�����Wnˠ�>D�5�����;����A��I�����v�х9������\�Wّ�͜+m�����d\�+�p,ZG�e�D�I�Dj�"����w|�TM+;S���tR�D�N�#�������ô�@�9��K��9n��\�<?�Ub1����I��l��M��4Sؠ�x��9���kҞ�Q�p�񄿏�S��a��֍���L_?.L��X�r�NDN�ԫ�z�@-�)��SS��������ܮN��:`O��,��M��X�a��O����P�K���^��ʕ���uy�+���K�a�2�cbΟt��]����7����W��>�'؃���K|��wgῖ!j�r�Õ���E:m~��7Y�
E�Wޫ�� ��ߴX�WSY��`�����/j6j���蘽]�)`�C%�����t��%�]<`����]{�g'M�e�%��5u�!�I�ú�P��ق�*�*�]cnd}T �Zi��,�~�|;���4�?a��"Ěw�1'f��ȫm�B<��t��t�0%�j��i#��&�_F+�4NH���g!;_y��5M�N��l��z5��(�ϩ�	�<e������ ғ�l"��E`/��Ȅ��h�Z>������⡴�H:� F���@}�0�BFox?�h��eM:�M�mԸ�ꥻ~�A�؞p2l����?Wy��a�]�ݓ&�`J��ZMK��Q�f�)r��0ҿ.Z\�/Z8>�8��i\����,.��> ���na}��=-�0��=9��G�_LM�j�V��5)#t�ǽ�*�yrbY�i(fi�;`�A���y�Cū�ED�lYT�A�!<g �y�L����,���R��l�V�D4��u��%B��x�u�-ܰ��,)}�J���٦{xPk�-�(%����e_���������:�H�$���B�x����r��>��Laʑ�;��aٖ�0�c̩����̺Q�M�ɣ	�&'�P�-;��4?g��.戨���7Ҏ�)-Sy+��F��
u�{~E� t�wZa��T}X�9��C�?uDp�%=����A�j�id��Xj7�faK�`�8b#(S���G��H�*qy?{5"�uT;+Ⱥ��!��|l]�C�H�z>T?e5t�Z/�)S�����	+����z��\�w^K�,�Iq�!^�k�:���H��b�Z`/(���;��Z��'��L�s��Z�B@Mx�q��$��*"�x�V�H�U��@�'�3�w�O�u}�K����)��)��ڗ�� p����"LD�
�}���D�c�꒸� ����}:�j%e�l����k�|f����q���(�C�}l��	tSZ����La~����/nV{������q#��٢		�g�?���?
y:C��U�8�Ò8"&;�D��δScsj}-�|� �&��i�Ӎ�*�R��"�N��R� �'X6�X�����,{�I��1�6�|C{h�8�kz�,�\�BZ�pKN���g��[��݆�Z2������$��9�	��s��K�Y�ZC�qm&S��_�d�V9p��~R��[��k2n��P��N�	EN���?����&
JԢO��q:1�S'�(ag�1[cI=+T�d���U�=t��F������$�6�ͤ|a���{��Û"�$UmLZ\��`~��$5xY:��4�h�P��^��X����'��}X�2�<��i�<Z�-9�y`^IU���͘���s����F�:�Y�&t��x����r:_�B�������/w�w�vg����'�Zܛ9�tFW�[��op��32�l��ڷ6㕚P*We��"�S�_��M�פ��1>]���T�Kmg�v��]N��)	�{�񠁲r6���g񶏤%���a���/��+&@O����+T��!^�j��Q�Ps����S��y�����������JSH(^ wzLE9��h�Q~����+o�����GI`�!���@�^1�z9b�fUscp~�W�u�(�B��VĎ�X;���n�B+�����@�H-}�y����Bb<�Z�����ڄt7�
&���s���f��60�Vƿ��<A
�<�&Z��G_~֠��,�ɸ�gc�t���J���=���$�G��J�&�߾R!J���w�-W]�
FL`�]��a�c�D�Ȗ�WN}��4|�$k*bƶk�-���a��n�:aYqɩ�c���O���ߙ��x�	��ӕ�u��2l	z�ӮYĂXG�x��qXsL���͖�'��Q�#FA#���8ym#�vh,"���,�4�K������ƈ%�}�w�������pmr%K���w�I0y����ɻ7mIan�+�W����n^O�x���`���u�Q@��.�Gd�8�o.DCgǭ��>]02C�'o~���P ,�q#Z�*�� a���)~h�#�\сO��-2D�$��T,���iDY����ϗB�8�"�s](���ˢ󇮩l�2'�w1X-��:fݾ�G��j��r�{��99�6������I�PS�C���ܞ�0�:9��%w��Cʚ���D�c|��T����՚Y�wjI�2��N[
N��U���Mj�G��<��=�tsSj��Dg�1#�����j�^�򰆴�����t�L���\ z�wHy�iʯ��3�U< 9E��eoQ�� 'Sp|K�jU�w�r�Brzz�ޚ�YU���[3KGw)�*�J�6.Q@�Ǽ �EW]�v�����%��m�!C8�49��x�sߒ�{mXAz�~�~��鞉��es-�ܱ��?��,Y�W!�K覹�uh^��Bě�D���J�A�Mɾ*�M`���̧�Ԑ���϶&VO���+J�?���L:�Өw`2�<��L6�����o��&�e�`2Iyp����Acr�^:��4���j+3"�ڪ	�x�\v �����vEd�g=`�T�Mn(}�cXN�����]@��$X�F�mv�I��U�8X!� �t�8�x��e6v5a��H��;բ^�C��`TR.9Q���WipϤ�b젲dg�&5�9��3�0��ޚ��=��a4���Sj����Z�{�Ϡc�Ä#E��&.0|� %����L��7�
l\m��T�SrےиR!��?iB[c��4��Li�B��O�Dp���B���d�2�E�`%d�}H�>Wm�˫�"����ɸe㯿�Z '�i R��hT����
��Mf����q�8§�;��֟Z ���"�j��R�K�x1������t������L�Yt���-�B#yE��/�UDW�o��,��!��{y7�xbo�Ftt�!��|�7�H��a�=�Y�9�	[��>�8ѡ�b8<���W��.?�
ߟ��'��O���_�o��j|��!��N'���j�Xɣ�m��'��|zIHgUt����c�-�$������bo�y��8��
~Ý���kb �z]��_G�����d��K�����@�!"��)8�����̬J�	���*�g�����>B���>�HL�� �]�`0F��� ���P�=�s
J�e� ����3�F�H���s1�^L�u2���؇��2��p^@��Օ���P�I�ԣ���E�68�5��)@]��J�	�խL�Z�2m�c/�[��CIU������4�C�;>(�Ly�Ծ�/0��2I�H*���d)C�!ϑ�O����n�07�����{�=`R�T��Mb�0 CYÇG�LWCE�̳ݙalk��a�q_x��ح������b+�
���K� P���)&�8^�:����%|\� �����a���f�=H�:���A0�ɤ>�C�� f���L!]D�j/��dĘ�mQ{_�R˾��b����]܎�Э�@�J%�^��M.J�Ϝ����P�u/&7d�UQb�M�g�f��F%hC*�%O0p��Ψ?
�瓈��/�C�n>c%jkc��:eϖ�$�Ə����D�"=A#�ќե֟���w�y���M4�L� �M�/����M���F������?��ߔ�E�M��[Qa�H�*d��R�M�!�b�^�$Y\+R���t� �'{Ozd�L历��@!��yW'��(����Յ�\� ��;z�Sq�
k��Z]+&����@�	&\��A5����z�2�1�3/��_��wpv�2x�9j��V�M�j�p�8��:�W���p�ٓy��e���
f�)F30H���-g��
�����|>�O�s�@@�W�i[EK����Iye��������Sy�ٻN���W~h�BIL�����~i��Ҽz�~*ۘ�Lf��� �-�jC�-��ɚR����jj�
�E��oo|���U#��)n���E.1ӂ-��W������E���O�os��̅�8�uW�a���uX{=����uf^úWa3;k!�ߙ��M���J�i8�c�h��*��ԝԫ��_��j�N
�9Ր�q�"fI��ω��G�zu|�s���#�n����p���H���wW=* ���n��I�rK&l�M�v� ��'r�7x��ja���a\�Va���o+���KI�`�/��y���3Q��U�U������u%3Ҫ]W�a^γX�~O�Z�u8�E_�og��˗ѷ�u����Y%��Mݵ>�ɸ7+�arP,��P�-����2�Qנ��sT�+y�I���R��C��wh�2����T�.D)$}BT���#�y��&���,HB	Я�ls1)ة��T�m��A�aU��Ea[<��d�%��L'���
�7?nsE}��=*�c��O��憹���>��u��*����_�E>��[���.�7�ӵ��i�f{�	�L���Aa&�����~�UGS�Ґ/�yO1�M�����IElm��l��2f�C�L0&���b��WEm�xɈ�� {A���2��SB=e	�ʧ>�q���'O��w�qkC�P9`�`&H��o�0�ڮɺ���(0�LS<C<�0����J� M$T�<5��1hNY�[b�T׊v?X3H�.���MN��l5�K�V"@��S;i��7hj���~�(���<���{�jFNk��)e� �ѱ�G�e�jZ+�s^�o��q�^5�p�ؗ""��L�%��pv��[0Z�w��Y�'��X����䅸��^��]c�vÓdhn�-AF�n)��'󞩘pFiE1�d���:�&�b�{��.9���yJ�m�>��<��k�M��N#���n0�t*ew5\z�A�R�zw��|� �v�B���g�J�\�ܫ	���9��G�W6�Gt9g��#Œ��5�H]�)�p�׭�I����w�',�^�V��`�>�A)n8�3���=s�b��U�B
�N4�����Ո������������k���\I3���-�;��'�m�
��׍��M���Y��T�����b��*8G����0y��~�a��7s�Z&R�t��� =!�c���G�m��#������(h�{Ѧ�k#.�'�4%�y��R�S��}y�Io��a��x� t��[�kX�N00]�	�i͇:롗xq�_�$�|E���SgY�@��4��7���P*��q¡c6��{Ҟ`S���������8V[��s�t�Ah��7P��>��-�*Hڣ7���x����� [�y��nm�1r�X�g>�iJ�у�i�$�����h},�F!��R��JC�鳀AY'��IT�\1�C�x��u�x�ve�&�n�6��-s�Y�Q�O��Ac�Y�څᵾg!�Հ�Ai6��Enm�����"��C/���sĉ����䊄#��<%e{g>[3�}�b�����0��z�,�����U�)'O���H��x�A-`f��VE�p��2D}a3���#�;G4Sm>x:��=Qp:ݒz��t+���	y��N(��>�C�"��`��h}����,NX٤���N��e��4*jyG,jǇTܥ�^]��8�Q;��э�w��.Σ�u�C)��Z[��wJkn�]�{h�4T�xCؐ�����!�$�Sk>u�US�2诲��"S7�v�Q��'�0��ӣ�aGHDoTm��F��p|J�>~��j��|T`'�o���x= Y�Y������:�f����b�[���`����9�I��^��Ln{���kDYC������ǂst���Y�ڦW�  ޏP�5�B̖��������O%|��ydi{�Q�F��I�V��6���'����d�-F���M�5ٸ>eNM��j�D�9(��>�#��ZGضI~�.�	�	��w�(��;��U�)1ϳ
S���K@�OJ	���w�ۭ�bj:o�����$pZ�J�r/g"e��N	��Ә����js����`�q�5��q��?Oˢ8ky�!,��a�3���3'�K�
��&���!���1�.5�J$m;�b߂26!J��}�Ծ�י΃��7��_f2"��|0�V�^>v�����mr4BYKw�*-@ab)��Εe�U�B����F9(5���ս*��9���0�ȡ���d������X��xжPB�t������rw���"�\rf�/Ie�a�&��@i��������zK��{���|�c�|!T�Z`��t���#W���!��{��YN����6����d1-��������Sim�-lz�`:N蜙�r��O�9��b�S&�<Z���a{���5�|$a;��#pl7�	�1�U�Cܐ`��4�
)������:��T�ΪB�$�2UL]���w����,t�;�r����f�@KMR�'*+N���"$`�^��^%s���0�&pP��掯` �� K�6�\�X@��7��&�*�Q�0��� �U��29����~��Mŗ�F�'����]�)��	O����Ǭ��Z�^�n���"�i�+���Y��	L��Oh�bk�2�	F�KH��(�OS�h�,�h�����u�ϕ�&ZxM���ب3Z��p��șԬ�j_�;�u���ǹ����������@DQ�*���5%�"���'
� vcZN:����ടM��-�刟1T�Md���?� ^�f_1�`PLP�T�y8B�W�(�Ofd�Zw��̍fVC��+2ݼ�Z�,��=�t΀x���'�������rc�������F�,���Z�xM����7"�S���KWJ5��&��%:�F_��s �B���]��߸`Jb`n���i��1}�g-�\�BHSF{]�60��JLg)��������Jj�*]�^�FM���8u]�v&=�n�h��/�,~blF���L���nI�ɬ���n<$-5�����Y�TS�|��_Mvr�8�&�Ec4]
�/�����G�@�=�K)�f$��A��IL�.�����`��� �0�l���D=7a�cQz���9������މd:!�ӣR�Sޞ�W�� 0�8�'o�"YO�w�����U��t�Elf��s�xߒ��f���R�ɳ1�3��n:��F�s�����p����`o()�������z��
8��3d7�.��0�����C���yQ�b�d-9V���`dh��r�rE�|gH��!�̟��Y����f�~c|�m��a��G��;��4���1,E<D��P�y	��d�b, ��!ՙBy���ʶ�V��g?V��Sۀ�T�e����i��5�,*�4�-������N�ܦ�ڠꀦ8�a���Ȗ�܊��-q��5N1wG^�b]�|<�YO�0ؿGc����Q�܌��:P~"�I�#�}�t�X\��X��Bf��������2\���}��*��||�������W��$�.���s9�v�J��b �IU�]�OE!�؃��U^����H9�Ƴ��ݯ�D�v~���T�p���ż&��t��O��ڽJ������z���II���f.��T	�� �z�]^�ߌ�pR�yJ�_O�� � ��6R~G[�Λ�0HR'\亾�bx�1�ě�pgEؘx[ZV/�~��٠� ���OVЎ+���/#ghY_}����Q�~V��Zu�����;&���u\�0���m�@�'�ieQq�d^ a�i �����C����5Ø�Iq~i���i^��m�,��.��K�L�޺�gk���w��{�a�,��װ��x���2j��Xb�q)]{̃���w�5��A��7�U�)��?��oI<���f��92��8|�i��t~�ɴ� "aeI���a�|(nDRI��|�N�E=8���
h��H�"��v[d�_�4o��H��$Sl��n�G��%j����8j���w�L�9�>y�<�Y�YH FJL/�����	�@AGˊ�}��r��C���a� ��
v8�F~�2N�f�f���r����i�v���h����N��+��w�c��(��� ��WQTٜ�u������OzgL��;$������_O�g� !U�T�F~�bڑ1��4�����;n��Rb�膧��?pH�H�,"k=���;��T���]P�ؠ��^����ĳ;S@v���݁�j�V���_č�a���ү�t�\M#2�䯭��d�J��E�b+q+p��䴁����W��AۂKs�xr4 �B��`z,����y��-%��V��.���:Y�#����RC�U����S�������xI��]/I��)sY$���T;o0�k���W��Μ~������mX� ����o����I:�녇��(�n� ��U������oYsgȝ�!�	�kZ�r���y4��'-�fצ��#X����*����
����\�F�+�x�@\�ƅ��ȋL���С���ž��_x��h�+>��t=BA�蚦_���;�吿Cd��۶d�G+~%�x�9�o���EGeӹ7�fy�tp�ah �q̋x�F�6�2k~ޫRx� ����r�>4Q(��$�i�e�[�F�D3�PO������J(yj_��I��YQ�+����|��u@����K�_|�ם$0�^Hy���!��r�ǰ��1�c��E����,�wS��3�u{M����d���]�	oQ�!i�v����u��b]yM:܋qQ�v�Y��zyn�qPv5>}���0#,���]@Sl��H{T��\�`�$�Q����>0���-�9��ݑ�t��G���LǸA���e�L���颲�}�G��Τ
E!3u��d\ g
��,@�D:�
��?��U�Ή��:! ?��Q������v|u1q:����L�gl�n���Ax#������SCf�p�,=��
�2���J�	Q�բ.����f��4ل������iZ��^W<���N'S@��)���4���������HJ��!eؙD3@�W8�` �d��/ o^k����/\�
v'���0�% �� ��O�z���Ɇ���\e�Ak�����O��d�(6����_�ܮ�\&����M3�bl��sdXT�
:|���%c��CJ=	���r���G�E�y
�+�se�+��ro����}!�
�
F��N+�shr�H�"���j4�:�|0���C.�s�1�Ǚ�
t�c��g��;$���0���Be)�D�z�r��s�����anJ@�cer��,]f����5K%�bQi�O�P�7��4���Z }�
�;�-oS�C�Y[�#�k�?z
WaЕtr}��ON����N�3(*�;�D�f�D9�״_8ZR��W���MR��}�|	��CD�8ԣcR��E�T���#����O*�ܙ��eZ����rF@�g�L��7�P��񰔋2���+����᰸h��/@z��.-��d�f����C�B���Rl.���ba������^��)Ȃ�h:�ml<�2���is��������e8�0�[�,Y���ǥ�r��_
��p���� V1�0�}l\��`�3^��o���n�x!�$��c;ѭH���>U7�l�]��
 &=��H�]��8G��S�Y����	�ǚ�k8����CΩ���L������b��x!,���\!vCkM
���l��E7Z�oU�|fw�.�xcP��I�kk�a�.`�,�W">�)�:��ՔG�t�E>�Y9�z1ׇN`HM�62I�:������U)�yH
�u�S�\��z�54[��e(kJT�������ڂ�VZ�s�z_Y���O� o�Օ�W�M���]+�P�M���")[����v˙B��vN�Hao�m��̩�`K��*�W�'�e����hI�k(�ehqL�*����)�t��N��Pme%�{��F&��眙~	9����a�D�;��AnO_l^�H�.i5�
D�k�:�]XҮ�p%�}b|>`y��fLH������bc���Y1��U��W��B��3���3 2�͕�0��c~ƣҕf�,�Ik�KDn�Y��>����'�mv��v��3C�����ӵn�*N����Q ��$h	RBK���g��T^]0sO��Z���m��,��on��s��!��]��Ê�w�C_	�����x����݋q�I�h�Zcc���s'�?a
S���t���$�����Ϥ-jN�=/*E�.�mÓ�v�P|�*�b��5��/�H�����d�_0m��<�����j����9!ߕ���B;�H2�-/�Bꫯ�V>��}*��!=�A����e}l�z.�h�2	?��Z~Nlzy��Qr�VMs�SD�!�g�X�2��"rl�ߧN�$�� ���B���57(�ˈ~$�˹ݍ�i���Y5K�Śc��I��:�t��3To�y�b���G�Sծ��\�o�Y�9t{=��?ߝ�2ճ�U-��4����h�C��>�>�ks�� [��a{	��ڵ�=N��P\-5 O���W�Ŵ�@�ӡ��	�&+����ej�F�.a�����!�կ�׆:'�/���ĠIdu+P��+2`cV|�r�D�)�DЀ;��8M%�&0��ф�`N��~h��N����T�+�-�N��iΒD.0g̻ۘm�<}�I;�9�����G/y+���V0�ldy�:K��4�ł��;�b(jCbMi
�=�=B?�-��=·��ɲ��� 7o�ğ�l�f
QHƲ�K���4�	۲@�MI>����Q�0A�'��.�,�nʵ���Qy�y���`)����	��Pr�����:Mߪ��'�����j�%\��3$7��P��C�ߥM�|S��ʇk�"�S��"lrD��<f�
Y��,�ZC�� G�+!�����O��;�C'z��j���;�h�OdZ����VQX�5�m�:�hDk��3λ�z1����|�+��]>�
�V)�L�}r��$g5uRp��!v赌���Q��T_�P����H��ɞ�^ãA�"�#��Q_�̌�'�te���7�-$���m�Ozxe�/\�e&�M�q1�8��爂��J~��P��}$'�n�2�5>L���?̿�H�x�UeՄ�g�x�Ub�w�O��[M��w���HaX�J��/x�_�L��ȼ_g�;����-?w���\�Ė���=ݿR�y
RHG���ѵ��fF���bs�-���k��2mnM �M�*��7�߉��򱥡��"Д�X��^��Hd�Yf�ccɶln���M�FlZ5���{a&�x18J�[y�J8a-�����m��9�ɕ">���v���5��Mo���п`B����>�:�kI>��]C��sΛ��z �ߏ�a�VS���NN�6д�ȣ-Tk�$^̚V��hXj�x�C�����`!��Ś�,e�i���CC�/j��"E[���e�*�,H��OTD���:E\�-)�Q�e��ah&X"C��yNk��U��E�~�:�tO>j�)��P:�CE�"�_S*z�~����iK�O2;C��_Z|m�๨dW��,I�h����i�o3et���2���o���}Na<j.ݸf�m/0LX��'���4�4�a� q�3~��::����~/H<�=�k�oȲ��j�ۖ�������8�c���CUb�N�Pц�_8c]n�u,쪸�u=��l���D0��8ny9���o�>�"�������4ʭ�TҠ�s[{W�_Z=�:�z���N7��߹��3m �5ׂ�ܭF��JAA���|�bn�*�bY��Z��o��{��0$)>5�bUhl��W��/��0��	!RL�ɿs['�h7�2pP]V�����c�Ъm�x�-6I����8�����Q�����������Đ�)�̎Pr� Yĉi-k���Q5�s �-���9�TB��r��Q�/����� 8;� �]���z{��_��1�o-I�*�U����m�mu�<k(��0��x:����)S�I=��A�������:'2�ٰ�b�Eӈ�WRh�JVI�(-PC"����&�F2��һ�*�8Rp�Y�:��>K���D�3�P���}(�sf>�4@�M��^�Yoz�� �ct�gi��k�wz��ajD�Q�����%%&<��޹`�,1w��7����29 GI����
�!sC�$�:E�a���y�#��e��1�R�]o^����69wM;�B��t�����@ǎ��>V��l~�VN���*����⹭(��ӧ���@E��GUjw��V�V�3=z���'��Z�4_�u+�S�<�-u;�J,0Fu�#��^- ��=��Ǯ��ǔ�sg�`u��^斥�u�y��������Ч���>�&�Î�sJ������"P��*V'p��q�by�w��������SPc���:�6��\U�.}(����c�lvs����%�@wi��췞�^���l��Y^�_&��W~L�e&������핒�J�Ta|��YB�ia�J�h����g ��:�v*�fO�1��U%���&������&�x�(-��w*�B��)�Zr�
"�]ŭ^��lxϹ�|��Jm����)�.ݜ�J�h�r�x]�%M�f�!e����6���D��)�x�вC�@�q�Iq��|��_S��<�#��$W��Y%�}�9�_��0�֡�E�z�=���ܡ)"3!t���Uh�#�(�˵�,̑��6{����b<@�1�����rY�\G$2 �d��#�$�3��m7��UbH���-3&DT7llN��4�ȘB4]�'~מ���1�PAzMw9���f��\�1c_��c��ŗVF�c�X@�)X%�u���훟4ɝ�V,��{DW}
W����5��	c|�(R�&;�Y0C;q�RI%�%39�_��w^j�܈8wc':�J���/�Ǧu�ȳ0�(u|}1kӺؗ��h`�1��[�d��h�r&~�l֦��\�C��0�.�����O���q�V�f�y�e�mnu`A��P��5�����~i�$���^���Qvv�U�Tw�#��a�5P�5ewt�E���*W�Хï���19�ۋ$�V�
��a�XBVu��Ž�l3gZ�k	���j�����1���<9	�\ ױ�W �KF�Ѡ�М���;����O��$�ʌd`���������t�h ?1Gŝ�+渹[V���k�Y�ac�ʥ��kJG �. ��O-�#�QX�;�I:x�:?��C������7��J�/��c����u��~,��&YMG�åR���p$�Up>%�-��jcT�^�4�Y ONފ0�c~�z�>a|�x��kp�l��#���of���)c��.y<L�@s5��_#nд���<;�*�>)U�]������EsCb��*��ͧM.x;�u-K`�eEp/k�Y�����e�II0f%{�MB�5���묊NO4��"�w�a����o^
�\e����P�ښ'�.^y���u�����l0�G=/�8�4ռJ��Q 
����kȩ
ےs�u��-�T���d�Ą~A�՟oC$�7���2۠�WrJaR�*��n�1i����[��,`��]&Ts��KUUF����󸠿�CU�h��-�ڙ۝[��Y�E�m՝^2�&�4�@g���?D����%%H��^Teu��$X��^��-��� �����7b�D<�l=&}�����}�h�
@OJҍ�MP�����`x��ʸf��d�9��bl��������'`b�0�3�����(�/���#7�'���'5J*A�j����2Vh,s{P"�b�P1�nTA�'[�<����7���8�c��AW{ Vm��N�8��c�3*4�;�!�b��y�3#�-���|���Z�e�㍮ _�=��ܱ���mzx�CY���.�1V\ɫ \�2.�B�ই-7�\p}��U�*�-�N�o�l+����'� �c:���U�)ׁݏɀ�I��R�����m�#-�4�X��+�㻑��[�-9�[�}�j�yl� )+�N�a.)���Qg
e*�-x'")&��C9�����2�!��8�C����;���d�?�6�j1�zHe��{E����hI��9��i���~�v�7UJ���n��q��nZ$�S����7���C�Ȩ����w:�+�d�S����jD�m[����-�V������*ǯh�?p4�!a�E�/����SM{J+�;2�u"%��/��GQ�]9_Ӻ�q������B�xL%uT����$3����'`�K%�n�MtJc��ռVf"����C'�M,2�'%>�h�PB����G���� �r�`?������J����9�bѐɽ��u��c����.;MKYi'j�@��$?!��u;�_�K�{G�A���|I�eЙ�ѤO�M�!�p�d�`����|���0]���̟Ǡ�6.)𝮗�e�D��ۀI�e�G�
Rw��8��
�߫��=�D�f��z����om�L�;�������ϙ�f�s�M��l�c��B5Ћ�Wm�%�t0FmwE��r�ثi��Q�>�<K �NB�bOWz�Z�\CdM�g�6�z��2~���ȅ&�����6��7��.�Ѿ������"�^sY�%H����q�f����S��ov��"�%M�I�WQUbW�M��e���m �`���I��g��s��q%s���-:\�3��%c�)��C+��
��ɻ��#�IT��d�t�	�2�����bN��Q;��T�S����5��4k�p6[������8��l!h���E���(�`�c�<���N�"#%�>��o��e��u�]��������٩0�P,f�s�.#�zZV���ty�/ ��'�� ���]K�C����WX�K����i�ACZ6!�q���5��i�>R�n�#HG�a�?$�Q�?�/�Mi�'��'�y�u��Q?ʐ�á�5�6ro�VBq�p��)�e�:��xD�9���p��� ��Sz��"�:h~���˲�/���B]���k�N����ѹ�^k���ܿ�zf��F��7��H?0kxAȺΐ�A�70�27&j��1��S��렸��M�����:�p/�L4���7F�8��*�l�f��(�m�[29]p�:���x�1s�+����E/�\͹I�S��U�0�L�U�:�Ckn%�S�Rffs�`����7x��E!��E7�@@�V+�6�4JY�w=ܟ��ܢ���@=�~\���������qͻv���h����|
�F�����IO�����	?Mu�ܯ1�	V<����_�1I'���m	�%�[
eg�j��!])�a�C�T$W�ٿ��p�si�ڎ����/2�<��ŕ����uҦ�^n�#C_�JkE�n�fm@K���.�7D�eW��W#�7���e�Ll[T?g��5{7��d#�M���\�/�;��ǭ�E�pj�b�w�_��L�`��.-��Be+$l��>5����5��2�rު�`� ��(�F� ߦ;/��*�����ɣK-�_�iT��ks4��N[�7cŞ�j�6!���u\�MAØ�̪z���h���m�oJ�NG�9w=�ċMפ��Dz�T��Z�Xi��W�%������C]�N(K�J�>BZсV��ꙕk��v�#���&Tu�gp+�u��n4������o�6�"�H�P����M>&���a�	S��X��n-�'�ս_�83 ����\R��hv�g�e�����o���~,N��l!����άO_�#u�^��7!i7\�L��F]Kۂ����*��6��m%7OfG�ܪ���+�Ki�B�����}��ۜ��{\VW�J dQ6f#��P��\��ߦ�K�Ϯ��`y :^���!�	�l76F�F���ǆ� �؏BXqv�ߨ�"]31$+p?�g���m�NG�K���+L�t4&��J���p�Yr�fPB���ur�U��{c�`إ	�!"��˽^gV�G4O��	ozД��e�/w��G��9��1�`�(T�e�.���23��������hS�S���ɎJP�MIq?�Cږ0Q���4�=u�K��=`��ޫ��'��V�[ \'g�αk��o��X��<�
���\,��2(M�E�B-�����H�ɀ�!�Q��0
{���P�g^B'�p j 0�W����^�󬱮!���)ҕiUt��%�ӌ�MagL��*�>e3�p?��+#@I)��D�<xTK�a��9�N'_v��Yy�>��A��Vsf ɒ�'����2���M�cF��)"�v'o1XD�G�&5w_��C�q	�#y�*c�S�a�G�'s(wk�ڤ�;���K�ZD�<�D��2@U)6$� t���<��O����#������\���i��w:�-���KEm�"���> �߽ۯ����t��+�u -���3Kd��x�g��BA�EyD_W$�Bɒ�f�!�ebw)��������7�k�S��M��b�uN�>Eh)�Mw�P�{�ؐ�rl
�}�	�
]>
u�3�ǣ��J��#�ML��-�a~F֭'�c�}"U��4�c!C��,`�ѤfwW���;�1Z	�*rptL��^�V�n���ٺk��	�1��s�D?����xXb�V"V�������'j�	�Zf)p�9#R��Qf�V��kno�R���Y�c�+ ����,2�؊��!�P��Ʉ%83[`�"�Dk(\	osd0��S���B��)���5.H��
ĤlҺ��T�V�E,JNG0���M+���D�wl��Z�����I��<2�s&�MU�IG�Wv# Nl�6B��k|�����G�ǡ0(-�\���9�-�EH?�����T��;0ݱ��ꠟV�\f����aR?~��1�H�'.���X�����i���Ѐ��]��N��^�%���Ty��R����<gu�r��I�UE�+���`Y�2�u�OG~8V K���Q�G�M�{��F��:�X�����kR�����B�)J�]9��8:�6�r�'C�?���`g��7���iJw�{�΄�N�K�5�A�ڱ�&hd�E��� ��LU���c�f�C�o8�T�j�j$�]���W�S��m��\�Gy%�D�)���C���'UC1}Nxk^�JB���8
^�t��{�T��Z���@zC$��i͡��5w��������W����D�s�����kV�d]@"l@_�	�34%���5ϒ��Y�Z�y䒎�����nN�݃�mŭ�mh3��/2c�0�NŽ`�f�Y��J�J�g��c��jj��?�Y[ي���0ǚS;�����܁�p�bH����jwayx_=��5�M��q�dfw^B�~�d^�T�u*���<Q�q}�n�Xgb��������fe�]�˃tH�j^ �|B�)�z]'���| `�}��L^�>��6�j��ۺ�0)(vJ��+v��p�Q���h�ZU��Z�ܕ۠U4�˪��D!�\-0#��+A���Y�2t��lV64���_� X&�궒�h�"��/��0�m�4�Ճ�4��p���Ƨ�U�S1�� ��v΅$���ê@@\���#?Y)ҞwY|ze�Ȑ����a�e_E�E($���گ�Ι�d�u�,9���+lO@y�)�l���sD(��(��h:�L�����Uq��|��{�=�$����^].�8}�C$�,F�6�Tȁ&E��)���ջB�C�"�&W\��Ϸ�KJ��ZZ�0Hj✥|�����J���J�"�qe�X2�K�E���a[�SN;B���K�Á-�KR���i
�P7�57C,MEF7��&�0��ϔ#��u�V��t�<~�H�?����
�a�u2����s�5�l���*�&m�u��!kF�f��U�^�My����d��쵕ü��]�3@�~�SV*3mV��E��#�ͳMgu�'� Y	;��s��X~z��\D�dars���Ow��Qp����_X=p`��+�2dIә�\B�o\�j�t��y�E� �)���FK�E�å�U��yA�Ds��wa�}�Br����;E��@�j_�e
�|I�u�@yJލ;�n�Ʋgmo�M;-���b�|z��[���_��%T�;�3hj��I��p��oD똘�Ơb�Ci��bNW���={��2��h�d��&߃�j���Vȏ�h�9�tۏ��c�A�÷��Ţ�]2h�����{��������u=F�bIp�m�&��Α��<���W�t^�H���;��vM�╔�@"�&�II�.
��lm/Fv�ˈXx$�}�9��8fʑ:^)�8�?_هY��	�i�\��L�ѳ��V���/nO= \5O�q[Bk� c��x��%�o;~��L��/0{6@T ҹ����b���&ax�8�
����9�ے�_b��|B1�j�veUb\��#�&�����y_8z��A�I00�mz��
��8�+܍c܈�$�p�u��f�V���?�)fݾ
jFJ�_���;��\�(E�瞕�@���k����?g�x�5؝�u�8��M>�	!Ƅ�8�R�-�U#���K��8F�@=f��=,]��Q��S�ῧ�7�.Y����-b�����!̮u������JJ��^6��Ĺ�ʪ�S�����,B �^'v��#�J�@?�pk�@떺�������7����o��� �;9�3j�l���z�5q�GM���I�B�ױ��B����ߔS I������G�h��Q�2�d
l�@Gz0/�%���簃XT#�	p�}שb.o��>i�!Y2}ۣ0��j.�ȺKw��UY�ԶЫ�v�<�.�Aхv��ڜg��; �l𘠭��Z�}�r�"��?�	b>��F��~��,����
��5(b���ⱴn8�W�"G����xFf�X�V�t��d몬�u!�B�e��|^�F���`�nZP >h���3wX�S��S�����^�C��Z6n:�64d�0�/���OA�}i���~�^`*H��@�o���q�UCd=���'��Z�P����[���w�hh��A��z�o�^��ˮ����N􂊡``?T/镾LI)
kX�k�cAG�XoAord�m-M!�y�L���k�*�p|'��,{�a�����_�ex�F+��`�H��4����DA�7}����<oZz��9<��˾���c�������k�������1������)5N��.�	S�=|���A��0mK��(n���-TQn�O�]eX�Xxڜ琯-�d�Tu������_!0�9�;�I�F�۝\e���#��Mj���}�0;	��D��R�D�����D�Lӂ�c~��MɽNCV|G1�I����Hy�g����Y6�~�i�ف4E�����ئ�{���\c㍂�<8��L�Ԏ�"��Eӿ�E��w��^ƫ�/x����
w+�Z� �9����9�a����0a=.��*SRҖ�l�:'*U"����ܷ��{T)��.}�%g��MI�Ix0h��<=6\�w�zs�Fsv�&�	�@�񧪾MrO	� *q�bi9�on`q˂2��H��Ѫ+�H6�r^�))�J���f f~_9о"K�^�b����t�(�������<�9�5���:c��s�#�i��px.���rS��h���Z��QY��Rˀ?�*���14��fv����U0�F�K��U7��LȎy���Z�(�j{I����yK7��k�Z��L�c6�΍���{�QvQ�����k�z�> H�P}s�2���t�����]W7�������"�:l�9ŕf�/�Z$�N� Y���+���Kdo{���Y�8h
��o�sF��E� 	}�Ǯ���Ls\�.���d��g.?�Gյ��H¹qv��g���|�	�i��=�+����q�*��\1t�@M����"T���&���x�!?���B�g�ru[O�Z���U�j�ܐ�|�֙�xYi�Z �`0���[K�:�$ǓA��z��;7��!�)�������0�%U/�Z&/&�ճ��U+i��K�),��S��qR(��9���';B�H�5�>�"��}���;�U�G�ћ��q���u �����5&ĺtk��kC����tL�eU��2;]<".���ݖ�5;� +#Q8柴W��;���\Ad���P�����4��ЮɗU�j�m�@����8�7���?�Xd�"���INv�gL�����`�3\���wa=c��
S\�:-��2�	�(|�f�c���?��p[�Ğ�����[`�t<~ž?�6u����$:�����)�Y�cw�E�+���_�+ٍE\23ˮ���%�s�<c�D�YĀꨎ�u���@����CD�_�6�F���]�L2�U9��t�	8�9%��E���G�G ��Q�����>� �k,��K�1V��f�jv��7�iI`n>O�0�?�4u�#܉d*�uW�p�e�]:]y��e��х[Wm�ҥ�hIy��q��^�GY'6�J��>Z�d����P�O;VZ�k_��
�k��ɜG ,�֘��(�1w�4Y�z��:�J�Wq�JMs��9��?��H?I�f�VwVڦ�<����~�.�w��hQ-���P����Ha1����7(�rP���L�(��p���%5�Ķ�ق�ۋG�aD���4�0Q�/���E�,9���M����1�x
�#�ǆW����z���5((�W@���X��h �@�r�:?G߶��)�CAX6D��l���Gj��J�q�;:Wb�H�͜��t�k��g���|T�+�ς� ���֋����M$u�1�D#��׫��x}��%��I�G�ş�ynS�ŚZ���8�V��_79c�-�2���iW��풏p���}�������� ���L�/�a���:$m>l�Q
"~��� ��2�_LgnocPY�N�90 ��;,F���������cټ��H�� � zpj�g�@�Q����{*s�K���Z��cۘ��Z�'Ɣ���\jk�!�fS3^+�&:��7M�B~���^Y�B��$E ��m�4��)��G1���=!�)�ܙIb;J݅�8cv�pX�Ah�3��0�'��4�p�2�WzJ>�L�'�8'�%s��ϟ�f�����/Tf�g>{8�*,��q�X
�Y2<�i�Ȭ!&��_2��
ǯ|��-$ƀ��M����u�ŕ`���\p����%�r�Sנ#)��v��]�lA�����k�؛����%h�R�>b�pGC}�?�ES�۴~=�A�4E���ϕ�v%aO�=K])§�t4;o��}k�)4rl8j�D���y<K@�S�ؒ�l$�/�֤��^��m�F�~%�y^D���e�,usC����cW�>n��D����g��1�ޅ�BCz��X ih�9�t������e�'8�y�i@B����nKq�7��ã��-rI���P0�'�Y`��D��,������d>�hv�GQ��P�t�%��e(Ģ��XOg��"��J��廅�
��C	Wk�쀅6jj�����>�u�2��]��J˾��3��>Z�]��0^�[����kEvkK.��aDn��=��k�������gYx��*B붃���#>���
h!J�QI��M3�ᆈ4�/�����kf�����@u�H����a��^�5KQ�В�}����b6�9��g��r��"��N��!�r0��� q�ѻ�h��o��Vw,�ϧ[�4�ӧS���ȞPc��eYƁ�vZA�{e��u������7}7�9 ��6Y+�i4��*�sC�x�"�#/�8}8���'Y�y��
�	�"@/kP����]��`�-�
�qs�oQ�[��a6����(I��8o"��ՠ�+y M2H�3'��E.H��v��Qf#������?^�b� ��XF�������I�62�M�J6B�'�������"{��W3]���ž��s��&.�$r)!%~n�K?c�#�9yv �4�)Ⱥ?�ձ�ҢZ��p�N�r�y-�
Χ>Z����%8q�g:��RYS�%mi0�z��������#篙inA��V��M�������N�V�wd�MY��XBA�ՄdH6�zDKhV��9B�xm2<2	W2 X��S��~sSU^�2i,�a9��}��a�Q�9��"鷠�^�P�?�����-�3���ɚ�X�Ʒ����Za�U�u,����C ������A>��Ã��/�D/P5���ƅ>�������/�0<�G���̅�<S��0��Z���2d5|'�V(O|��.�s����.^t���z��2 ��	�Lm�^ಬ,�X���7vA��$&�}A������;�ur���ø�����H)�g�?>nc)�����d.�Y�j����<ηQ�ZmRح
Q���,B�J����g	`�pJ�d�U(E���vw�����-aq.�Ɇsc�5���s�?����M��\H�4���E�8=g&��XbP�t���[��A=��K?��+˶?����e��!��m4�x�ȅ%���}���Q�Φar�/��=�R�I�!���鬙��V�Ѐ�a���/�B�C0�:�Q���P�X8��$�*���	��xNq�fϢ�Jc��N����&�h����F��Z��b3�+Sh�YB�VJ[=P�cNĥ�F��V�[��RX�[1�y��� �Ӂ3�q,�Ly���d��;���nY�����V�p��Aj DU���6Ol��i����|���Db�R�Ԕ�`|����w@�V�r�������@�0��ʨt�l5�.|1�IZ���C	�-����i�؁�����# ��r���(h$PP/��^�����9�O$�U���<�,b���D�k+�Vf���%d��n)� n��T�PR&��ȸ��a�{fΦt�������"�nRI$��b㣳X�D�C%�t�~0�F�P�w��E��H���M��.ξ��Mɍ��P��b��a�;������c�Q��]s0��FfYR:�l�"yL!"Y��Y�zտ#4h�~���Lv�r�E��n�x��t:���P=%!K�����7>'�ԥ���]��<	�T-�m�����ꤊ�Sb[*�˲	��m�ވ��rT��6�>�gǌ%��OeL��ʐ�s��x܋��m_���3|CK'�1�Au�x�)��V{�λSr��!q/5Qp[���38lB��K�s�*�&���Wd�����f�ML	�y(�g`��Z�.�ȋ�-x��o>DX��+�[W�p�Pf��{���K�.�3D��JI��걳M-Wc�C���x�ȍ��-1g;Ae^\U�7�Ǉ�Y�����-k-���v�������mB_��H��r�Ѕ�G��N3r�e���p7<�*�6��p�����JodR�x�8���#e���{�JA��bX�rv��'��)8G���-%�T'áZ<�R�
���(��gރ�X�&�Y�j������7��e�픏��S!8-�+�EJ��j�%�ޚ��7��3xa9w��nXP��.��+�`�	w���;X����L�s�)�du��~�l,M-�i���^3XFh�����YG��oe��?)w"CI��K�k��e֠���&z{c}�;m����|O*��0fR{��Z�*H7 9&D([
>f�*��.{΁�>��`Y�Z��;�d�/���u��Ǻ��i�Gx��X��PR�};_H\��.�fY7�ȵ�!0]/)?�
���JΝQ��O~
}T*l�@q���o�m;c�7�H~��d0��<� ;�	�w�1wb��Q*#�ޤV�Wh��7�ŗ�yM0�̩I�)�w���s���-�g�5{�����`$Rw�=���������R����(���՜]���hn��?���o�z^�/��fk Oy��X�9�q)�w���K� �ܜ#��� �;!n�q��s0���1ĴM��f�4!D���w��7+���W���Qҽ5�K��;�$A#j*J�S��#���%�"TN���E?F0wo�L,Clש�k�9Z��W��e���.����AJ�C��KP`��&�So���1uI�Ο����׍��e��rQҾI[�Ϸ*��v'���t#Ap�z�g��}�Bup�;D�d���_?�B($M폒y���V�]�>!�6qM��IGmf3<�m;ω�0�����KL#�v	�;B�")+�gDÈ�g���^#����}ɂ�q`�����<d\H��?>��¿��Dl��K��dڠO�����uR��`~.A�ˉ���+翸:��m�L<�kg�x|k&�)���I[��p��e�|�(��n��A��BȲ��e.U��0�Z[Y�(a|'�f��{p� ee��ou�`�1��m(]�
5$sC#弗䖁��,H��3�u�̻��#!I�k�ʊ]�&�jϒ�B9Q5������#
~�F=>�@�\�cmޅ;<r-�e�˭M�sų�:��%��Q�F�����UF��;H������;B�8���O�?(��	_Zb@~�3�6��^���N�����\���h�����W��,ѳ(�Ѹm�׊���E34�bϿ��:;�|	��2���?��o�/'*+ɜ_��VD3E�k��>��%����y�=o�L|�+��\�w9���~��s2�W3d�RXv����Ĳ��CU	`ד�/\����Ρ)i���3�^�cS��os�A[_�>�~���R�0 ��W�����(8P�<��>�:������A
z�2[�Qg&�}�c:e1[��?Sot5�	�������$XO"LJ��g$�-DKdw^5�Ǳ�	=����GR�@k�� ��P$4�Y��ۿ�%�Z��d�J�SURx鰭�=
35v�o�X4�_�-m�Mfy?�������d�n�5	�I�����\�,�e�!2	F�E(�#�;�̂�DN6�ۉ� 7��5-ʱ��J�F=�ɻ�X�P������c3��C�)�f�ƶ<s3-�CZ1��C��m�w�O��a��g��OE�EPc	�GH'�>l��L�X7k����N�~$��d����H�����!:� �K��:�GXX�WC�B2�l�7/��j�e�7F�݇K�
d;���Nr�.�l�>4�/��u�Q�dS&/����Q��%J�­iH1X�Y����ҫN�ՙ��'&h�4�g��x4��t6ݽ������h݃�����P��Ɗ>�����%�E8�C�����x���������6u&Ղ���b�كB�\��@��fq��N1CE�|H���U;���Ű<�`�>�Ն��?$�sBG�8!j��c�s�=��eba����՝���Yd)7wx��BG�����t\���di)1��_ǲ���!�O� \U^Js�_�-�-���_�~&=QU���S��_l��W")TԂ!�Z�J�����-3E�?�_��QK�j��D����v/�����m[�>��?n�`B��&b�|���v>�Ww�YZ\f�<!� b���)�a�MϬ���EE�Ն���q����u�iT=�x�@�U�� ��w4�Y&<������tF8����)=��ڷGg��iS�E!���Ǒ֫r��}�@�z��_�U�tCr��a#���M����!�̖[��e/�{(ŕ�w/�_�,�-s�ve)��G��<�N������i ����O���q���▨�N�/]w-��Q��]'��)���2�9ʶ�y�̜"<XU�/1������5zf�����|= [W��m5�L�*m��|��a�*�TR#x�)�<�y�wk��[�U�WRB�$7cf�P%�ѫ�E��y=��~"����I�ꉽ�}۵�2f�N���O��1աqF��My���X��A�Sj��L6^����.S�ߤ�c�>+ţ�Q� ��X�Ч��{(��j�T
�����4L�-a.H���{�Z�`�ZR>l:�h�Su�^�=�q��<#�5͔���&�!�_�1��)�e�H�k(��UUP��f�M�.c$Ց�� �ƍ��*��%�������w�7*��cmȝ����3��֠H�u��":��^�TZ��ɏ���j�S�#LBYχA��W��x�02�1HTS
Zp��;���m 4��7�3{���u�8��JK$�ۧ.�Ea�6�,h6hd7ԙ���7�4�5E�?`�c*��5�Äup��7~E���c:'a=�Q���)����ppv`��`���E���XN9�l+�?� �[��:"��<��#_t/8́�bF��f��Ԯ�P��u�	�� w|����@9	��$���6�2\z�X�\�Ms��]aJ��\��x��s iU�Vp�6m(��cԙ�k���z>�.��	4`�M�,NbQ����/��~XӨ���	Ǡm暤���p͹���6�-Y*!`z�cv@y��:~�`�d�iAp�����dy��=}��L�~p�މ�f�����P{,���a�:9�����G���IF�\��2�Q'y}g��>�rI�wC ~ij�� &�驫aߣy��m�����>����TfT.m�����88�<�,>g���Z�V-��	���;�9�q7���~���cWe\��(eQF�����B�D�ʐ��L3�'�����uڽP��9�&��c N%B��|Zj�
�s��rd��>Rj�uF�|%�-��g��C�����iH�/6SM�n#^̪\.��SB�8R��`��6��lGq
fl�����<ĳ�W�W�U��B�����bm�z5�ѳ�C?�����W�@�ws�*sߪ�Z�<���3#���TPOd��P��j�6��
��츎<��{4��J@q�4Y�����j@��d��U(#ku�
v{����^�Dł���]?��u]`�,	q^#�8M�W���Ʃ&��'�G�uJ�B@u���	
3�Q�q��D*�����X��S^�]���"u���M�FÏ?M�+�1O�}�����o�g�3��%f9���ogaHz�	n��6vD�1�*9)G�'�{���V�6',��������,���Y����G�v&h���1�R��ip�h��R�m�%��"f�^ؐ�z`ʩ� ��� %��l%��Ms��� #�%��� �B�dЭ t-g*���Q7�w��J�f�X�m�r!�=Hl㸆�T�Bz+ �e�i�z&�\�4E6�x��zp�ڃX�ݞ���i"�"C�U�3���&��Ѿ�q	,�)ld����(2Q'������=j+}f�ɚ%�&��#+��)��0����$�z����o�[�Y���<���x�NM���)`��c��IQ��B`Eh����:}��&(��5VG���Z�{�+ٝ�x	� �5pa1zm��"l�|60�8�� +��ʯs��M���T�����/��o^!�%��CQ�H�z�� A����k�2G�+D�,y�D��
�����B ��Z�&�K��8�DM�g
��i�hr�=���ӄ`�W�I	�<J��u4d��ZU�V`(�@�Ci���p����A*X�T9�O��31�EI�;ݨ(9�H
 ��^D ���oW��0�6ߤ/�����Y��m��:��y�0��T-|�[�;�cT��#i$W8O��.TӰ0&��[�b�����Ods
�%V�o�X�����3�l2.b"���l��us���PY���Sߵg���ٸ���X�[���Q& 6��Ta���u^3�c/<�e��V��F@����%�Cq��sӱ��@�v>[��ja��FZ��OG�1h�_�[�d����s����Eq�0xj|Y�Si�xcC���o�O[�Q1�tkyv%)=�O�z���,�����M��T/ƫ����&���D�K�������s}�{�w�ԵdC[�e⨗� ���ݡ�!�y�w��);�V�=�7�t@�a�����P?���yd����J�f9^~=��Q��a$4~�N�=&�4J�T����S*b�\�4�P�Wi�S��kZ�p!�8���&�×��A2��z���u/䤫8�Є?���2�逈��}!��^$�0t`��ҝ2�×�����h����r땤��ؿ�7��7�:��.a�-��tTb�Z\:W;�V�.��cr�=8G��m�7��;��7]�ಹ��j����ɤ�S�c���/�>T2�r����-`�/���)�2J��=b;k�T��~�)6���_�ߠ�'�gDo�x2��G,YS�ӎ� �1���d��YE!���ߢ�S�l�<�1��<m����$�_���*}�:�p�Y-Ed{(��Sov��,��I��*Ǜ?8��`���!� �u��3|WvY��E�E:���&��G���j��Z/<T�/m(��98��4�S����"w�Q�Q#x��ym�@�¢+}����&�KA_р^�uo�-�p=��`��ˣ�ˌ�<�����n��U���gM���b�<�]�Y�hY����c�7���W]���J�"�3I�OO{�vz��#d�R�[��|���lC[�����'�z/��~��(��r�9/��&��.;TA��"] ��̓rb�Y����g��f,n�I8F�
�%m9[E@>��0g����]�����l��'���ǰ``�p:v/d��}f|��^�\u��kP�Kn)�	2�:�S����}�ڱ�/��D��ۭ2Y�~�:����ג���,PM�����<�Nt\�Կsk��[ݦ	�	(��m�H.G�E��U��V��� �=�� pd�w^���aӊ�'#��!P(`y��٭�~�� us�n���?m�"�gE�L��k��?��Ԟf�T��d���VG�g��6�&���N�EM?S�1L^
'%ŪoEJ�i�nÀ7���ʜ�3�~%l�a~s-����\���EC_=���Pܿ�YY�r�����Ex܏9��3^�����2{	���v����K�j<����?�_�����G&��g��=�Ps�M��� �a���X[�.I�X,"�h��N.�b/��]A�T�����(ڢ#F����8��ä��c�D�F��;�oíSQ��,Z�����rZ�_&�=�QU��*u���V�8�F �Y7�Ek�1Kc>k�tv�II��oU/s�v&���F��>�����G�S��)��t,���g˴�#��E���40��Ҭ�+�M=�=�̓��[)]O��n��C��B�=�Skg���V�d?�M�@n�a�)_a*}��Ci�@ ���0³��S[e�^�o&������j+��l�:{`#F�`5�α9�J[uA|���]H@�1gF��@��%)��D�t�~��3g�MY��sa��/)��n�]�X�����n�1�o��В��~h��~�7��E�Fj�X�"���q�wk��T�:�$)�!N'�r�&�6mg$�RT[�pڅ�
D���%؎U���LzŨ�q\^5ȹ�"��P�Ҵgn^+T�>BA�Kx�-R�����/<�"���*�t0��y��_(T�A��d�v�SeZ��|����)p'��-.�I]t=�Nc� �����"Im���tӶÝ��Ӣ����
��Ѷֲv1����hg�0m1�#��o�0�֜-P	"���^|;Eo����6�s�@���%�_�с1�"���@��,5��S��l&I\ARi��q9K�V���v?�	�^�7/�V򘰜1� g5��� �} %�����/�E=ƃ�%�m��6�FT��-�ͮ�Z`袨��xL3C�܇�69�r�.����֐�rCSJ?&'X_�|(�\���X1�(s����˲>J��;�k��4��0w
Ճ�BKx���#�N��3:���@���f�k�Q��t��<�l}Q[}i盓�@�/Obȥ����D��;MAT�y���\�V�G׸aZ��T����,Y#䟎���Q��9Uj������[���d󾌡�x�|V����������QCOJ��t����hx�#��uT��a�^F�)'t�<�1N��]r��(1Z%�X�fɓc2��|��J)�)#�GO��:�T�y ��Ds��8r*Y����53�Զ�yI�@���G�9�5��.:c�E=?���&�|�jk[r:��������0q��ʥ���,���>I��"�g��ہ�=6��� �ե��S�|����JS�B�R�-j�X�  ���%���#>���chȜϓ�@N�d`K
�Tb~2���	*��� �B�o=}/d��n�����)��S��xԏ�H�X��@��m�&&��K×%�8���{�lԪj�Nu�}���!��ػ8�{`b�fK[�O��/���oR։�w���
�F��5���&~GY@�ѩ!�axt�@:W8^N'��y6I��6n��B㴸 �V�k	W�/-%���ʛ"��-��Pz�V��G���#p?E&�}�z���ؕ���њ�����3z�Q��(H�2����]�H���jc����̘'��~�LAA���ݙx�O ���*!ƛ���LXo5��{���4�UEq ���/�C�����zy�&�C~���dvZ6�14�E��&z�^����I�W�Y�s1��I�a<q4�P�k[�U�6@tn� ��`Rrq�^��h���m@9�M���ۤ�iB@Z�Ω��H7�2[��V=k��k��|OK3���v�u�cWf�s6%Q���`8�j�'{~�aOR��J���w����n�>�<�;)��L|������I�zt�V��ZQ<L&:�k�Z�~O'[s�	�A����$E�ff��I��聕�~~�_}a7s'��Su[�+�!��R&�c����[��_��҈����X0+���Թ����<�!��Zq�F�U����ܸ�j.���>���>��/������-<�f�.{�dJU۬څ��O���>���)_�u�w^%a}����q���jᛁ~���t�	5>utf�`vy�B�k=����Czi�P#vB���o���$�"��Ta�ͯ��v����Й	}��mzB���'��,�O-&F�:��ُ������^�2=�P��`��u9��6H�֋���t���\�Q�-I��a͌M�>Bۢ�+�Z����������R	��L%xb���s�;I�gb=Ҏ0�ـſ_���y�dF�h@H�
a!�,ϲlo��v�]��w��;_�F\�ΝV��|`1�.��E��+KQ::���Q\M��}���B���B� "S�����Z��7 ���D����ܺ|� �Ǽ�*��4a�:�Y� ͧZ��Xˑ�(�F�A���%=p_W��?�ꢶ��9k�7QH��Ϥ_w��'C|7�7��̙���(�^C�UXבq���?�o�	�v���BC�2��j��$c5�+�U0�G'�Th���j���a3�����
d�YB*㒇��ڈ�kI���]}bj	�8��,��G�˫�}�D9��x�~��"�p:+rԯ�\TcߟɈ��kqR��rФ�� �N6F�=V���yG�֙�faN3n�F���;Y%ZJ����2� H$a��u
A{Nk��$"�i>A�o'e{��������36@���D4����|��i��_�n�&��F����i(eǱ�T_�O�=� )�؇��)�R���{>��ٙ�$�xx<!�A��o�FS�M�&���#��T�
o�����o���+f3��̪�J*�̛4X^�W�i�m��A�m��_�kX�8��t��c�v ǴLX8�,�D�z��`*�)����uq1iM�'�-�d�V<#.I:��f<�[?T��׊#���D��R�ڋ97ޱ��N���K~�/�L�Fz{�����0�c�w+��t7,ԅ<}�vk�ן/��QJŃ�0���6�t��y��6j�����<@��s�y05R"�n0�[��G���҃�*H鼛'u*�
����V(��U^�]P�6�j�"�΋ �y�y���cRy�G+sF�59Hp�NB\L�Z���f��cl9�*��+�4)Kz�⺟���UcB<X�?���fH�c��$/Y���S�_4PEۘ�_��O�Ɖ�z�<�w����ĵ9'B��|5
�Yo,˺&�nP�O��o~�	�S'�O8�!8�� >��.ծ�*�|�XV�}}Q�9����I�~���({�m8�Z����][��}'�o�pk4%�kH�w�S{�1��l�j��%=�1��N5����حoΈ�a�ѭl9��ގ����oG�`x�Z�	�d�[����W֐3?���q��a�L�Ǫ*�7&���!`_C����A�H���!�)�6̻[2���>h����m�-dFr��bv	3���+)�Ⱦ��~�AK��f�Rn��M���I#e=<�"ܩ"J�gʆ_~��ϒ����6s�W�g�����kby�+c]�1.B�8�i����潹j� �z�HͲy�4L��A�-��7��>~��g���F�76�I�[�;�ޑ���Qz)�*h�N82q�0��jΉ��y�r �njD0�z���ւx�NW3$�C1{2	��Y�VJ���t�������&�숋Q69�Q�ة�Zam��\eү4&�C��P����m�����A�땞st�!u���#�ʀ%��)�q���!��ֹ�:#ϟ���u˩t��(���0cĀg�ܖ��'�G�a�Ǿ�'��Ɍ̕ŧ-KK�\��%�U�^k&n�����������}��i�+RTOeI-9����[=e�MrԠ�f�<�>�=EZ�|SE��IR}��~0�;'��<*ߤsM���*T0�2*e�+�J��b�����m���A\L��
��ޝ]���"�?c�(���l�J�� V����� �x���.���Q	c���a7g�dy�ܑFwS�A�����������%����$2D)��g+�9��A��z%8���q?��72&��G��D�>=3���;���N���W�w֭��	��Y��^y�#�▔�y{�ݽ�&�o�~�
���=���G�ul��l<yF�W�t��X֥N&3���+����j�;�~L�g�y�����fk9���t�� ���3vqA��:�-M����v�^e�ÑQ���a�۵Iq�$+��TQ$>�f���ғj���݃����阰s�$ݍ�c
�h���㖀�j�'��K�)���y�p�7fR��dtǯe}Ei����r�	Ŋw,�-�y�O�r7�	�{#��~�t$�d}���$�:M���]\�,]U1����F�ͱ�e:K5�d2���+I�	q��\����6�qI(/���a�.�'="�Vq�a�c��y��aJ�i?z��!cȷZ�~Wq�����3�]����]��$��JZ�O��3/1܅W��b:����y�HJ�X�ai ���j�5ik�م9 ��6��w�P;�k�q�MG��z����v(S-Pl��0�xʨ�Y5e%�g;ճ����x�3=J�p3�so_�$Z�=K4$"��Xk�#���b�m�,�Fa��ῳ�U�����*�^��(6D� �Л�T	�a�@(�s=P�`/|)�����|��q��o��L�Wj���ٰ}c|1�� V��
2����\z'�~�1�*1�+b֍TL�@���7"��$){)U�#U��|�c�E*��H?O��Y��١U	+�?3U��a��L�V�J�v.k�/��Ag����J�'�ӟ�����JjcZ�=�2\��;�4�x[�P��"�Q�v��{�w(V/��2�|Y˯��;p���`k���s��D���v����t'n�Z3�^���LSe�u�@S^��=G�G��B���cB��׾�dXʀ�M�E���i�Ƶ���:m��a�R��撣B���#�qjǏ�5�" K��j��_�Y�/!h%�O��0]w�>�홙t�,�Z�?�	�[B�@hL�.��ڼm�Z��X�P����<x�R�	�S-��ly맃�c;�r�`{x5_mjR�����C�m]� ͯڣ-yn_qO���e��i-���Ei����GL2�m`q��:V֏4-�5#1:�-�	������]Z�RA�u���D\1?�3b��4�����^>Ha���
?����F_�E�J>��dB�<pD�Q�m�՛0Q(�P)�H5���"t�O�̥�ݩ(?���!�;*p�ft~�4*X�w�c�I�קaW4e�{C���Vւ��e)��a8�+xMEg��%wK���A[ 3��e��f��/c!3��O2{�L�4P6Lp����G
���M�X�q-,`�'y"����u!�����C�_�o>��LXj���h�B5��<ZW�0ɛ�x3��&��2��1���_�_z<� ��`[XJҙE�_@]�\F>}=��G{�>6hĕ�-����&_a�p����[�ZNW�G��Ew7
�ԕm�s���TF���@ʵD{�aT��ީV�vr����m��3�'��j����z��i������=�f�C���q�g˺��}��+��WB�����G�^O��WM]�ِѳ�#�q��Nz�`?�;D]T��,z��0���o=1N��0_���a,EI�T�0��>���r��5~*L=�5�K�7$zUY���}�2������$�v�ɀ�@T%�}IGE��X�O	�,��!$���\���b~��V�U[�t��Bh��c�c��2�z �@F������5g�U�?%�`������;�駆2�������n*��bO[��� ���Q|�{��U�X�ޡg��Mc�l�y�����LN�q�y�M���;Qe)z+�Mwb:E{}`o��o���PZ?Ī��mJ��:���ϫ�C��T2;�#Η�"�A^	&�x�q��b�І+xO�t�X�q�_�� +�]�C���?�3�T�vWW����"'�F��ԟ���xC��e��G�Y|�`���;��Q�|Mzq�T;�P9U5�"�U���S��_.�f˛d�r��7"�ҝ�ob�N��߈8���,>��=R	(�q�G7�fEݠ{�BZ	��o7��5�(z�hy�lNʿ�h��&���If>)BD�_�JD��!D������H�k�!-i���Tnۗi4=^��?n����$*5K �X��K�Ҋx9`��O���.P̰P�b�2�*~�����ݿ	��[:����"TW�]�ϯ�(�����P��P|ˋ|be��w�v���BэX۞��T	.�݁�U���~�؎��]˶�`��k����k'�oPзd�-�ȮډH]<��8��i$_fb,p�S���jx���(P:�����HM�$�GP�u��ߗX�d<#*�URg��ܠ��x���k�	�-��2�K%�i�T��^p�\���u�c�9x�/����X�K�dy���6��-ԏ,� ��Mn0���Mfxj�%iWvf��#!d�	���ڹ����8�}c�[dz���iolE����]aQ`�X���w��?��
De	���`U�r��D�����A�YuSw�dO~:�m@�$/3�#��{��̩��F�xc�ˎ?�ٺ��/���Q�cM y���}3W��m�a�4��L4�p�-�����ϰI�IdƯ���./�<"܀�#�-�UЦ���t̋��)����4�S��d�;~�h7(r�{ۖ�C����v��Oi4��3�Jv�ʼ����,'w�:~�E^�Slx�_��ߞ�c�u'�D�2�%���D���kh�O�[t��ɄE���3Sn����??�'N�X8�7�o	<�)�A�Ix)�
�>��E�4�iv�J4A�$gb\�P��\�U�=�^���o�cG��1�4����3�)�d���x5������Yya�ұ����6"O$y.C����Ǆ�e�U��^,�����%a|����|��3�_��:ئЈ�E̍v�E-�4-GD�J�+�ҵ�(u�;T�Z����P���PŲ�>p�0�G��=?��Xkv!J��50�W�������t����Wa�h���[���']�!��0��	��	b���6ܜ!	m@����]��]�d�p���1+B�,�<�AO��O��מ�� ���ZjC�����o�����8'�M��a_�b�x���͋(�	�|O9�{*Iǃ�`���7���?�>���&����Jf_�ӗ��&�Et��X�$̀&�;⭀V��:4���ær� �k���-6x���H���;�_L+�=q�oQ `F��6�W0;�S�/UwP��uH�]�₼���ǐ~h�c���aѾ<�b��v6aE����Qe���������1	z�s]%�N2�]��)p�gD�p��;�n�$�����~%�
M��ON�1�����h�?�xD!s-��m#�?��ٸY�+@�M���հN���!�	L����|���V���k{��~�,�D��C��U�*��6`�Sj�hU}]�p�j�C�D���8&	���zDJ%ӏ�hVV�%�bO��7��;`�����fBg���� �3'3�bca���j�BP�<��y�=ae���e��N����v�U�����ŘF��UuFک�<1g�.h�0�;I�l���.�q*<�[�IX��$H���LᲓg��h�&�d���#��!�)tu8Z�.���b1��:T�?V�(�$3R�Z��V���ɗ
Ŋ��Ȅ�j�uc�W��:��|���P���M���\u�ܯ�9���7@�ly�!4�l��L�#e�@����|aj��+ ���+��N�w$��Ch	�Y�P�c/O���yj�E���4�)�g��\�_V8⣧��)O��K{v���g�n�!��zs|��hȡlT���B�'u&6�^o������Uh~Z�9Z�l 3i"r���z���&�7[�)��ة���^ݖ�Lst��g�a��>��8R@-f�����}q�N���%՟F��Ld�ꆱ�]VQCu-�J4I�|ܧ4�S��9k��Z)�f�u�E|��#�FE���v(�Dw���&=a2�1~�����}Q�	��Ņ^6�rQ̬�ˤ��:l�
c���M��� �~�ˀ�AK�|T���D�Y��� �DPAV�ŞP������wUdXZ�?g�%��3Q�}������>r����& ����P^���Gn����[�'_�{(�ݘ.krqUL�jr�nB���dG@Zv��� �&�ѱB	'	;�P��S�+��K�{��.L��K3��,6b��m,*�S�c���c�\��r���2s�A�kl�ҹ�m�O�HAOT���&@_�Z�C
0�I�;�����-8��˧(_�ઘ�:��� �liN�����WLr���m�;�������#պ���󊆣{��!�{Y)��.��,��,a<;K{!{r�3J슦��k�3��� hjeHtFTw��D�Ĳw���JTk��k��Z�ǖ��bn�=���9�~�PYKě�`s��6�s�F���e�DSX6bd��'�D��LEL�MlRUP(`%0���k����6�6��p&�Bu�;��V�R�<n��]�� ���c�:-�<���@ѣ�=`j�VU`�ѳ��Κ~�,V���������6�$�y��x�o�	[�ӮG��%F�~�2��)*[5�����]>ɨ����}�!��Q�3��-��:��y� �����WTg.HYF�U�G�(��)B΃��a\�duĦ��@UM|��˞]��0Њ�pj�z��:��O|EA^���O�:���+�L&�|�[�+��Y<�@�	���	��Nl(^)���{8�QW(��C��^ť��=�'���Z�Z7�KP�K6%���9\r��!�AzN�΂y��7ʸ�f�l(�AJoy;P�4/$W:�×!�ZT���S�M�N�}v��ڵj!}�Gڂ�l:�a����(�:jh,v5��/∙�?EG����Kn�ʤ¯.UH�Yj�P���sՈ���i�\�m��j^���$�J��Xi�}Q�O����eH���T�������~hP/V�kGb�A�����WIk����L�џ9�<mx�TN�sРB��/Hrߍ��3m�w�St}E/U1�ҹ���Y�)X���h�x�aj��H�E�6QJ���4�N���:nM�^�ڼ������L���q���A?����*��U�;Ed>�.J�XJ�+��=�����R
|PXd