��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�x}��j��S�b_�)F�1�(d'Â,L.��ꙺ��e�˭'�{���)�Ilf\�@,�y��Z�n�X�D�P��c�����=���]Od�w��yD.΃��o�N�o?ղu0��sS^�ۋ�0�[�@�i���W!��2�b�Q��~w��y?����N+��D�����Y;oM�8�u�*�i���&)��9q���t5�Gcٝ �z5⓸g����6��?�z�N�#�E��e����kל�P�ؘ�AX(S�8��*z	dG���ş0�f�,�~������gJ��d��& �I�k͜�kֹ;��_[���]�]^��pk�:������Eml�/=Iw�0�^e���ס�����bN�?:�|��+�-�Ѥ��4�B�3��x�EK��*���cG1>^��-)<���64xf�J�Z�����E֩G)�+S]�rX��!�[H�ݧ��>F�v8䜁�>���+��0���r9�R�B^JM�1�Ҁ��p��h��Sd��� ��m9������(�qB׫�T�o�K��L�c|�΂i޻	�!5Pu�:�!�B��Zh�+�l�,*�t��i��D"�0Xk�ԩ���������0��f$�ne�f�+��e�rf�z�.z��=��ą���I�.�_��_:٘�|�kz�"K���ԜBrzpv�:�d��O���̕�����2>o�ٱQ;R���Ď�?>����/�>V��<�`ڹ���B�Z����[,������cf��H��Y��-�\'`�*cC�Bƙ_�޳�-� ��.ݛy��~��,~�zl{�f��Hw�e�E��E�m�F���\}+���Uv<5����F��A��p�~��
^@^�\�OFa�I����n���lw��Q���Cj�������L��ة�-d�$.��)J�,�;�+���TN6�{��`|��h��T�%90��xIwTC����n?ʡ���ڸtFO����+g��[_��3e�ml�(��㮦s1_��5*�	��*嗉��3W1�d֚A��ʵ▗_c��0����Oc,�:Щ�}�C�erT�;��-f�׽��#R��*���B5�xt5s�"_زpb���	�<��5VK�^�%5q��K[jDW��sV�*3�)��a�7w�8�� /ſ�NRn�)�>�����r�lk�٦������5��Y|���r���q�	���J��5�xh��f�C��fP�`aV���-���QJ������o��1�۩3�j�,j&hn�m��K^��pd�Z�CF�j �Kk$*��wh�v���L�z�/lB�����"s7~#2�����67l����?�g�5�*}XIm!�iV��bbiD=�=	�8Uu	�'�'�d�́J�E p��;��=��2�^�&�^'F�	U%���!�z)N��ǶT٤���l�8-�qIrfZ�/��5�����q����jg������M.�{x��a��������HV�e�S�::����i�77I�S�Ѻ��::��:_��FA�����?
ٷ턯��?6r�KT]�/�p�>�xq�;H)��m��a�N~FM�H �I�RV�l�&����<=���72�0���0$LKz"����!x�o�
��q��`��G�1������X����R1_GH�' �Q�R�18�^�aHN8<�3;S�T'Y�F����%�{�G�Z�iN!4lx�f�p�I��$���{��ʫ� �ck����Tn/��ש�Vj�P��'Z�rv�B�7��亮E����n�ݷ�rF��jm��f��2�Md8P�2������Kp�_aaA8eGB����M��𤽛m?3�>��O/m^Gi0}��r��"�@,F��� ���0���\�+�5ףv� k	X���O���x�(�\��p2�d����%q�ظ��p�P����ƛ�8U��{���U�('��ń"���ʄf����wDkR�Ģ��u!�����M䀈,����L�5O*���XĈxm'�U�jd�$��"?lM*�VBj� �' m���6�_��"{���
�H1;���ʞ�^��UmU_���C���,o�u�U�=r~ߗ��\�j�YQp�e��R3�V�C�To= B��A�I��275^L���`�7���W�W:���^�Ǜ3��v��E]|a�e�?w5����j���f��������
��Y��mf�F�����g�Jl�6n�8n���%߽�[4DS�����x6"FB�5��ui�r'!ē��Q Wܦ�4��F�e�m��j���ƷƢ�"�~GNvi���H��ϊhf.&�?�#�n����R쇋��@��L���E/:�M՟|���6+�o�G�A�����$F��愢�a�̄X�J�$���x �'�����='77������O�bNV��9A�.?�
v��c�FH�jQx�{��<��4��ت�9'��A�/�
�q�gWd��$�8e�K��`��-�)mXI���C�U���_�js~�������/�C�hqR��Ֆ�y����DS%�� ������.����U'dq�j�_��n;�]���;�LE�O��t��A-Wh;"�T �b��d�]=���b�0��3�^��F�&���j^��i�N���[�e��G�D*mj���ZP>���qv�D)�pM�;kc{._�:7�����}}�V���L�+ʭa2t�+��I߶���l��X3��Gc��E���E�^:�K��Ch@I�.[P�;�L�@�hK�R*���*c/&<�LjF4-S�i��KccJ�d���Fv6�vE���9)n�M��h�)��h�Gb�L�&u\�/Z�+�A/�Y1��1��D�K����1<C���x��6Prt50j��G"D=GEEǔi���#�?T��;Yo<�ڻ��� z�"	Y[��ϸk|���@% �@j��A|�6D�*��>k,�ݖ�ىO���|�:,-~�k�rX��ө�Xr�"�3wr��g$1��.��Kd-t�E��7���ܕ��R�k���������َ�?����DU����<�b�o��V��FH��\��j,���@j����	J
���&NśD��{9AB�Q�î$WtEf�3����62j����	���,<�iQ^�]�ٯ��l戎� 	�4~�:�R�_U�h�cϳӶ��A%��LGI���Z��y��u$Ds	��|��H���mQ��*������P&G߬fi�����O�ŭP���yo'��9Hor��nq"�Ru'�B66����:�Z�[Q����vB��}T�����?ˑ������^Kw�ٔ�ɺ�e���~B@�h�eV�9�c�0�o[}���n���y�5�)� Z�KUOӨ�Z�m�l.��8B�+�΃��a�+��:F� ��,�0)��3��URQj�o�}A\@�����d�((|��g�MN�����W:9�M�������>V/E���J�o'�����Ϣ[x��˿�A�%B��m�67�Z�u~��٭�x�xb���m҈I����	ٔjך�`7p������}e̢ފwD�����������~;w&]�CR��vV^��[q�� ���!	p��o��#�^�_)������
K5u������`4�CDl �lai?L�y��3�
���礔Dct�b���T89·�G����U~���B9�3���]�����|�3��*���9��?`6\���;i��XGV���C�w�h!㘫{Kw4�G� �v��r�h��gӅ^�-�
L�ܻ� =x�����
J�bJݩ��������xU�d�}��z����� ѲI��r�2�[�J�� ������h�t͞]�4H@����PO��'�9.?��	8�ɷ[���ZK�XT9�K�Z�ϝ�Ƨ�9��mw�B���Eg@�L:�����R������?�Q\[�E�u��E�枕�����yی�2��Q�:�ߗ��~�:���,���5B�Wʾҕ��|L�+�l�0���v�ִ~���Sn���Y��}�õ�RT��:�ǰƮU�(�TM�М���M
!��$�Ӌqx�q��L� �o?�J�0I~���ӟ��,�6��
 �>�@�Z=�5$j�σ�@�-kH���VEO�-}������wY`�>�z�\tѪ��8�.�k$����r���Z8��B?�I���k��_�^L V�V,�`�;
;p�_�nzH
� ˨})�S]x�iNb12�R�o�|}�gd-����{���8V܈��ǀ�N�;K�,������R2`V�/bA�,�|�1� M4���4E2z��_�d�ϛg�>��)5�����F%�Z�o[K���{U�)��}�x��J�ƶ�S�f]���I|s��9�bM�zB�8b� I5� �t��;�A�E��U��?�yȹ�'!��h�K��뎤�+��W��]y�;���N��٭�f�X�t�ęz�P�N��32r�b�?�Kܿs*�7x��a�#i�������
3C{��/���Ü[)<�O�i/&�%ԑ�
k-�O� ���=f%����Ce�4��4�ݬ�^�L5�J�H�,����������v9������7������5VI�
������;��=�rÿ��&�5O�*�=��D4]y^�r6�Y�'�Mpt���)���>��)�<��E���N����eT�.�W���&k��<�Z(��d{A��6�����yֽ��8��q���2R�îV&{�15����H�tZ/	�p�;�<H���H���'p�cd�s�0�~��ۥ��Z��/���T��WI�ۺ�M�`������#Q�g�cĂ�b1-�P���U���O�-03Z�T�kL��L�{�c�MVB�A�|���|�]�XZ�|�]cZ�!,����+����w�>�ʙ�`u$!���^���Gj�G��}�b3:�8A�"xy��+ŝ�����(+�o�x����Q���c�F�_�t���<�j~�u������;���^�Z��3�gÀ��6�w�X����*i�-G{Vk�� �1�1��a~⑅�a$|:|����ݢ����GY'�<
*P	���d�%�$?���ȟ��u���4�v�n��[X�k:V!��_�,l`9��:~:�"���#��dƉي��T-�ɷ�r������%�t���������CT�EW9Vp���xd��v�1�W+��@���Qo��edآ��4� Bm:hٲI|�u�R`A8���]r�A�IF�A�>ȿ���g����"�Y�����Ynj��U1)������V��y��V8��(0BEF����Lx[m+�e,�[p)E��B���C�����	��#vK��:����7�9�!�z6�=��^ ��%'��R��,�����o���H8$�c������]ӭ�����-����S|�My��Z�Gw�9��Rټ�����C��Ů���^	���M�NEc�;�>�R���?��XŒ�Q�'�<�I�M�}���m?2�Ͱ�~A��ˆ�,^�%K~��Z:k�4��<F�.f�Z�d��$�F&a=A�*��?8+��q\�C����V��	���D:O:��ú�
�o�k�=��{�N�u�(��҉8��X;������5��,a��G�d��-B��(�w��O\ھ��6��D^w�5qbvÍ�Ӡ0�2�/���%U� ��x�!  �F�(O�B_��î�Ԭ{�5���.=��yD�a�lD>�Xo򥏃���6�LA;��g%�b(�m'�O�$�T������'m���^������:KT��S��������#=H2����+6K�g��$.&�����̖6ji�����G��y��hsG�$b��):��⫣�--��I�ۼۆS���.7$�*���m=Od�\ڰe���K�gf�LU)J�,�bu��ħ�k�A#�]\~�}y:iȖ���y�Y\QOǰc�wA�Fa��^�sF%�@����I�}*Z�oIZd�v�͎q6�Gfޚ:aZ�襗	_��٥}�b���C��N�C;�2m@5J�N��P� �߯�ы����e!�=��;��;��&�d��BS)��Kۊ��ۦ�!U}�)��_`���ܾ<q|��AGT�-�����uo��+Ny{5Noz���ͤ��Z~ld��$|_i@�h��Qv�4�r����X7�K�٥��E�(I�S;���%�xZS��R4?���[���D�R�C&J��Av��"��]¢�ì��Q�5�/W�B��w��JZ��z��̄(�v!X��2Eԥ�&�,$p�p�;�}4M�d!�_��e�M�6)��>�Ra������;�6�]�%�7��S8	1��0�Y����q-d��!� ��(r���0��L]�苨���4
���� �\$V��Z��`�p*G�'/���5�amH�&b#h����+Y[�W���q�78���\���K����J꿏��k[g�2��3$� �[O�Ԣ�՟*�'��KDl���]�wPS�l�]���P������S6,nR5K:s&Y��P�~2
vh�,Ev����[̀W���SڝlaX�A	ϟ�O�z,G�i��%I�1#��_MgX�C�~��W+mɷ͹,ӛQ�nk�lZ0��/��%Umt^�<&oXذ�l
C����T��G���f1xyzԥ�R�`��8Ǹ(7����հڭ�V3xH�)ѓ�A��tEM�����,? =i� �?�b`e#��Lp�%��q��'�ǋ�Rx��,����
f÷+�ui�����w�g�*/i5��9:�\��Т��_��
Rt�紦�d�M�R�$�n�W�OiF�r&���F內	a.�����p�C������3l&����'{zQY�qD�'�oO�seǋ{B�I2y�`��(KBia��f�X�~�Z�}�Ç���Y�,�@�E�>9�k�<`'s�1�� t��b#��m8�	��cr�CE�Ќ��q�<>x�e(Ǯ��W�nգ���(�?c��ﰳ@�>Wo�kת�-2����Y�g͏�@?W��=ɰ^�N3[Q���۴L��ds`NK��s)��A���,�E+�P��ܴū�Ge�������_i2�lyl/�U��\1TF譗�c?���<�����-�c�^�Tq�%D���hr~��R	����-#�K�-�W+p�\����/�(e����_)���&�_�Bp��IA��|�Y΍��w
�eBj�M^Y���o�5��F�{aj�]�C�) �j>��8Xy�`��k�{On��{���{�Oį�#=�V����lK�H[�*��2��H��E���7�=���|0�n���`!+BW~�[z�4�d���)����[ط�Y_Ľ��'f�����|%j]Ր�|�W)��F��\G�<'�	������Җ��!�@g�iy�� Y
)t�I�q���R;Y&~l=������-�QZ��s���1�D�*h��au����r��b9����x"��=�N·Ϸ��Q��˰�PK������@ �||F� -�n�z=�tX������(6+��֒�.�Ă«p�G��d�RG�$�|�DP|��&55U#:ܘ7 @��>R�����}��B��pf��`����Y��ƣ�<�j�0S��H����kqG��1�X�����Y[no�������s��}������{�(�d�8"�(Z����q��2w�q������1�2�����}C��x���`�4���C(�'��MK����� E v&�7��Ԫ w�B�ȸ*{r>6�N���ު*�i�.�ܾmS�]܊v���,�-%������_Ҁ���F�=q��y��ަ�w���,n�����]�
����PT�zKt1l�I8W���a��='#'e[����u���d��Pt���B:�.��m'��'��'��Vp���:�"V��f�qָH����;��p�S��R�0�.���\�]�?_G��=�k�b^�����R�
���[���y��faLǓa`M���YuW��@���,dU�f��w��,��Da���x�QUc�7��:�����u�sa�z��1�p'㌍��~W9��0��\V�(]`e��J�v��Z��������ܷ�89�t4ↇ
�,��W�|M�J��}�O��ę�{�@��j�Mg����-3@��w'-����m�����Vt2/"�`��}뺨엦S���(9�[�.�+&ō���y$#q�� B���k��I��,~WB��20� �(��#�I�^�u=�~6:�	�H� ��]T�dc7����GyA�e⮅���,;µ0�m��mD�8i�$�y�_ha$5�*��z刂#��%��;tx�L��<������/K���X�Ah�&�eEPrhdpe�
�V��T����s~8?R>ńϒ�����OOkc��ǐ��o�S���
dhm|t����?6G]؎(%��
�KyȒ��k�D�̋ 
f3��Ch�I��8�S���SIp�-%1��a��{���{�}uמI���,���*+������a��~wǛ��	�Y'B7I�Ќ��_l'���\B�<
��[@��bm��c+^�tf�6��Q
	�i���	�����U�)��Y���o�B�ޗ<6�ef�W���d.�1z#��2Y�5���E��ߪ®��Z�A�}j6D6ۉl �/d��0Us���o^F�F�zٿ�{q�D�~E�^KzFo�Ts�!r�+;�a9R����zjY��5�"�[L1�!��l�ɮ0"���!�ș$���]�2U����6,�d�5��{����{�??B�y�z����q�WP5�6��t#xyђ��VK�.���bB��]ʅbO]��D�C�|�].��')m��aGbĐ[w�̅�g=�
����+�m��)�V�wvE�1��������i5���ݖ1��ɬ�,���_�#����i7rQ�(����i�V�f�"�[��?Ac��0�O��v����	��<��2-	�e\��>1���$�,�j��b2�aQ1��O}~����h�ו�,��JA��B��a����t�lu�=U���}QfȮ�{��B����45��Q�s%�o~{o)�4((�g��Ӽ��yx�zUb匎��6_zx�����ěqb�z���%��>ЮR#�O���.+��w�i}P�[QB�Thߗ��?Ѵ��*��6r�5��~[=�{nl�\��.�C���|k	�~��o*/����4��D��=Agfp�/)�Sؿ*�'�t�H�#�z@全���G�G�r@�|�7ު�0-�"�|y꺀�	��p܎�ʋ��.���'�_��3��",X���0�x����A�9��v��K�goK��0B	���t�Vt�3=
L�ˇ����P2)���5���O���f���#�g���̨�x�8�L��.��^���W�:L�^�Q���1�+N:f����le��*��E�b��#���i�[(�p�Ա�&���"������*�]t\�F��m�.u����cf�
҉bi�^WA<�:8p{��~ yt�ܼ�m�"ap ,4��
�6���$$=��0�q��R��*�\s#����t���͢:A#'��h���e�h8}S��8ѵ�����W���/<�:ן�b[��=�O3�o�i	��,�:��7ʭwիvu�YӰ�Kè�s�Q�}����$�����{�mQ8Z0�~[<�����
�NXC��4��PfY�O$T�1��S�!�L����e���I��e:���ۑ
��&[�F�LU���Cy��d-])y��7�����`��^V.-�y�g�����{�(PDVZ�O��;&~��)Id~^=���8'�:-4����A�̙tQ��j�v�*�t��[�P+3���=�@�l:
6[�P����GpN/Zs���\ �`\{e×M�[��n���R�rw�Zt�"��[�ԃ(�f.Z�$0�|��_�.4�s{�#ɚ�;>�Ӯ���z��>�#đo
����r���� �z>A����Is�o��3_	y5G�����~*O�o����e���N/�p�BK�E���@Ȭ��Ta@�H6W�{d�d.~!{Ed��Xb�ْ��v�C���=,إL49�e���$�TCo�*��z��ԷE�>y��1��/���e��0vJ�1���0����j��{���@��
�hN��yB��h6����Е�N����lߣ�����Їiɘ��0��_n�D�7Bڂ�`r-�P�Zߞ���`�MzjA������"O�Y$Vn+7�֯$~o����5vsB� �+��4�#���ǓkmL����E��^o܎CJZ�vY.r�����, ��=���	�.u;~����Y���vf����^Q�H��"�+4t� J8�u��ߎ[O�]�A�UFV�u� 
���F�'�����>X�X�SD���+��#���`h
$>�*�>_)s�"+�rvq�!�lz����#����yMD֫M�١�W	�/��`�A��߸�{��I��5YJ1ļ�nK����8'{ {��m��T��n�7Y��m��z���Qb�3��ȻZw���u�vŬ�~G�{y�s�yp���B�7Q^��d�uըh��PM�k����v���ܨΣ@u���N�sOE� L9�ϫ%.�>ɋ���>��-6k�fl�"��q�&�6�1WJ�Dj���Rz�Ƽ�>Q�8�C�튛p�>�O<=�Gf
�ݳ������J,�P��mᤲM!����T������g ��s��%���o��T�1�+�;h���rs�@>:���E{R�rf=��!�W�l����^I�Q5h[@l����fؠ�I,ӌ'0t/퍮���Z�e��nmPiZ��p�l����ȣ�J��S���j�Q�����cP���gǝY��T5k�u%���ɜ
^	���*[�\���=�s0u����1����=�j��L{$/wʽ-%L��K�7^x�F��ݽA��F^������xuA��]�޽a�T���`�-�
�'�=�>�l�-��h|���$Vڀ������7�5���e��2�o��q� G9�u�k���[q�O�j_H��H���RlU�L79	����?�,*^f����7_�㒐ph����C�{��]I�%V�0pE�Z��!G�}�D!ޑG�"k Z9g�? ���`4�ܴ-���6�B���m''�<�����4��U�qg�!��&}h���VÊ��j��W�*z�Et
Z��� Ͼ���h�vlb�r������ʻ�C�X�x4�ض0-{>�1U	1�T�F/:�[xV��m4���l�M�w��)�*�H���;��k�4��J<�6�j���(�ߒ�B����]��S�E�	�;��趘�䬙m.o=\1V��A��O2�����ˢ�1� �Ks�"c8�!��}���[��"��-qN�FW��[�3�� %S�^�*�j��B��x5 4w���7�u�3Wd�1���:�^vOm۹�e���`�HI#"<H8i����.���슍
?:G�J[�w$8;Q�x�;��Ւ�����_�P�JS)�GeY�@|$]�p��tvx��g��*W��{���J�s����z&��4 �;����`w�uzG�@��Q�-��ܘ����7��g�C���p���U���b?���I���v9�&�
%��;]G�pa�#��[�/;�� �N�j��J}9H>T
H�B��?�Zڏ�`l�0���\"�6B<kIValvCh�fs�z�B}2�$�(x:��Lb�v����W-Ț0O͘F"�5C�yFԭ�����"�7:mIK�B{/�]&�"������{�*��>���c<��eC�4��m��+[�T���"/S��\�W�I�jjk��=�I��9�4���BE��`���"�x������M���Zy���
����(���k�&[������O�[�jV;�jR� 6)lS�/k��U���r�&ދ�L3{�"=u�[(7�W7Z:�CI\��J(��,�?��������p�H4�!�/eV��9i��c�(������
�?LT����=��wZ�u'h'c�#����G;9~���!1�-� htϩ����f�?F��m���K�ﱜ�#F����j�i�&����O7{�����C��#�b��J�k0$�^���۶�=s���9a1�tp��s;��U�F$���]<��ɵҕ6���O˺�� 4��-[�z��ī͍�N t�Y+�o��I.�!%Ho���!�ޞ9�L����� �Z��9��-��ಃ]���A���~{o@�{��nxNX�Et�+[�7��N��ثpGm�يA�22�TZ�,H���!�4��
�T�h���B��&"E(�؏����"��(�OUc���w���E?	�?�̱�=$��v�S����ml�5���d�����#z"q�^�P .�z�g���Naw_�r,Us,$'hx����M]HWاW�E=`��wa�z�M��Zj���.�M���YzLݒ�����[�+�w{��� mn�\�c��vV���'�D>=��eʗq���N�v�7�{ch��R}&Q*�N� ���q�ƙ�)��Ձ�T]�����Y����/����N�6��������u��������7V��n�C�,�DU��9x���X�X0��r�G
��lA��|���y��u�����\6嵕�_K���k�Tu�te���l��2�YE�tpg��c�~ſ���uo@[#�8X����~��1����[2�7�?�&N�L�Uw��A8���X(ǞBF �J��@�<k��f�5��5���q/�j�:��WF��#�_/u$�[L��+�E
��}�]���8���Ad�9j
��p2���i�b����b_��Q���ӧ7�ys�Q��[���m�%�P2�3�g:x�c��6��@!��+��_or�~�"l�?�Q` ���@�hd��AR�|j�cl���OCc�A�y�q�&Gm����TZ��˲j;݉nЕ�����&��y��s�u��wA�����^̋Qk�y��k�~�v�=�C��#8)w�>�#7����_>�aU�(�ϋ)G�uf0�ʙp�;�f���Jl�jͿ��Hba4lp��:P l�u~ǘʨ���u�yʥ�)�^WR4֮TB(\U/�
 ��Ôb��F�|���P4��H���^���h��?�n��g?C�M�q��D �v�ttOG�䗈�	~����UQ,�NiҼ�5vӹ^�;��/*�i���˝�9�NUD�M�N���ݗ�d���@�O)�M��mk����h�c<S�����֐!x}�(#'?��7��R��S��%���A����'�j��1�P����%�I�ݙ�g�"�WF���U�N5��n(�n~���g�Z�O�m�ѭ���BZ]�:�~R��K��7L.mNg1����2ן|��{�dT�ï�P��#��}
Ф(F�m�.X�oH�q��Qʂ�yuo16���W��EY��e�N��VN�kL	mJ<��Z�'e����v��e@