��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������-��
1����yr1FUb��q�ej�IϢE^U�nA��a��"��� �AMF'�k-���޷n;m�o�}Z?��$Ĕ��L�h������g�Y]�)�}�"��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�?2zֺ�i�UCv�~��t_.> �KX�d��@�����O�2H�%��
����)�j�6�Q�؇0��E��:��r�;xՐ�>��~U�Љ��ӎ/s{p�|2}���/�&u��y�4�蕵���b��\���ի߿����{��(%�X���`���0�B�͎&	�3��������x��q�2�����-6����5)�:��Jt���a ���D˄*��V]u3��	$�RYu�������Os�Y�7��v��n3~HGC��,��,����A�����e�Y�'̲&�Dv뿽�3
[!V_�2!�#US��_3�i}��<�[�㤪Z�g(�@͊�y�=��Ie��2gV3���N�	J2�?�����EX���Sz�\%R�a�(	�Gy�j<S��˖.��� x|�I[bi�@���ȳ�"Z���{�� ��d䫥C���g;>����7/ ��_q0�:����YP�Z�l�������) �څ�B��Q:�j�Յ��K�Z��� %�C�.٭M&<³�Ag��ի�_9vUdfA�(�~{���{O��/�ĥrv�������톲���k�Y�W"H�p:�J���A��,8�dy�[:������7�O�jy�S���9�l����&;��'�iI@l �]�4,�aK�ٶc�3Z\�؟v�����Nk/��y.`�\3�I��8dڢ�c�j�@y��otΪ۝'w���~_�qb�P��P�,��w�ɷ����)/�t ���9b"5��g��RSH�<qPA����ru�Ĳ��ʹے��j�M�vo�鄃D�l�e������y�;�U4����3�Ӵ_���n��V�2n��j�r��{6�?��'Ĭ����6��|A��|Α
� 5�*�검4��Rk��B`��)ȅ,��d"�6�
���<��x�3��m@��q����?8"u���|%4Q��0�ؾHތ/��wZۯ�_\��������#�"�]Ĺ�ط��U6�e�#a�;���GJ�g-ࠬ�á�������
T����l�%����v���6cBi_Xܪ�En#�)��4��]T�2R|�G��cƆ�ߢ��Ԍol�y=:���Kۅ���}�8�U
�����d�N�M�Mn):��*[8-�[���xyἓ{�� *8�|9�%��$��V��&9��	��j�Uf���ZWI�&!�vإY�����s��{Q*Y��Yf�+Iڗ]
^<��}������!ޥ2�T��|}4�@���d�;������N�g�U-��E���O��h=��h�J���P�1poi;��#�X�/lG���0Qh���GH*���:����V�c5,�������
4��)r�ViNza���$��W`�Q���|��Jp������/븶W�tLxd�έ<��z��/�ݞ8�(I�Q�?��m׎)���$.��L}8Z	~5����asm��驑c�*d��A�g��[L�/�����2�t���9�A�.�WE�=��#�&�Y���Оڀ���������$�_q��}����3d
h�uu�(��cޮ����ʼ�
�Oc/I�@����.��Ҩ,�E̋��V��Y*š)t���٘�3���鑙�����~�Ul7�۬ �z*�\��`ֿ=]���w��3���&�=����W��P�^�޺6�� �~���nhW@�.��G�l����������@����j*��'��"��W��*_��A�A�a+D8�0����p�v&���F��
n�8����&1(���4�k�F��`x��{���>M�5�C�g�X2WGN5Q]�������0�g�����Br=a�սʧ�-��"L=>#Q�5퉎w|��h����Z��7Ϫ�ˉ��Sųj�GW�z9OȌzE�AG��˕p	>�N5�V1�/g�dة�5V��v4��^Q˕���gV��� �p�3�5Y��������4$��G��w�9���`P�%�;X�[��q�^�K�2�pǜơ�J����"�r�Ӓ	��Ԣ�=�xM�����}`8Ɖ�!�S�/@�W�a�_�)Պ�?��� ������Ӓ	���a�&E�w�r�:�L ��P{�r�ʝ	�HEˏU�q�s�{�(h��9^B�n.a�-@��������3�h��������Փl�ΩO�s�|ۋ�����\�[v^��s�uc=
9dxc�B=����i� yq^���IH�95���##[���B?Ž�~c�2����X�a�w��̑C-�gΊucMv��	�,���Ju�f�	�W|7�$�,s�GW0�.�?��`����f�c<�0H}j��?�r�|3�ݗ?L�b�����š`�F��Jq��X�^����̓�Y�[*�!�d����������d�7�ie��cfZ�0���h�w`��{�|�~o�H��m&"���o��UCB�|���7���4Ɋ+�)1;�GQ �]��U�T2|{���eڦa��+��[L��G��Ef�o����cE���ԧ\U_ɦj�pf��?� �"6T���fI���8�𦻎_�3�IY �=�Ri�C�%4]#��� O��PX	:, ��SIp��SВM6(* MJf�a�Ԭعk�\Գf�����@OKd#�C��+�n���J����_��F�@����
���k�޹g�;�m��9����a� � %��:��j������o�a�4D7�oI����ޤ&)O�!�A�U�� ��ݖ��cH�mz��e
t<A�A�>��m]@\�+

?s]Sm^r�j���ri�����4_ �S��+x�����+�Ƕ&�.>�W���$}��`s2U�i�m^�$x �l)?ÇV6+"@�.W.�oF�B���_7��˾n;�)�yZ�Q�u�&쳴�r�
>�|L.�N�#��V�����Ÿ��*F;f|G�/sd��E�kK���b�.,ݨ������n���,�e+w��V���]��NQ ���N.����P�� ����9��\O�	f���s��:|�}�Q�wj���%��/"vA���ri��%�@�]��dHe�q�����+PN\���?Mi���zNڸ�7{��s�n�~T\�AZ�x��<��7ɀ�R9���%n(Q�ba�&��y�x�G=�\"�탵҃��*���plJ�z�gw��Ƹ"�����(���+�h��:��I|�#�<��r�`#���*z�y�SwQI����p���Z�`�L����kum[������#�r��ZY DxQ�<"����U"H��H�5:�:�c�:�oՃ��؆�a<�����L�0��É��eF��,n�9�|�g8q���� ���#s���jH��H!�"�3~s��
W'�|�v��O<��u
��� ]���?oB�is�����P�M¿������1�؝��aڢ��RïI~���cy��^ޅc�p��=f���@lӆË[�]W����VifV#���F�B�v$�49��Y��Fzǝ�%$����XL �[����Y�1�~�E{+����T80
�`��/�B��z��΄��P�^��w�-��OeN�4��k�a %������_Ջ�C�Fr��l������ ���ܹ͵��+)�4	
K��lX�\+����&9�x	�Ӳ��7�-�.��+��n���:�?c����̛Bb4�v�{J]C�.t ��HX�.��5��,��6{._Ash�K$H��no�=`��U�4Kđ�#��Y<c�]��׽i�&�=��Fw����F�L����Z�m�{�l�e|Ȼ�-gQ�Z,ÿ�l�����#�I��{� '�=�ac�"�����;o�w ��\�o��ˡLl7B)V�ry����<�B?d����#�`�a�@�!��A��Ѳ���aGx����E�-x.������V����A{G�ʢ���t���_|�![�`{.��$b%���o]���&r�S�xJK�9�+Z>������+�#��@��^\ۀ"�k�@�����S==D���i �͹j���&vJ>u�0��33��|��?�0���j�7>�������k��Q8H����X�oy��Vԏ��M�qj�T$}ۏ��Q_d9'B�+�y�E���^?Wq]���Nms:��\h����z���!���fMݬ0�
Z�k�heV�Gl �⳶zb���<L��2�K$#�~0������_H.5���'m�j��i��9���U͕bj�������x�~��lW�����9Q���u�����Ă;Ա�r����9��#�*}7,���hm���.�1=>���2��x���T��f����&�6 d��H�F�_U�D=��:5���W�#c���C�Wd�*7PwE�m�c��l"> �'�b��/�E�u�R�Zg�@����<ƛ+�����U�҂�z~�@<�Ϛ�����B�?q���'�e�S�"7w�x1"�>���������˿7��=y3�4�G���RG��a6�;V�~ת�Ic��f�y�ۥ(��C"�A�¸b���_�NI~fߵӝ�|3#|>�A�X���;Ҹ�s����.l������H��%H����pS���=0f�b'�d<��-�BxG����4�4�t�G%���q��T�R��<k��/�+�%9}�����3�[�I����=������ؿ�|�l�9Ϲ�y��?�Ե���̼������S##la�Y�fic����^��y��k��4/��3�0y�!2���[p��m!so%�i��(�cqLs1�P����}�O-=A�(�B��"�ܽ������W�����֧�s`?��ɻ�`Z/�]2x�� ��9�p;� ���˰*���.U��
;:di���t>���1�>i&M��=�@�_/^��2;��;�~�l��F��/X�6G��Xq���}�p�SPkk�.����-oY��]��J�-��~�0�5L�ʩ�5�j�8?��gc���Ӂ$�	��t��
��=E�L� �ռ�p'���������/�^C9��S�������q	���q�|����C��p�=X�	�\�=���&��������C,6��}��E�q�Q	�A����U�\g��k�E��k�|c<�������_���Y����ྣ�����0 ��+}<�>���dH{�~R�M�5ß��KĽĹ�-o�4(h�C�C��n��<���JV6r� V�Z��<F�Rժ�%0!���ׁX�������(�ZN̥<��&�����H6ü�wJ�2��n����ǿ�=��?����rQS2�J�����ѷ@e�^N<"Πp��n���V�1�)�k6��R*�M�Exuno�n�^ڲG�(�Y��c���͛����2�_)q���jk��$�� �_�;��8,Nm��]�oC�
��[�����0ӵ$�����������2�W_y>-��?�T�����+�9m�.�ܸ���Z����9�'��c�� �m{$	3kZ��W%�s�2Q���L�Y�\�iB��u����B��׈y��^Q���f�B���8	|���`��36&�2�	9�
i�x�Ⱦ[|����Ιw�`����u�݋Pj�3���p9��[+�Y�m�K�x̺q�Ǐ	kL}QÃAq��n&���/��M���gI���oN�dp�{5:,[
��Pi�W$zu�*i˴��e�e�Dך��+�l�˅K����O�~�2E������;7tC&�>�OB�Ñ#��K)ew���9���/�Ȼ~��� �����(́�F_�grc���jN��s_]��Kͮe�ue��<�"�%�l�fV�v�:O���Qg�~z=H2�Fm' ��`2��o�d�aD�OG�1ׄ�k��K�Wm�N��"��9M������OF7��NȒ`��h�= �z�Lh�d���e��
�5<���F~�By�p�^���Ç�\*>A�:zkSXf@�S~2L"�� ��ܴ�^}�1��6���y$�s6��f��%K$�8�%����n����O������r����@���m9�ꂩ��Q�{�q�f�6�G</r��Շon�`�2���W�p��+�t���v����V�0��ԥ[���Ѓ_��-�]~9P�t�y6Xh����0���s��W�
ަ@||�=�IyO`l��K3,�f�3�f&y�I�*P�3�1O�a��(�J���Sf�ڍ w��4�R[�߹ ��j���������=�M4T�T��U"��e�?�?uܗ�k��U�{�!yj��6�m����{��n��7f����u[:ld^�eq-���P�A{�3t�lC�ܼ�s9��Ӱ��[��i �O�j��FW!'�4��h�J�e�[���(ۯ<s���4�0joL=��Gg��c��J��ק/O�Y�H��OЌ%�*���7�6�S<�.q��;:u���
�hӋ���5t�Y�h4���v���⽜HQ�K��c�y�{w�\F��m�q.U���v�j��W�)_u!P�_���B9q��s:�U��egMy�|��K

'����nb�ߓZt}�ܡ�y�q������z��[���׻c�{�0Yo�u���~��U/ם0��W�ELt� fE���n.��jM`�Հ����r˜��v�38��~�5�{��\��$��k�/�'r7���Z/kL����H�	�H!e$���XR\�\<ݘ�ެf��� �;+NƖ?��1�
�u%W_.o�V6<��id;��Z�_�l���A޿�L)�oF���BLF#o�k��f�s����f29!�"�EJ����F-w3��m���5w@[{\7%.��٪C�]aer9ٟ�E �o�`uU�:����l\�υI�ky��=�^��pV�&���r�l���m*ޠ65�Q����4O6���y܏{WǬ�}��{���m�qy�vR&5��=6e�V~.�c:�'��U�ڬg�C`�)�TL9#������Yn��pZK��9���O^;���⋾|�S�.���va����-�XO�NU7?t�MYQ��9�W�s�YC���*��=o�m����7�l#�2}�����&C��؆�κڍ2��a��OLXg�~ѽ���y���L���f$^l��C���K���H`v�Gz�J��;��� ��ӔT��ԭ���p�o�fj'0�q6���L4d��!��$�e�_s��9�4f�Q(����U$�mQ6?ێf�<l<��s�"�L��|,� �u4Ư� �I�}uOC�2�#�`yc|IVĥN�M��Ή�3*�(>#P�RK��*�Q�%{ҹ�6_㛲��Te�
�=�	C�����]�ϻ�v� 7�l�'U�2x�xR;���s�s�9���$Ͱ[L��r=���� 4�����P�
 ����b����,=�XSb5_����M��ְ�%)�mW���\�!�k��l1�qC"�I�ct�L�R�[ճ��o�ihɼq��.(δ0�Wv�,Q�+��IP}���V*˹"��ۇ��<v���]7��pۢ"H���ˏ#��D?�s`I	�{�Y�����|�aj $k9Ʃ�ll�w� F�D�~_�b��H�;�m�	�)ܺd:c�c�[��R�r+F����r�#�|:��	�^S$�#X0���qbUx9��kbg���ұh����
��<���A\����*i;�˰n_�7%�.�3~�(�C��Г)-FY���e�����\Y�����LD!�MA�Z�ckt }1kK�fm�c�:x��t��.���~�I����A��p߽{�N����>d���4x�����bт>��]69ڬ��ߞ�^�Mן�ɜ�:���dv�*o@s���P������9���]�ȃ�媑�3�x@׊�?��5�-T@^��ݫ�i�?�UN���c{����?�H�C�;&$� $՛T��c׭Iqa�̓�Z.>�pz�%�{��JC�t��ҏ�U4��$� M9�c�OQv�kˎ��z���]T�@���O��}����D������)�*���@��|{�*"�s7mf�� 񊍷ط��C[��ڞ.���>i0�i���#F�]�y)���cw	ŠG�A3pj���Z��ŻG���7�w������@#��Z���\Ҩ&��DVU�S��XS���g�*_Ze����x�^hi��&�h$2ty��!���B���9b��M����LI^[h��~Θ+�o���[�jk�3��>�ӅT�� ��&��,p����.fw"�Z����]�-���,$�or��sž��Dl. �{'�5E��)�H!��]��ibz�� 	#�������J���#��ߩK!$�|���q�.8n��l{$Sl�a���f/���׌��r?D�[1<qs]��ﭬ�z����'m?�~@�C:�_����V���}/}>�_q+x'	��JtI�Y���\*�N�@��mMAyد�}Vcm�r_;6���̺;�����l�=�ם����	C4 �g�	��K�y\���x������G�B���2)hE��:;����|O&%��{b�����XD0�>4b>����s���756��� [hsP�Y����,4'��g��2�����3 +K��=�C���e�?O$�.y_L�d�<����^}e(�v~�X�dv�Y�7��9�M��
���p�������t�]bP-?R?7D �TB�8@�<�c<$K��v̊��(�W�]m���I��!�j���4���)���X���#����j���T����PF����K��k�(Kw߉l_G��e�� U2���l�g�>����e�X���=!u��#�~�=	���ǾZ,-`��ؤ4���R/���[�5�$��Ӟ#k�zd*hF2�A+o�qk�Y���'�E��G�}h����W��A?��|l74����a�\U9��x]�M%
����L)�P.�Kz7�I���_����W��Ҩ�=1%����'-ŭ�1ĭ-;tu�]xS����l�B�%�<�=<�p��#臲[<����b�t(>��g[xj�9��a�^�J�Ae)�;l���Fp�AJ[�R��a�?�c5t���rǈ�[�	�~J[󸪘;��"������bq�	]	w9�c�,��>ͺ	"�+<������D��b�I�ga���V=�����^�8�;�-�[.�e��s�#fI���G���%���4�d�Y������׌�dsD���l�7�lVG4f����?���t?us⾜/3�e��U���75c�t�L�!G�#�[�f��9��8��� ��+���n�����SĲqq�稏���m W}/�TJ�D� BD�0��9�׎	�kN�5�����Շ��-���P}-�b��j�6��U�[�x1�xzą�д�u0C�P��
 �P�?C���{�sq�%Ó��ݿ,�k^�A��P? 7����4�?�}����y����[��k���ڶ�_I�l�u�����Ϊ)�޺����[�P�ߘ��?�[y .d�� ��i
�4Bk3!а.�Y�itd6�<d#<�����'��f ��Ǚ�	a<�޵�֮�z��X.@�(W����"`�e�����~�n}���T����Kh�p&̩u�aE���(��m I.��:@�橲����'���0O�h�.��$�����a��O[O��!3?�>2�b�\���'�
>��t�5�<�0���O�`��"j����
3��:�O���^6�W 񆷩K���?q/y> �h�ý&�̤�ͱb�Dr�Ps��_���n�i����rUm�*� q��
�^���X�Ƣ�(���;�I�®c��rBK'
��O)�+�x3s:�丬n�keGa�V��j&�+Zo8�d���@	Ա���%w�0M�SUm��?I�B�X�x��@`w�^�(��;T�_9���,|�8��7=T&frg2<UmN��':N�QPD��L���J^������%�i�_Z���qD;�)|��������K��1�i��(�d�!��V�d�/��H�\XG�$-`Wd�V��i~u^�T��`L���i��j��9�ͰmRob$�5�ne6�Zt��2�]u �|?��K���kJ�Ш-G�)/���#fʌY�E!�$�`�4H݋��ۆf{�	茏�a�$��'��P���p��R;����%	���7���O��ʴ#1g#��0��nR1]�n�+-fw��0_�w�#�a�;��(H�*0�O�,�S-�4�駱@�Cp�`�B)
�6Rئ�;B�|&A����G�LD\4IP1 ��;�\L��!!����FD��DϢ4R4��;�e���. ��Z?��=n�i����qaa�������癅�Q<��%Zi�H���l��-�k�M��"���u�W���OG���94���U�C�,�u2D'��w@�֌��J\�E�Xo\(��1n����<��EHΆ<�3u��vC�iS��_���w}��(�K�X�������n���c_�X��9}���<\a��dl� �FJ��d�Y.� ©Ӕ�7�#c}����}�Z����8iR>r�>8GS�j��gC�۰�!�ABs��3���ɴ����vav�q�9��u�A�폰�ږ,`'}.�]	���mS?����.�ĥi���"�17a�M���#ǅKI>S�U���LpN���ܳ��#�Ɂ@�鱘�&!�XE�,-7��<��*��ٍ�ht%��KH%�x�� P�i%@���{������{�cj{D���^W;�*��D���Ì	n�8���+3YϠ;��.���9q�-U �J��zoU�jO�!��z���E#�s�@�Vd>�������wzG�A@���4�Q��#�4���J��N�5��O�b�����=��°I��.	bE����q�ף�^p�y�)BA������z�XO�e�"9g���+R� ��a>��Z�ݿT<�5��Xeb-���⁶��*i��X|~�r�U5��@b��l�� ���.s�~��9e[����Hs� �I�P�$�J��S��ʵ�	k��P;�]�����<Q������`�S�.�c�Cμ�L�jGè:�� �#$�:o��KFst������/=wr�,�_���ݲ0oBŧ
��ϷJ�@k�����A~���q�=�o�Ia�5���Yt��N�%@��B���F!t���]��!��1VyӇ�P��9����JA8m$h���Ǟ��N�N5��|�ͫ��X��v��`Ԛ���揖����Ϫ��������������'QL�@�X����9CxZ;�����l����H#*�o]i�1�����r�J�������]%�߳;�ˠ��P���E����u��7" ,w2/�6�Lx2h�|7����2ɴv��4�