��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������-��
1����yr1FUb��q�ej�IϢE^U�nA��a��"��� �AMF'�k-���޷n;m�o�}Z?��$Ĕ��L�h������g�Y]�)�}�"��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��ʺ�5o�1��Uh�n�}�.��80@b��bb>�WD71��.�4U��|��=�kvߤw5��� �S��Ћ�EB�ޡ0 �<��rV�҃��Uc�vƷ(~�h�y��O�f���@؜Pa��,���� K[B�	��YR�Q��Zbz ��;i!�K��d~;�N� }��qZ���J�g�U�4>���`�O����� ����F�'�[Wי9��I� �٭�Y1�ޭ�!Sb�zn�2 �ޘu�{�ͺ�I90���>��(�>��P�A�i���
���U=U�#U��2��{U����n֑�+Zt��a|h�����a�{O�A1�&>IAkg����d8���'��ac��ڤ{D��7�#x�fZ�x5���Ax"�}�..��cT�H0U��\�m����v��3l��,]�vA��Z�M�w�Y��o���Vn�b1��r^�M��0�9ƴɷ�_LԹ|H{�N&*v�C�S�INf;�7a��	��{���]��I��\2<�����'�����.M�Gw>w��$����I���G���UmB�J��Ȭs{�h�¯��I�@زs'�]/���
�#G��q�k�>�)ց&��vI�4�
��S���Y���$��Vų�4��v}��߁����j
��5O ��w��d����ӃnB�9;���v%M2��&��k7o�"�U����V�\��H��r5�����P��\)��IJ�cD%��I"q/���q�Las/04s���	��8:��G*��
]�Vh�[eڷ�U�L>=��)�r�����s�+�bH&��:�7�^M�������$�M��kl0�޸<�CR�١�O&�:�EWl�w��!=����PO����Ϻ�?y*��[�N)P��J�î����B؋��3ɓ"�Y�>�!L[]�~&g�����h2-�\��r|�m��������0t"��l��#�}V���K\��	�uG_��2�Cy~S��Q:�(��Cc�%����a�c�E����i�V�hh��* 6-5���ׇ��-6Z���|������J �[(��>�Ag�9�6XL�<W&{?�=ƙq��=�������$>��)\�Q~�Ik�=y܁C� �%���#m�oQp��3��!�<* �.��=���}�V����*iu	�����Ũ8F+V��Ҷ�J!M�����[��<_�y?��C*<�f����Zf5\��]?r���{�j?�8U�C��]�W�0<l�	�ݱ��[���:�U�$,�y��yp[�ѩ-9�=V�L����7q�)����nP�mBX�\��eݸ�˗���oe��� ?�\�͔u��S'���
	>��E�`�;�磎����W��߱POM#d���I`�BǙ��kR��G�ޘKB�,�q�d\��f�P��ޡˋE ��r7&uC��~4ww y1��}�{`��2�����z�q���%1U�A��MP̡ia���.٢�7'��6�~j�:T��X��������2������g��[~��9J�q�X`�1�/�c]	�s�l&�}Ou���R�$�3�n��9yl/�*�X>���_��݈�O퀉�����ڞ�K�m|�!҈b�z N6�x�.���Me%x�%231�F����v+�O��e��-�U�8^�:
q�8�+�4���l�U~m�mbڟy �s�#�z���jGϥ�IV7��T�!�Z`�E|@ Ix�ꢂ�/>��DӜuBz@��{P��r�ڿ3d$<Յ��Y)(N������ǆ�q,� �o�/�r������kٺ�|��.$R�/L2S��m��)��i`�`?wϭM���n��o����E����f�eҰ-.D�֖:���di!#�Z��H�y�C�a����h��Ю��d8��s��P���tib�'��)�k�vHQ�6��||�H�[xZ}Ν�o2�ISw�p>V?�#�&��I���<�S�q
M�c�0B���-����c�ٔ�𶋉�oވ<��}{i�b%�����Gs@H>d�V�= �FL�r����S)(@��	�I���Ň�I�1N��H[eKU4SiX6��f�� NȾى�S�"�j�({���{_��]?V���Vs�#,�}w4"7�Ue���,�D����oS��g��.�. +c-�=ʕ��o��c4��m�B�Y�gR}�
��)hS���u#)Q,@$�,0Bj`�z�ϛ�kh����a�l�,����ӎSAF~�;r��L�FUP�9Q�4�v^�nonD/��l��qF�P_g�DY��|3�r�o�͏Ѱ*$C�0钿��������f�Ԁ_��>�=Gt߁:Ooe�n@���)JV?��g��F�fJ�K��z�e�JA8Ts���t��I\���m-J��v�N*�S�c��J��3��yC��\m^ic9l���e߉W i}LY"�߽�1���l�k�.����:�e��|��#�? �2�N��8���ݱ��˔W��'n:������46�?��;l�ה�Yr�'"-Em$��o�����r*���cܣ��RP�TupL�~�x��/]$��F͢�����`�v�;�~��~D��2@��[w��ު�r|�nsqB� o���A\�מ�<�Y�Н)�k	��<��LT����?)�X��]�.�R�&��F$m+$�_/O NRul���V�ַ�!X��!+E�c�:��;4��j����XG֡f��@�U�Ȯ����=�8�P+s#�$��8��R�8�n��e�EQM�	����ՐVAp�ԫ�j;�\�U��sXm������+�@ʕU���6md��|10��>44w�cv�C�O�f��
�x�+��U��Z����H6'ؿ~ۍ8�QMK�
 �^�'��s0�ͨ�n-��):���
�d���J������m5�_p:��$ Y6�gs��@�8 �ԊD�z��(W���i�εp��U.��SkӖ+a�x;�c�1��l�3A���6q�JJ�wЋ QX#�4F: �c�"�W]t��~��y����hF";��dE���$h~��uw��y��㤘s���,�AVMǯ���$���:2r���ɕ�,�%��;P$��[��!@R�X7�l����F!��=�c-?���Ǔ�!#+k�^�~�?��O�D�D�X�gw�d�ݸ\�����
�Դ�f5geEmn��9��D��>%�,_���Sٵ ��J[�<G&�p(A��Ϳp�� /n9�������.��'<�?9>�xx���|���H�P	b7����
��-��-gT�$ؐF�|+��?�,����+�Tr0���a�.\kyʌz��ѻ�t�+JgJ����/������Y6S݀�B��Q�y�������^��ZG�r���=�;2ZS�&���u3;�6�goJ��Y"�|E&���u�d��zK2�$��a�����k�,Ǝ���#0M��"2����'k����hA�C�Y��	M��ȁ�J�ؕ3�X�-+��w3�b�;�ó����Y]�n��h�X���@�E)ϩ{��@�Z!���V2�c{D����ַ	s5"��г���m��c�|?���({��C�I㑿:vN-�B��f�#&�g���)b�o��$�Z�iq�-�|��Hx���l��+��������&{=�ha�,K5��Ok?���e6䲣�Y�� j)O��h�ʞ�3Nj��o��ɒ~��<�>� `��	�T��B /���{,7�~�K:qh�t���}I����oаΘq�&y�����N�\����r�)�#���"�	���/'��c+RH4\Jr��3�Q���8�?�5�I(P�D��Q PPU�xa���%�40�5+'4X���խ=Z�+5ϙ��N�f|z�F�a�I���캷i�ƅ���ei"�i�T�\jDTO�{<�~=�7�� T:<�-
a�o&��x�U���瓀[+�X�$"p�煥$�y�Hڍ�=�M�#��j�Ep(ʻ������3�m~w��������&�׆.kl�����{�6����[���t�1o���k5�m����_Ɨ	g3��<�En""��J���E���U�>0��y���2φ5���7b5υ�O#0��{��=\���&������
����:9��W��V/�v8|�p��������\�J��+��6�K����o������� ;|�EJA0�<dU^����fD<�Z��φ�Q�\�1���L�]��w�H3�di���*]���&ú�}�����)�p7�����vTz��?ɯ�	7Ȭ���\�ö�Zus�Qfbx�d0�?���|�������T�\EB#���Og�ǍX�$��ɰ�YG��|+q�}YM��Z˨'��.��!�K��X�#�p-�R-��K$^��@d.���y�	�&rnR�6a��v�'�@�}�%��%Q�9�mr�����λ��������x�I�(q20��2g����j�:0��n��s�9J��ʉKTx!�IL��B#��g����b�:7mQي�J��蘼��̈r-@�]��H�Ok�:Nx��Z*��K��)��� ����zNh ��M��b���0*���$��İf�� ���s��3]o��������{B����g..B B"bA�ٿ4%����o Cs5��z�a6P�L!o��Fzeq�Ge�x�π�s���G�X�q���WK:F��5�g��7�h��rх��.����|��&�Fކ8����5�E�[��VPzD���F>po37����� �|#��J��#��m@y)o��P79�� ���C�?��|>-N�Ys���G�	zY���[���!�.-	�W�Ȯa
y���|?>��ヴ+�4�o�����f��e7��o���>J�#��5�lc�� G��8�SL�n����k5/��9�����׏���2�|��b���� Jἰ�Zz��=ɣ��BK }!�2N�q�DL��|���	��{Z��?M%ϓ9ǋ�������ia�]���c�i[�� �9�l9.��mMc��^��汫_����()�S��{����⼩·�G�U�T�os0]��fn�^�I��<�W��b��������9�V����
C�W<3�9r��Y�����K	��">��T!�s���n��VmSs��g(o{�n"�W�t�萖������2��z�t��-{ٷ���I�I���ޢJ����2��� �NC~ܧR���
����Q�n��H�>?�E쫁Z ���G�v@��#G5�ھ��/Q{����bڵke���&�/9��S|<�ٴ�b����m�q_�@��TPC�(�j|��""��?�S���z�~�_iҡ	���L/H'�!���Cʌ�;ysi�Q�gY�Bh�～�v�0&��*A,�e��`˧劾����g^Zh1�l>�6�k|\��v��IIU@g�=���F�J��I��H�>��ׂ�z����D��^�4 �䒦�_e]f%�\� �A�a>�t�;���^Xr/��}i���[�]:{I
|jJg۳@��h4�Ҹ�[qĀ�D^��X�4\.ʦ4��)u�z�=T�����k���ː�H�c�t�lZ<�$�D�|/PSt�8�E��=:-赋v�L�:'��m.ީb5�`:W�	�/l��GUK�l���~����Ϳs���!ri�1t�G���9)Ō��)�9la�Q�?=���;��K��s�D �������Sw�ƃ;l6=�� ���[�p?��<��@י^e��Ԙ#ҞL=�7��E�&kDF�(Zk\�jKVJL��jmq�����4{��`�*Ǝ�Hj^|K��R�Eb�;í�kf$��d\�@tn��R��|���V\K�[��3�f���7�9x|	N�~��>��o��ƙ�����.�b���	�{6�JYM�ZyG6����4�
<J~��¾���\��)����[�D���}�u��c�k�A| �(\�<�=zi1�Z_��^�|f�gx�tu=�W*�TN���
S�¤]�o�
�_�#�f	3�|C����"�ȼ��A����뺈A�O�_���M��/@�^������G��=�ِ9�;'��D"��~������?��L+gp����L/�.�WW�s�1��8�>�4���U
�0�ܟ�)��r��]��{V����g.��,�)O	h^I�Y�/���Y=�F3�ϥD����Ǧm{`�u����Ƙ��Q���m�C;q��l4,r�xK��b�ޠ	�ܙP�H@��49;˲�������k"|%.��VZ��s����� 8��U��#�L�i�4I/_�z�uqM������E�Z��zV����/~{��k����,Ѩ�"i�B�A�A/��iBI����E���c��x7಩����_ot]�S�x�C�g;@��U"�����P^�k�2#����j�	����Ŏh!é�q�_\���Qf��3��*{h;�@i	���[l'�D���\���a��
(�{a�3ϼ}�������F��v����R~�N��Bf�Fӻr�W�j	���zU��Զu��jSͧ�ې7OtQ(	��xd���J�#$,���p2���u�JR�����s��Eq���Kq��B�V�ځe2��O�٧;���`�82c�tyz�tI]V�D�8�k〉�w�sK�k�����1���b4#�P���7�2>=�Ě���3����Ng@��>����ϓ{�O��
Xb�Ou�mYU������Zށړf\�F�ƕ�{��b��B{yWq�}�o�(�����'�t Z��o�� 5����	d�j�9��ڭ9���<"���B���[f;&��s�m:�r����M;U�������f��r04����_I�i���ڐ�V��1���+� 5?�f呐"�-�§������"A���W@�L)�q��u�ŕ�>���vG�tL���M�2�t�>FDY��^y�2/$�jL0��m}��tQAr�;��z�r���<�2��/xR���0�b�7�|�����W�%�JJ��&]{M��.v����sa��u*w���LXI�{#	 z� �˕Ϣ|�'��o��D6�� v��+@^�Gd�?��Uܪ������JNxf����4WS,��.��Sߒ�?��q�nT�#�$хC�y�(Z�
��Nٱ� ��L����p=VG�,�}5w�x�Μ���[H�yG���)�O�$gn̺f��Z���������a L�`l�k�9q�v�>��k`����v&t������B��6�5:n���Q���)2&[Z��GVd�K���q8�xᾭ0�/�h�1�»�TCj�op�c�']�:�.��(�l�
굡�]���='!���҉��^�6�h��Re�,����;x��-t#�ʘC*}Z|��)���8A����
!�1Yu���=�oЦ8Ԉ
'f�蜱��w�0R�Wo�α��"��ǉt�tc�ҫ~���tEMbji�{q�4�k��e"s�Y$��=�[�܈n��[��[�a_d[Yi������9ͿaÓ&i�:�w��'�Q��By�jS�
�x�bF����������rD�����Ղ��5��4�k��se� P�jJhN��4�V��-j.#�&�I�{@�(6$��W��9K|�;�c�C�'���d��l|OZyĹ�]4p�W�9b�PhG���ƿ���>��;q��9ބ��.m�u�Rz��U�n�4+ ��]7�K���W�L� h��G�O��������$_��r�Xt�8h��)W����oӖM��S6�����Gy�`��cIe��v�[��
�=(Z�Im� W39:�(R���-��FiѪ�<�m�l�]�D��@���k( s�c�[���jY��<�_������ڣSx��:�B����e�0}�DK��9���혚��T���Wp襳X���C����������}�P����ű�� װ�2ol+�i˂��M��������{�ͳ����v�tGʷ��1����dݏ�#�5s1�0Ca����2%���k��s#�3e0��Cd�8�!�����
�/�X̫/�^Yi�M{/
��\�HӠ���&(��T��{/�"�&�G����f��G�^o�T�q@�w���O��N��{ϒ���f�߷�2��s��m(��`gy����7���ui
�Ta[����m<����8�*����
��K��d�.����Ez˛��Ph3��x�R��ES�r�F�]�'�z ���wH�0k��Yyo)�<e(�T����6I_�b��G���M����&��ʤZ0;8,�J�.P鳦8�d(�w����3�J�ٶA:�5��Ej��cQ�+�_����I��c��b]-��E��A;�#�T��ODh����������ҕ�(!km__���U����~0% N����Tcz%�����e�6�5�~W�
���{dM�^+amr.T�g��n����}xK�Qv��v(%��F¡q���\w����L/�Z���������ߧ�!��4���뀼�8�{5Ka��;�f��ji�ʞp�d<H(������M9Z������i�X7w��}�Ӕ�Q�`s�F2�Y��`�B_Y.5��@<�KGu��ƪ�¢�A�x�W�V��i�g!e�S���+l�S���;0�5q�Z�E���Y�ʾ�K۠�_^Fk��C�|����Χ������k`]��Uh���'���#���A�� �@?~��D�nM�Gy��!/��3)����0��ֹ��p�NO��?�g1 VT��D��u4"
�r(����z�' +�)'*��(sĮ6��G�D=к�Zw\N�Э�� �s����1i��qª,F�Eh{pc쟰�Y�$B���0ɽi�1g]V��FFQ�n�u��|��I��
��p@�|�Mo��̺�?�N��"��Q��j'\v�^�P