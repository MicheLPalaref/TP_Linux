��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d้�^��r-�>��s �8������h�Tw#���#/�x%������N+*z�ăZ�4;L�
�Mrbi��x]5*�j(\��T\�6e�C�G�x����UKD �8���*�`�U{�C�;
���^�<Uw����^��DB/j��,>��(�)��}X� EV�o[s�J�~D�����ӘFy��P�1�ɂaܾ⓭X�����j�^�T��W�w�C/�ļ��7Ow� pa��rᘸv�9�(<.���Őh�Kڬ��k��;h����lp,PM�Hs�5���Z��]Y��2M��1�p�w4� ��\G�l_���0�U���'��i�H-��vv�?��04�m�=��3�hh|py����s?@����zc~�7�lw��Un�b�$rx���!!"ۡ���.��V,��h�� ��Af�v��{{2} ƨ������2,:�q��Q���b"CA�4<�Yk���l�x-�7�	v�fx�}�qD5�:��L�k�ת�s��E�+��o��Ɛ�Ճ/X���7�	[�s�k����(�L	��'۽ԓ��W�0Eh�݈Gn�S�>�C�rԁ����j-��Ԍ�g& fN�����[eb��"��������^�4�sa�u��)A��~6�Z�j��ģ� ����[��c8*�_��#��'P /8D�1R���w��t=�"����F��t�i�Ƴ{�;��xC��N,��hv��>!U�q!�Hp��RY�	���,8@j��z����y�yI�kҋ[_�K���_��Mc=��6�	�GQ��!�<j�0�-����Bq�A�G�ph��fX�����<a5b�:��6x2�K�)����'Z�zA<�K�6m�野��fYq�K�r�=~)�hF�.��n9Vvw$ȭ#�(�z����_x�"j�ˆ ��B8�b�2;;n�Q��>rE�űLo��g�,8'�6�j"څ{Q� `���כAR�T��>U}2F�X��3L��"45eMF/��"S*��;&��ÙJ�pi|�b��C���U:6W�N���@Λf��ja������y��o�v��K�&ڄ�!b+�D�?�xF%����T$%F��*�ju��}�ǃ��}�?� jǽ�G��y�un>�'�_<>�L�s�]����E��.�S��H&���݄��SfuwG8�,[0����{�OT��qcZ`p ۤ�u��:ݫ$�7<'�y��7�i��֥���Kw��ё� �d�@#f i��p��mt�������v��q��r��E
^M�?���c�_:^�P��>ލ����?wj{��Sb����p:KFG���F�%xt 	�+W�N���(�G��;�E]Y��J&��lU�fX����G�ռ�c5�ݤs:�ʠ,�
$�ѵX�����#���g�8�J{q��&S���>p��U�%�-'#L�Jy�9Bb��t�Q��u!N�/JLcN�������Ǖp�M������� ���?�����s�]Y��GZCd*U�}~�'�DIA9�`e�?�K�E~e��_�є#�7���`���4$A.k���_ivH:B�	!�& �Mfk�3��,����=�~�p� �j�?���I��踌�C)�吾�X��40��P�+�=���Wժ�Vo�Ы�o����<�
���9�@{=�H��ׯl�g~��ɏ�d�j���'��j�3	%�!�\`%�nf�.E���pX����1�A����E�ט�����,2��w�Z� ������1�&ץ������q��j��\Yp!�G���W���`�W�^���wk�k�$�d��u���I�z(��G��朒yV��S�H��@ּ�:RU!oʊF��9r����+��2ʚZխ#�w.be���N,��F��߽�b%s�T��=濁}|�|Z*X���E
�Wִ��%3-�d�]Rz���nꇁ1
���'?Yk�vݥ��S������~����B�E����<?�2ɖ�-��F)7	��V�����] ����v��q���ا��� !���DTW�d#/��o�����}��>����t;f��s� �Z"b�� �¶�<M�nC����-ʗIX$��+#�ơ��s�$���В��]|6��cm��4X���Q��$'���?_+���a����X�|�l�VQ�(��4�m9�{>��{�b�*9��3U�6�����7yӏa��G0�:��%�T����E��X���V#
�)k���aR-k�k8�+���˽@���Uy��r�6�LL��9t�씝��Z�e+/Aev��b��Z��o��N.{�
D�G-_��2��k_�,JZ�ԠO��_��`�#���3�Z��p�x_LB��c�RJ���֔a��ͩ�q�ƴ��I��l	�O�Ap�	'#��+�ɠ�p1��>�/�0��9C�����	�|�`�5����]���uP��ȅ���s?���@Խ|�ѣ��C��9��︙2�,\<}���d����a�R��/�2���>�Z�����5�����_�����Ж���uʿW�a�c�~�{k�Ѿǎ�vH����wf��Ȳ�q����Ϫ�܅��j����m�@��*Q�9�W�� �?�c� ����uo>	�9��\(#%JGE�q�[��t�.8�X��fY߃*'H"��c���T�韡����8k�z��`U:�4��๯��]�p��Pw�1=KH��>��	@"�'��z&`�.+��_�oE�R�%�oҖ��\��w��H�1��D��y<i����d��t��R�e�X4[�Q�|ـb]�g.*nb\����uA0�l���`��o`#��9�Q��G�~9(��q�B�
���*?�S;��Z�}OAz���rF!�o;����#�o�"��!�T��~-�N!�O�����g���\������й�lP��T�b���9hp�U�I
���SY���sM��;����3��ĕ� O�j�|�p��pv4t5	��'g)W���?lNeR���.���p��Y@@6�����%l-�u5�	q|��c�AjLQlѯ4Zד�Z�a�n�<Z������FU�R?��Y�{<��_�E�ꔞ{,���^�c������%źi(���W-�TX�$]q2P��d�.1��X��S���O��옽W�0c��8�n죗A}V6dG?]d%��b#KyE8� �Vt��)���D ���m�+��)����vѴ���CdҶj;i~����l��0ѕj=�3�S�9�h21�վ|d��T��<&ęa9o�Y������x�n�ƌ��<��8�jQ��C!����e��Tr�1ak�K"����MOO��[�Ź;G�P���q��_NN�#I�	�Y���^���
�(�������\��u
x��P��4D�Ą)Q�}t���\�h�1��7�ᐸ��t{��4Pi"�����	j���0=�G�4c@u���Z��ii�!Ό�m�_�X�Ÿu�`C��p��k!��I�"��Y��g>���f�;|�Ɠ!��w<�Q�G�[�1��X��L�=vؼ��5jj�*�}*7wؿ��#ac�F�E����`o{��b6ֽ;�5�Typo��Yj��@O�Vh�cX�;��Kf��aJ�'��H!�W�a�mU-�*���k�+�5Ⱦ�b&v�1 `s��^�Q�N\e�!�]dw�9���*�!V�gt��t9R��^�X+�9���`}+?�#�¥��/��4�ӝk����:H�z�.�R��k�۲��5��X$^*s��~q��ƞnI�NwxsL������7��r^e߼��\�B�Ch�EX��G���:���Y�C&?�9f����n��t�4�ɠx����N��//�ڐ-���M�Q�=p14��O���dڦ��I���t�(㒁�P֝���Z�E��]W�z8��}&P,2��>'�F&"ح1E`��tLp��o�e�w�X��%u���M�Ԥ�?�FU{�l"��1������L:(w��&��<�ɋ`?��lӶ���lG^�1,1��p��kr�0����j��"��.<)ʊ����_Ԙ4�nU�4��`�\PK�yȥ���[�:�?�O���e�5)a��3�"}�|�Z�f9�T�Th�=Et�(��9��f��-=>h]�,)�v��qAQ>-$��m/�HM�I��$Ց��3
��G�O�W[�#1�T�	��
�xR�Uʚ��J��!F�D��.�5�V�O�Q�1Hp��Q�(��vo1�4<1+�l�[��뻞u�އd�'j�A�AI�Wf3u�x*y�X*?�s��Dĺ�of~��S��B�̆�0�l�F���sm˴\�8R`�"\8�3�+&1/���-6Qut��a�(+Mد(�Ν���ލ,��<K%C� t�����4W��Ȫ'Dz��)X�ʽ�����8���}S��Wm=���ޙ:N���zF��@���n7^�_��\�$�=K�⯰�ܖ]
���#��H�,�^�1+a�R\��ې=�&	Ne��,?�4���5���Y�D#i�G�S}�M��㡖w��)��3!0�G�a�a:�PK$&��! w�m�اO-�� 5{W��>�osUW���ĹT���':\�q�tp�:�&%�yA�I[
��(:&ʸbS��vf����F3��S'�fX�������~�j;"z���p�?�3f��!B�~q�#�0���/
�f��s��:��J� �v�Q�G�%�>�<��bMN[���J�6I jFXH�ݡ���\kᆾ�IIبS�.I��[X $��#K�*���ڒ�ޟ_=�`��b`�����B��F�x,oyFm�"AY�>?De���i\Lo������n���;�i��^xz�p�����M��c1�BwH�$�I��uQ���H����>������8t��[�vy���X��To�)�%��:F	a��i�pƾ�$+�@T]J�$��V����V��񥄁���+K��H���N}�K�V�����R}����"Ԙ�m�e_��
w"�`�����ɪz�ϔ>zm�,SL�-�חo3| ���jΏ�"}a�B
W+N�PI>:�{��]p��8���q\eF��_rYn��d��v-�.!do�M�VUt W�I�wכ��.�S�9*t*+��9�5�nݻ�U�Mu*������d��_���� ���Vs+��w��D|�{��Z|��8�s�����ؒ��]*{,�t?d��v��}�x�n��}�+�U����/u)�S/�f������Z�R���f��犾Q��u��e�Q��(79�.����r�)�ݰy��x$X��uOD���E0Xa�}�zO�=���m��&Q#��(��Ը�6���2�K�w}#��61FM{oRh�����9�Ӂ�qW�t�Ov�"21�3�V:�3-��U�� 3��/�c�e�E����|���a����ci��L�MMڂ|FLޙ7��ї�
�<PT��c4�||�8Ӯ�D����eK�ghI�u/ۻ�΁i	���-�+8N3h�M��<�W���ӷ-��rJ��F�јw���K����hr=UR(|<�F~flw���{_���r�{(eY*����*��I�=��+pcÚnA�KqE)�A���ۀ"�N���h�Y�D3�?�\z�~��v�~+Xj �ح�}�M����"ڞx:pH �G����2�MKT�I ��{O������3MU�xS�O$Jx����4�ѕC����<ķ�b!E	
��F��D*�_p� �EÚ�:��2z?|:�m���xn��1��_V����sʠc�\[=B?�g܁��_c�M!�v	�=�b|�"��o����OV@�����Ͳ`���r�2�s}85q"MN�;.+Hr����)�.��m�e]�{�p�ZP�Rp�F��\�ݝ7�/3 �Җ0�8�!�7���V��6�c�yi�(�yE95��!�,����X;�
�Z�2�̺-g"��s�b��O�r��19���d.�3d�g�B�.=�N��0�F没Y
�ޡK�Θ��(��?�r�uч�ވ`�0g�HE��i�X�G���N���U�"\[x ��Ms!���iܛ*t���;�ђ��W�����T�g'7�X^�����  '�Sv��	FVV�Hv "1+�&�R@�'	��K���#{Z۹8��#?3�M,*�մ�k���5�2��]�k�t��tL�G'��&�.���ʪq������|�Nާ+.�X��X��|-�؟h��*�]"��߭`բ(F{�(k[v��I�����>%�y�M�ψ��	���n�x���߉lݲ��X�.�[�����ψ?<�� ��}(����Hp'泵�m����l�H��_��~�����.�����`��|������Qo���<-�v�	%�>�h���{�L��\�ڜ�
��� G��K|���̎��FA�W�a�����;9hh�"�_�>��]�Be�_�'j�D<�z���
�ŧ�Een�����ϩ�_�|��wL:A�{�Ƙ�/Ĺxa�Qm
B|[g�L�k�`��I�ir���-(�z	� ��wS">��D����aș���\��;�HP��ȳO��[�e`�\�F�L�ڹ��i0M.�P?�G�����V}�:�]�K7%�Ā͐.%F%�4ry�+4�|��CW�j�\u��H������W<�]E��!��8:�W�CήF!��nBT�����D��ӗ�^�K�Qch)������"��ȁ^�W%A��S��3�>��Z�*Yn|�8;Z�#T��oW;=�]2F�z��f����@�*q|�5%0�1V��2$��٤-��Ox�l��yu�i�N��t	�Ҵq�H�z7�VM"7M���P�+��H]��}w^Z�\�a�5ݴ.��̱�^BPQ�&�!�~�m>Ȏ��@���;qd $w�N?��Y,̩�9����#	͚����e�?��wp�0�7Ia �y���a�{����G�q��T�,B�ף�ޱ̕���j��`[�FǾ��CҼ���*�	-`H���3��ݾ	^���L�-�l����밤�������B����#���_��x�e�$t��}�G�Z�|~&�/yl�BBʴ$�y��)������'ԭ~x���a�� �����U���K�o�Tj.T~/����./B��ؓ�B�V{��iQ_iP�^���/�u��8�Y+~bg�#����UC�~iE��$UUY��;I�lGv���3֯��[K�d�Ox�ԯ��ךj� 9�i�x���h/��m��f��7��n�]~V�%�{��?(2�:��}�F��Kq�����&l6��]�?ʹ�c�/{�WcS9��3����mD�װ�v����w&�	��3Q%�;�e���S٪����@v�C9��C��Э�~%ق��y����c���"���.�n��|��j�^ޯ�^�C3yY���K������[ ){f-�</N��� �[`I)���EU�k2o9��kj�����绗K���f-0����&`���uv������Cy~��hx[ڃ!��)J(�����9Df.������`����7�%ѨTe�:���ыi���dM�9���X��;��RϺ,��et��[@l�DV9/l�r8��R�:��������zF��ս��8H:ؕ�|���7�:�u�Adv���m=�B���;>aE��qe�������&�Z5@$_	p6Ov&�Dh0�8��ht~�4��6t�g�����êP 3Ka!.B��������78t2���Wv�������%��J�Qx�sdiE�����tّ{;���2QE.�̥&p=����5[�-ot?������7ϳj?�jx�7�r�Ì�l��_�݉,�j�-̃a*'�#,��r���/d|�L�������Pxw2o�i-,de���[bҐ8�����5j����j��d��'_;�L8z+�U�lv��WY:	#e��w�w�:�3(M�ʩ*P=)6)X�,,[@ea|!�@�߀�s:�)/��7����������u����d��`ғ��_g+K��;�����W�����t9~=�U�.����c��x��s�p@!�@)��^��ucn[jq�0�����	��t���dx�/9��2�p��w���[�S�R]��<��ޫ����ʸ(5*�6�8�0�RQ»�����Y��?gA��eR��\�x�]sӲ��X��0L*�e�6�HX�7O;��/����v6M=���A��)�5X���}�h|?^ȕ����<��ƲUCC����.At&w8��;��*5��9���`6��)�`���|1<�(o6>�8X1Y�w�'�ԟ�6S�G�K}5�iΛ �D��kK%5G���f:�Am�ܾ��f�<��Qq9��?����L_�a�s�S����y�����
�+�*�������1����2V�G1�L H�v(d�A���fu��@��q���Ч���v����E��@�kD�p���u)�4��J��=e���%��v� t�b��#��R��_�`7?����+�+3���s��;�7�J3��Lw�K��׆
�:��YֺDz�$''��P�Ĩ�
t��2~���V�����|4�w����)Y����В��iZH�ZT)���d�D�
���H�Or���{�$�EW-��PP/�	�g�$hſ�d�:�A4WP@"�saV����R ��W�)
<�pн��C�(3�[���N(���,]D��Zکݬ�����321Ś��`2m�):��\�l[�Jp��P�Q��ʝ8_Ge�(���
�#�P�*�3In��Ro���է@<R���3Jg��3�B�RS���I�#Zq�bad�2�'^�D���C<���9��ϥ+Ǎ��By�$���-���5R\ʟ1P������zKuxl�f�v���i4H\���}��5�^�OaC��a�K�|�\[��ZR��T��h���+� yz�s�e����t�ې[��N�vՌ�]yū����\s����J, �������>�J�	(ϮocB���:�{���;G8o��kq��?	��ZruQ� ��\OՎ�LYKgW���îf��Ѵ�Ě�f�>�}�V&�ʓN����֐�H�h'��͋w���l�<��	*R�-ߒ�.���l8�:n�lQ^7�����2^�=�-�c՛�6�:�~q��{?�����P��;�ry"%�*o�,�\�E�R�[��gm�ͤ6�"�c
��i�=��?͉i���=�k���S(S20��.ָ���NKV��i�E�i����6�9gح�m\\RT%�������$���l�h�Ktc����E�g�.\�=S�I��uAq�{����z3����] �DED��t%oҏ�$�E��A�Rn"�C[㻽�<,�o�T-�?wԇdkI/�'jp)�4 ��L^�	�@.�}����&:�p�C8,v�=jM����Cap?aYȋS]�4»;=?*j��7a�xX~��4/z��;v	��Җ�T'�EE8*ws�I��|q�Jad�D�"0�n���*N��6S_��#�'>�)ZvV�F��d-�M��ݱ��7Q��Ō��/c��]��Bj"Cs<`�(*JLx:�=��J�Y�b˾t�` �GD��^JD�����}f\)~J����8Ȳ�9��.�S'�A��e��V>���oRF0&w�g �e�z�S�$.��f��X�ud����)< ����^̭a(�O���A	qZ#���ACjR�o�K�wnE��V��ZͭdV>[�!�;���dn���܈����ǱL�Um6Q!$�͸�΃/`�,��]�rt�B��)\tX.Q	���6G\��ӷ���T�=G��<#0i��E��⮦kH�!y���E���\1����)r����MݟG���s}�r?�$� ��F䱨��Q�Y�tV>�ׇ�*��M8�rm�Ѩ�#��7�RON
�B��A�ٱ��齀����g�d�;ZKe�?�����l�P	i��#@���[���yL�<ҏ��r?�t�@��"
�A���Q�ʾN�/ڪ{}p�o���q�(�v�v��rT\�:=��{��Q����=��o<*�i�X8�����jɶ�:@�g��K��0w�-�q�@2l���j>�5����I��[��;��³:�����g=8�4��,�۰����
��,SZۃeT�#b<�*���U�}5^ьv�O�����X,�,&�2f��sX��T^`�Y��p5\���]�t
�$+Z�r0��nǚ!�$�?�|<�F{�I���� *_̙
�7�0~��$.&��9`*d.���^cU���h/���eWހm�Uz�[/Lc̀9���YOO���Ct�,}�.}?'놚r��W�p�545��RW+M<tbpg��Ƌp 9["h$.Z����<E���z!s���G��|��<"ot^J��j	�����mI��NE�*�t��a`���}'>���,'� ���w�l_�gO�6r���6����)���g����R]ec,�E����@&�z� ��*�5|zK0�fYk����wkō��H%|u%5fF��r���b58�Tր4w�5�P8��t�>���f��cW���̀�J�&��*���&0��N�	՞U��)ط�(B{���t�H����!Ƭ�����������'�+�J(�� �HݟXU�j��d?���go���Ů��̾A��1C���cW³4�v�b���WǦ�J<\��E6���<�kX;ENPe�6�qOڐ{/g�p��9p��`�c����h��N5W�nfdӠi;]U��u� �f��(z��4�ZԚ���[n3��ޝ����&9��>%��
�1��!����
A�2�A�I��o��x��� �JM�gsa��7�mIn�յ$�T��O���֣�>Å9�]��LC�oN��g`�,y_�ϒ,=9�Ȏ6Qn*DV��-���c��H�R.z���鱄«��Ӵ㉝�R+��� Pp��n��B�[���%ֿ������}w|�[�^���'�K �| �tl��@e'�3�S�Z����D��+��̱�'k�h�'��~6�ˋ�D#��J=�J&�n� �wU�F�I1w{옃K���Z����d ������gKfj|�q�҉@s�m$��'�~�����F�/�N�]ӅI'(�1܈߈���x�**Tce��Z�ײ��3Ϟ�#��$�W���V\A��-��\7'�CWs8���	��Z�5��RbN5��n�,�U T�w�"����#��UXz�ͮm?��6�+�����q
%��p�˪��:�q��ϢF��CG_��i	��l^>n*�#���>^���E�d�]<��V�Z�Γ�މU���i��+}�X�.F�ߤP�M[	�9Zi�@������MK9k�{��z�#�|ti�J���t��w�����tսN�A=!_!��7�/�ڨȕ�Ao����Q�7�f��}�a)��3�j�JEQ�å��0��qٽ4(��,�oQB��iuf=6�d�:�C����
>��5X�~�J΅�$C&���(���Ư�"�gS�L�[{���b�<� u�uG+�ں5�Fp�ѯq)��me쇏��`���%���*�	�T�2�Vt�B�vz5
��Uh�	���d�����o���b	�k�rI)ݤ���Q�h�E	�D�&I�N7p��os�{�T���[����e�OZ��̞��w#4�&��²1�Yr�Sy�4z�)يO��3��ٯ�R�Jwd<�[�e�AnF�"�����0k:�f)��<���Gfl~�L�	J�����|���w�a0�i��qT> ʩ�rH�T��g&CHS�?���j�����E��6#y_�7�5W���+����`I��J
w���|����\P�:%T�L{?��4��rw1���CNv��b]E��� �<!;��p�
�ElC�	�G��C�ӣ���u�� 0���MC�!�͝�a��{����x1���?Z�H������꾏2�!6��zJM�C�{h�g*{������|t�އ�.���/�L�H+�������lve!�{M|Ƅ���--�]�B7��~����G�N��E�h��7M�j�a���$ުW�3�ɗ�Iu�y��GVg���O]���x�6�̓ưk���w�Ըq�W�"�$&q���(�!-��h3W=���y��>}o#ڃ} ��OF?�~'&�s|I��y�*=x�a�ӹ�� ��h�xa-�ڿ�>��E�� W�d����N�.�;ڝ/T?!]�U����Ӟ�H���EUK`O��|�j�ug�-Z�@q�+�^\�e�CU����xm�r���)ȧ�rT�0���I3�p��P�O�z�;\35�%4?�Šႈ+�8 ����g9W/�Bs�j����6��1>���Zc�Lp@Υ�*y�W(���	�6	�f�5�N�z5�kK�T�TJ�&����X�^����~��1�l�,"� #��ҟ��'F D�J鬨Ų��ɺ�3�I3C�ݤz<�b���mU��1�7��ҕ-�U΀7��e#�N0�V*T�1G�����r`�w�''hn���w"��	�"�6���5�6�hq�f�D��_�)~��Sjp8�7��&t����ș�/���xr���gp�.T?���[Yh��w|���0���M�;r3ٞM�]Xj#XfL`W�g/�:�=l/���)G+�2{d��yH����>#w�r��S F��еK�K���F2~S�O�z[ �i�౬��sa�P�2��ĥ�c	�=��Ïm�ߏ3�Z�f�q~�B I�X�kI���5
�"2&�;Jc=3Hٷ��߹`�4��ЮY6B��0�F?�f��bK�ㅡ-`�y��.ģ+�5kʫ<���9&(Cŀ�wI�w��%� ���_�=�0�0�]��Y\/�W#\�XM��|d,X{�u��_8`2 �[#U.SB���7#�6��� ��h��	j<]-��F�$^��+^z399�`��'�uV�9�`4(�i��U�Cs;�!�3F�z�[4�z�'��.�}j_�KY��g�/U\6��HV�jt1���RRO6Ra����|@��;H8�'�a�A_�L�r"C��?�F_Q��xt3�o�1��yM�G�w@j�>12M��n�����E�
�H+�!�J�Z��:#z�k�nvSΘ}{OA}坻ـh28�<v����Z{;�:F�'�ڒJ������;ߖ�e^s�-�>
��|��&��٣��~�wB��c�U�X�^�g5�3f�C�M���.V�v��+T"�P��&�QJ�y�^H�TO�m��D>�/c�U��m$���7Uύ�T!�
p�|�H<Fw���������F�^ص�H�.�=2au��7�V�Eаp�0�^L˿;�j�VOT�k9��Z>]�jћ{g�3m�{���v����I�Zd/ϐ7�3����zi�YX?A���\�f����>��(��D%���[�Q�o8���\�d���=��[D�����������&ƾ�aBL�$��1�B,!{���sbɥ��/K�5�6�⥁s�HF폞"��(�ު�57>z����u1!�����>����t����[�0.�LO1��HV�>^y`V/�W��E`�}=~��Q�L8PE||�/֧���Ν���Է����|_���G����n��1"�W�^�'[
���$�aU~k���&t:��8�=����Pq�1�vro����ah�d�}�].&5]�:�v6;�F���=#'�ʒ캪W��cͣ��Qu�w�Ԝ�pF�H;f$�e�k���$n@�sz�Pd��T�G0V�����}��g73;Z���6v%���e̙۟���;�a> �C�V����F�{L�f�������RgGq.J)<�rN\��j�t�1��)B6��Gd����z&��`?3Cx�h"=2+n}K#���)Z�k۟�'?����!NU!\��a_
�NE6 L��']��s�E!��4�V^.��f��r+���:�2�����Y����7�;�3E��\��.9q�w��P]:��v�U��v��ov���{�R�g�j�GR����⫵��'E�n$U)mO��zF�ͷ*4sY Y�]ߥ��Y��o^o�MDk�]��ӹ�,Ƥ!w6ʪu\гԇ0����� �z�w;��;��w���<����^.�Q3��´ �M��T.tc������2Z��/��4�kA)|�ÜMVx^���A�:Um�#h�OY	z��"1H����p,KI8�t:�4��r��2W��[�����?�g�C�ԉ�5�f~�Ȝ;���k�FW� C�`�^B��O�B*a���7�q|���A$��}R��qc��P�
���G��"���
Z{PKn}���&�V�2 ��T�)�����{�6OJU/)��G�)?���Ş%2�٧IW��2,����~� �%q��Z�E�KM#f�;�-Z ���{�Üj�"
@���V����N����{f��Xu�Q�l�Y��4x�'[n�p��p��r�R^�z:�qeEx�絰 %��[h�ъvV�ݚ�:灁��Ϸi��5	&YT�`�Fb�ՍK�JYFSf!�ڢ�=�]��w����Jy��m	��I�S���\�zĸw�!� 1$�n�v0Q����nˌ�z������ 'D�[5u��E�=H�=~�	/���v���6U�OL-�.>��m��+��EP�ۃa�(�X�ޖ�~�$�8:����R	"�9��̫�I#��!h�G�0��e�qr"� ��p�VLϑP�Y�B*��f1��	[�;�?P0�1�70䯇AW�0De��|�%ަ�VU�!�xd���\^����ϲ"Gv1�0J���<��碒�}���om�
^�Y3��c�6n�!�r�rvS��)[4OJ��^���J�v�p	)��!"Q��捞��������ˀ淀�7T�ܭ������|����w�Zۭ]�"����x	��8��J�^[q����H�ֲ�����'v���b�զ�m�5Y6��.�)�����<USq��Z�H޹N�oH%����s�M������Qk�\��$G>	��ؑ7:W��J�RP���1~>!�yx����d'����3�Bҋ�٢|���G�3��b�X$���N�1�E�.��г�ڷVt4�Ӿ#9+�9��$S;,��7o3�%KYhm���6Wb�!O�CWt�D�E�=P}��"�����}?��λ�������V��Y�x|��E�R��	�������v���S?�?ط_�\���ȧ�RS��GTN�w:�fS��&� Ǯunv-\���Et����8��d3&��ێk�;Oc��4/�U%�CX��a�	C?�A��K?YŴr��н����G#���R/}��O
V~�iwZ�pt�.o�6b���A�J1��Y���Ui�^�	L��r�So���lUxϺY���
�������R#y�|F̆��^�lI\�L�@�����w]��23�=�[�|�gPڸ+�$n$_����SLka_�Xϧ߂�GC�����7���^�'NV �Ѕ����+�.�ePmk��UP{e��xw�?���dx��h͓�I�6����nT�k��*���j�J&�p�&K�=�1�WβL�j�e'�[}���K��B[H{� �v�.{�� Tf���.?J��=#�>V=����t�6H<�Uf����Cl�Ů�*(!���W��P� ׵c�u#$�/�����lGiTtW�xOs�*���u:�U> y�¡6$7���P��f���kyeHk ���{_�>ʼS�Dρϒ,�(�pA[SݚG�]���ms�$ӹ�>a��kN��l�����Q�T�A��?�h�O�7��&Y��/u��7E9���h���͍	��1JGt��$#�N���S�:,c4�� ����Iwj?b�_�F,f��&���S��ND$�j{k�Y��$��짴��4���Pa��T���|jܫ�k���bh�Ý����eu�$qJ5��`w�ߓ,"|C������ue po�O^	-��6�OT������RW���ܔC��C�*���,�ŗ-3N&(��eA$g3�{a�nV[ �zg��D�A����w�Y���d?����6��ߦ76���|��(�>�Q��׎��5�1l��.3�d�e��4��Ҩ�ā�W�YGM�UO��N�:=��7פ�Lc.]���͢�g�)e�����-T�c�z���x�a���D�b�(6D��oc�!v��	ٹ˔<H�&Ǻ����Φ!���l�Ҷ|^nD���z@��@]t��?�����w�3��ўL8�
=�.�[�G�l�V�.n?4a�5&��&�\c :��]�aH04��!+���,�s���R@>�c �@.�ϱO��՟��O�CC*Z��:'А�w�RL�H4'�B%�@�vAfʉgHܜ�ZW�k���QR����F���-F��4F��h�NI�1�7�7-{ok'��Rw���0x��9,}9�P}L�"����]h�ڧ�Yu�Fрt���8�\1eft�vSr%�M�pkG%���!Yܺw{!"=<��I\!����Sp���1��s��#.u�<�~�����B��&g��%.�b�3�P��6�4V���;��9�`�Wx����#B,��#Ia����k�����-�Dv����8������^��W̩������)Op��~-�yrD��
D�H�������o�MJ�=�]7� =]Y1��wM�#�g�DK{ㆰ�倧���z?���V��Ӡ< ��/m�'F�z�.���E��=�G�)�G��[�G�I���t����K�۪	sN͠�qԂ]�6�(g�M�X�"Y�5y3�H
�&VS�R\>���S�Z}r8I�8ʡF��WMTWTC� yHE,�ӟY�N[8�4bt�ԣsAB{l�f"���Ă;��e��&([���)%�E�V��i��H)N���:S[-5�����=[E��T�����m��,܊{c��pDU�O��}�د�W����^��d!3�?���w�ÀJ����r]漵$����v��twJ�=jm��_�M�|��(�Z���A��pR�3F)���Q�+�%�1�{r̷�tu���u�3bO����%Yݠ��As�\�����>���|��D�t��k��.�["�Z�EŘ���N
1|Q�m�б\���ك�1�v ��Ƒ8V�3�5.b�LF �v����V�IZ�<;e��B�`^�P��Ŏ�V�;�*�
����ǭ�ʇ�I�3[O�6��!#��V!�:�~��P�z����n��V�)�b����������|#�N�h[ �>FL��$fa�l�my���D��_���L�8)j��w�!#o� ~��(*��]jN��}�pS��>@e��)U���,��4D#���K�9.�e
�[��b\د"�9��_�F���>y`��H!�;��W�K���uI0|��x?��8��1��&����_���h�_�F�L�~��b�E�N�� �R�&W�B��D��6bg��{>�;;'Q^UV#B՗�ɉ��p|�gc�
�§�����=:(ˤu©�(��
���t�7�nE8M��\��1�1~68=Ĕ����
��k�pk`�4��m��o�ѽ �	XR�H�L7r���o��,rn-OD��X��������Yo�|�����N� (
nv=�&7�ROt_[�Z��+%�Bp�D{(�F-{#�^��/@�G"B给�̓5���er��ܚ) }+�3°Wf��1~\�C��є5C�f(��y��'D�9٭cW�c;[���?^xf&Cp��p��S�&0E��@�zG����܈�pJկ��	p�ͻ��xWd\�?�6�VX���&p��A�-Q��xSf0�t�L�
H8*���	��W�_�A04��7<��7�*���0u п��BN[��9�nx��Y�J��!���]�u(@��.P"��h��+�q���~�����V{��.�I�ie���;h��W�>�d����q@.N8��[�-�6��&y�ҁV -<F��n��B7�����I! ''�~��'�&�E�f@�)�BS��&�/�6�^.4QN�����w�������9�M��,�Ri3P���)�$�F��g��53�j/��u����KH�s3�$�1t�/���c`�=���ہ�jQ�W%$�A��{�wg���1{�����ܔ���|o?_OH����q5�u��V%.����/�@�7j��t2_GDu1��}���E��j��!�d0h��o3la/L��j��J�P]�	��c��QmKy�é��6R��zWA�R~D�v��.1\�<b(��V�7�Nh~�Q��w0M�����k Z�t$AJ���Q�8T\!o�g��.���o� "ȓ���>��5��6�<m>[���.�B��*�R,$N����-�?`Eu`���c�;r_Yq� 2<e�c���30���?_��b�i�^_��"'�&�r�H_��wctG>�z>r	C��1H�Ў��nl�g*�jδ�Y��΢��N� �p�+Y����_~�r���*�HR��V�6��V�u^E7 |q�2��A�le�é��<w4�˅�j�b���k������̐�Ѳ�yHo�R/	 �[sB��#8�)#[�X�aI�裷n���\KԵ�����c�<�������`)b=�:lϴ�UP��M� L&�:��|�ƪ�c9~�J���Π%���N�-É5c�G��$ۓWM�j������KNr�)��3z]%�W�L�O�e-1/���:���Y��	V��JY�a�i+R�.���Q�k/x�{��Wɝ��(���y����iM{l�n(�	\{�2;|a�xa��eY���S����-�k�x�EG*��YY
ש�aP��,���N -e�SI�f�~5s	8̂ct0�rM49��J�qC�1�n|0����E+'�[%����J��Ds©<`�Fo����K��'-"a�(�����v�Nq֯|`T���	z�_���!�=2�|\�D$(ys"��٧���}^��	u�!���5P�9�w�²/��� L�5Ƅ|!
|�@ӗAe�A5�'ȹN{(/��uW���Jd߲ՙh�*,XX�J�c���(���
$6��\i�� Z0]+��Q�?�d����p9�>u�yN��S����  S
){{`��tц9����ߌ�V�Z������{X-~�	X����`g��i�C����U�����"���4I&��c2ȷA��w�y�qy�&S�}�f��OF���#�B���lo.?p!;�Ӭ�����	�#J��E��$~�/���n%�qTP�y, �X��t��ӈ�}���:�?^��x^��} �%y����~~	��ZWG��r��[�4��C�H_=���Vr�O���gXf�&-�U򋶹������p9��6j$`^��U�k��B��P�j�דrz��{�+2>��H�h���t�C�K[q�X��8�Q�x|\�6��NT�F�a���C���(ܡ�|®3�����0���N�6�=���&�s�K� ��d�ۧ��*k2�� �k��cx�8�
�<�fI���E�y$�pcPMC���6x��\�\.S�d�
 $=�Ȅ9�SuV�/?��U�u#)�U"o��������"���b.
o��K�EU�����省�dPv<��'��S��de^�&�5�T��ʞlo�f�sb���DQ�3I75�K��݃��B�xb��śvb2�X�u_=��s�K��&���U�,�����N�9�g�9S��M-D��f��#2}�Ŕ=�����X��%��~�e*_����D~tY`��8��Cm�C LC�q=�@�[�ˢ�OLw���M��KZx=� #���b����v<���emv��2�R�2��cyZ��V�u�z�Qh:�C�����M�@���Y��6Q�wFj�9{����GV���faٙ�N,��*�MA8�I��ۏ�*�g4i�u�̔nz�>����ȝ�O��l�I���3L_��I-�DDfY_AO�WDuJhY
�8+H��R��L������$&567/�#�[��u���	�=��\�p�i�ah�ʠ��/d��_�+���K�T�{%���"�6s�E��8jDn���a���ǹ�G��>���!�5�l���XH�.�T�8_�����|X��Ć�*����ה�$�z~��g�܀��㜢��[~��o2�$)�@k���ϣ�D�'yfP�Z*%�z<��"@��2 �8�00%�=��*X�j*�?~X�ɵmf�	l�zc��/��'��Q�gU�-13;���*>�Au|���Jw�B�؍"�<��/+�@�&T@�&�4�5ą�_%!
'�婞��J��F�Ä�4 ��7�bT'o��E)AsCDR�=��<ExLçz^������<
&��a��U�dp�k��Xӕ����N��^Ӻnڍ���Cv<-���p����J.D�\d�ٗ,���(?��(
��6��C����`e׍�4y����`�n+Y����۸�V�kӺ�F��*:&ؤ��/u��מ�k.\h+�Q�c���%#/0��%H(���+�V�9T�� �/`B&.8A(7Irl��2ލݺ����7ʫ"�������(��J�b�%Ũ&=#��խ�ؐ' I�7��pb �n4��	3�yF�{��ee%�q[����Gm�j<|��?��(6Jic"N��QuͯC�aS4�r4bjj�
�?�js��������c�>�u-S��T��+·K9
�/7������
�SBf����+��ڠE�J��ꨔʉ67�#-��r�ZX�m�9t���iοblN	��|<����.�7͈'@�aL�w�aL�j;#.Sz�s!�����~���75��@�#A�{[���jR��w��'��k����Ww3ck00NG�?cJ�����~{q�Mb_?T$�����X`�؊�W��])uQ! �� �NH�t�u��~��&v3<>�yz6`
V�7|��+	:GX����D�7��\��UŰ���@�����Ӂ��|5C2�P<�(Y>{�U!�)�L�{�ը��� ��B�O�.mO����6�M���u�b�y��HPɣ�@�����O�T:�
����;@>�����������#4He�H"�m+�-{��O?��Ak6*T�:C��\��Wp�Y^��:+C>�����54S�Ĺg�)�O���<}S�#3���o�H����u��s�G��^xcuն�v��,�EsbY΋l��|��3!/_kC2m`A�"T
�8q���E;'�K��K�،W|�hIݔ��V+��<9)"�2�Ӹ�&�$�n��$P�)L�ʁ�,���O3½�b{JT�<jx���Gt^i<C��Ϥ� �$��BmE&�l�I"���)�Y%$��� Fbͱ%�ե���c:7�E/|S(���N��J}W6���0qL�M�?&Cչ6�aZKDl�Y�k<l�D�ԡe@��N�ԏ�ei��i ����پ�Мg���(G���etc���R?���j��Q�����/�B=�j�@�$A��
�Z}�e���������.9�7}����H�5�[7_� L!O�@��A#��rUs�Z��u`M���G�=�5�5�m�o"F����V�A�h��xD鬛,#y`j_�B�Z�?a�0EP�QC���B^�xI�s�)K��*�Eq�b�u!�g`k6����,���� �0� ُ[�K��q���f��~�?>�\�{�^}��2
3X[&!��q��{��<�X��� e��Y�sX'	p���1��Wm姵$���V3'� ��_� ����>�d�F;��I��,��(�.ʬ��?([>TmU�M�5��t�'��v��@w�׀���~�aXM�����=x��\"�*�Q���!`|c~��X$�_����]���1MI�,��8���-�=�sfS9D�~|`��@)TR��@�z=/[���@%W��� �ܞm��k��q���-v�����w2�9Zܶ��\�Z%��n�lⰵM�����9C �x��c��i����ʿ�[���.��$�,��N�g|?j��Ϙ��x�T�|�6����x�pN_��J3��F&&��\M�#Aa%^�����s��\^��2A�����j>�*���P�����%itТ��&cvg����@��u����Ⱕ�FQ����:�}1�%n�L�q�f#(�ĸ�e
liJ������?h�E1�Hi���'�m�=�`�\{~`\�0��J�e4�A��6ND��7�C��%K�$=��۟�HjMQ���R�����˂��F�).��5s}+�
;	o�IA��ןiZ6��?�W;9=Oo�[�) �&<>�AP��ՐɪD�Ob�
z�V����m[j��M�O�4��=�.!Mo�Mݣ-�q��Zne31��תL_(^��3v�8��eH�V����֏�S��"|]qo"���M���v)�Λ	gg�SDn��"�����q���k��;����	FF�u�*T��k��7��R�S`P�=6W���`��:���J�t<��#d �i�~��Æ��8�O��*�������1��4���'�0i�Q�*�X{�;W�/2tP�;�*��}ᡭ(t7kGf/W+�V1��_H�k�et>:΀�����q{����ĉ�oQitw��+�����f����?r7%jwx�{�!��rʹ7�#$@ ��nX�yR��%���w`��3�j����d�::��WVU���F	��A}}Nk��lemi�\θ��-��3�@��c`{��
����u�&�����%�:�f���A�����M����Snw�x�Փlv̅�V��پ�[�� Y�RX���8��g����îd�Y�/<���1fR��Ɯi���Z:�l��=Җ��ғe+�g����x�7�A`��VMۙ�2C�+C�L!e�����!�;2�;�3_�Y}޽I��4�x��"�sٸPח��))�:5bN�@�iF�1�[wb�u��E�{3^��`���vJ{���IH�$Vg�����t[�
�#�����I:gl$w6uS�̻�5���꾾$]���u�;EC&�6��Q�N�jM�t�6��2��W�Ŏ}�F�����d��捦����ٛ�e���	m`S��n��J��%r	Խh�D�(5{V�i �%�+�a~g�	�i���;����9dl�+ǥ�URLH��.b���U|�6Ԇ��e�:={����*9�/���"'%
��,X�.V ��'�g�s�6�I��˙���`Iԍg�7�(��%-����.J4�� `���͡��n"Ij������t-G�f3[�v#L5L�æ���)����l����E������8Z��oˏ�dՏ:�O����4��o�\�z�>.���w�WRB_�����6-;'B%�����-5������t|Nճ� !�s�`�"8.�_�UνP^����M9<����"��,Ki�s-r�9PZZ@�`�Y���"L��e~#,Z>ؿ�9�AJ�
�5�w�σ@lT���۠bDU�|1Yԫ�g�_�*vp:���K��A�k,WA 
n��GT�!���eu�k:i��; .!�t���h�V����g�N\?g.�+`6lP�h���Ϲ{XX}5��Mt��b�wQU��hC�����c���5�L��}���i�QND��=���{}�ddf[�w݂껡�qWJz)�VRn#d�"���R�H���l�B�5Ks��L"�??��qy����z�A�z}��1�Z#�3�=�?؇"����Q	W��t�GBk�Z�JU���hE̥����wB�#��Z[�Є�D�
����ѧ'��v��ɂ~�J�I '��p�G=�o��hV�	��[�?�7'�rZ�
ݹ�I�1z���F�c� ��k9Ì��;�;9	� �c�o��<iA��A�����&����h��>|��Y�D��Z�p���,��V��y��5W��x��S�{���j�7�����5JĥuN��h�\��E�����u�n�^p>�[h��~�����'��+ [봱�"m���Dg�������F��Pn�ϊ� 
���S�jLS#��
hջV̹�}�/���X�=�F;M7Q낤��r3aJ��A�]�vwkSw��Β֜Y�k<#�Jfy��@$?���_vnu�D�h�p .ѪF����F��vb�֑����=��x���1�/<���$�^g���Y��<�܃��s=��S=.9��!��(1�[�D�vJE� ��-k���~���;U6����m:0���r�Q�b�t�5���qϊ&��%C'a|zg�F��OFe2#=�K�� b�[�eU�3ˌ��G�F��y�
�F+ɠ�o�0+P�:�YZ�k���1I�͗z"�����U�Rs�.�w�&](��p�'�d;:���z�k�����[�Z�X��F���I�)��8;d�Di�W�K���5���`�#��q��lLW����A��d4��$��C��G��a3PM�4�Y$>dxː��5Ƈ�	o���K��-�+Bigk8�2�b��"m�_���:�h|1�8����c�t'gQ�m�n�X/�T�cԛL9��لiF-��c��|]$��SP/����}�r��t��?u�v��:�	�G�2��Tui��{��_|�"cf,��6�\}LvFr�l��j�������j�|\��	�א��{U�h���-�����}�ý�o�99z�������}�<��FT{��s�
�"�n��\�*P��jL#��@�޶��T�,�z����ӥ�oX�
�~���sw{Rz�gd[�j!��x��i���i�����s����Xs(i5�y�dij0ە�Y��;@�T�H>s��Y����N!�TƔ���B�/�N��O��g]LʈL����gk,S�S��w5*vd��,.��Оm>��bb`����us0������(=;K�b�Ls����$q�A]��c�ƄR� 5oL���r�0G+4�R,��n��Z����W��D�Q���CD�,��x.ޚ�C��(�R[�9O�}t�T�^�\ fx �$�;�6�/G��T�43����cvKӼ8pV��29����4ܓ_y\��d����/��UzX�%~2j>'.D�N����'��u�m����@TPgU�H����Ќ����V�N�-�B�-�g��g��ݳ�u8�&\���`���,�> ֲ���*X�Ҡ�M7�ذ"�o�5��E5�U�RQe�Vy�i���%��ʾ��������s9���� 8�-�^=�(��Or~�[
ɼ��j6�������yh�n����e�e�ڹ���[|�	�NK��rq,��ݮ��.���UD#���~�A��!�7ۃ�^K���N3�(�Qu�B�MZ���Ha��=���H0&	B$��A���ꃯҧ~��!�=�Ģ5�8���p�3fA�Dm>'�~px;�h2�D_&��|C_�wPSE N���S=�M�����k)�/�9k5fH���g�T����S�}R;�Av5wPI��~>���+��K�a���k��������̮�׽��ڌ=����d�2��g0�q���{��s���-�k�=�xC�#%k��YעB��/x�F�?�(�k�s�/v�t�	|���J�>����o��)I~5����hxGK׏>?y��nM+��U_�y-t%�S��]�;��a�q}̬�L�}�����r��K'u�Yݛ.�?��(���;��!ǣ�q���[��7�K>�C��iIK�KP�F��(>#��5"�Gn`SG�
R.�6�8��a�J�S���Jpr8����/>���%�P42)�$(�_�r���Ԕ>�Жin��	{�X9*�0We�E/��7�����B��pk6@�2����;Ƙj�2i:��ß�_���WXڦ�'zAX��9��B�����]Γ�S�U ���tqf"���a�6�H����g3���$�)�I9���Nn~�l�W�Z�uNrP�k��,�$�; �e�ӑ�{�^�?��Ȯ ���2�'��w�N�U��+���B��X6C�{��P�]c�8�����/U�7˄�ļ�D_BA�:ځp�����e�%N�Qp��˒��ȉ#`��s8��+����A�uXY5�)��8FϚݽ]ۊ�j囅��Ď77��!�M�����k���@)v�ų	���=}2�Ů���M��;o#v�e�O����n����f�(tPV㇢,����G~��Ơ*��D�͚֩�G�`�o���� BN]��)z��=�tl�~��p�A�[xg���W�ò��Oj2�j.l�7ۓ�KM�5�E���ř��Zo�޼ځ^����	oޟB���L�R��--�����ϳJ��j���0�VB�W6���Qn?Vo�r�q�c���,��)bo��y&G��~Ý�O��er���7���q�v}.I<��YA^�L�Ĵ����#$H�$��4���#?8��;�9m�����v�	}%�v��S���-ƙ��㺌 "��Bd<��9z�	�~/��(�]����(��Ru_Z�Zhg�^��׿/=|���!)ؘ�(����.eJ1U$�U�`}���K��ɩ=��jϪ��߆2�`<�Ť����s
&�O�V%!}���TNӯT#�>���ެ!n��]�- %������q+��5+�C� ��0z���Y|BrTM}�u9�y�Y�mS�qgLO��ױˡ�u9p5�SMby���c��o@����-=��D3S���ꏞb�)��ܠ�K�r�ŌrS5��,��I��d80b( y���Y�\�[���~�bf]ig\���F���8F�a��
�Ц#��gV_߳�É�*�� ��yD�� �p��ڡ�A�\%��G*��|�;���.�V�|.ߎ�V�'�Į~ͣJP���4u-��*�JZ�&ݤ6�	���e�q����0����8��+lZ�Os!��1��Ssx�['O$��������QD`ͻJk�0��������юW�����ĹaO�a����IO�ޡ!��Wl��w�'Kr�A�������޼���v:��}�7ҿ�B?���$�5,��TЋSq�l=�r�{V ;���d�k�gTb��m�t�\W���H2�9T���	�e����)�� ����3�v93�T�o:�M4X1���(��+���Ay%�T�KꋄK�0��}������Gb>��8|�b�;��?6���j"掵w�}���;��,�jo�`�ǐ��p�i�`�q����|k�=[>��ZS(w5��db��5��v/S�84tv�B&h$�
��vw�4�~�pT�D��X;`��N~߀��i��6)����"{N.1&�	�U���!�5�g���tt�#q)�"�-3�V��]�)�r}�C�s�|N�����I]%��']�[�d4/a<t�~<+y�GGzU;�y�����[XjM7,�M�]�b��j8��:���ڨ[�{+K6?"��k�C��:şB���>������@�c���RF�L	.�����?,�r�-�q�v
��O����V'ɱ9k�C;�ݒο۟�M&���>��E	��;��C��-E�����O������%�<����c;����>A���Ʌ\/g4A���+/����Re�`*ĺQ���̩�G��`5<�\��O�W�=�2�?�T������Z��w��*[L�*
��K���޽\�f�m�}��η�j(Fe�r�/4�F��>��a��Fu䕂��$z J,��5!ܢ��S������6E$w�	o������BR��gA���t�?��&�Kp]EsR��h�����M61E��3�D�,]nn�e�lw	���j�C�#�� �)ҷu�0wy��@�.�H�R���2��@exHE�$��h��#�n�o�/	�9�dw��?�� >���L�몬9��s��ˈ�j	WLΜ'x�*Pϴ�+��9q/��ŉ��T��*��܀Ж�&�7���3���U�2J�o6�u���J7y�����9&˽�Be`�x�Z ��^�q�'	����|�w>؉�D�	߭�r2f
u���vVJ���ȑ{��:+��%��~&x�{��W�b���x�R���WW��:����6�M���n�v��h�EI��RZ���Zvsn�JXk�?>�����\�<�cW.�#�Z};���r�Z�����B:A��i��y�o�� o��nHC9�Q�h�f�X�nn�Ό5��?[8Y跥�U�I��8���e�R�dv��>�K˰�`��S�;C3����|۽T�̋�+�'�L��c��X��@��]��&��3%��������\��fUˌ}|\}_�'��>���e�ڻ�R�dQ�@5"拁�}}��x�E�粨�
q�LO� p�I�Wu�bGa&'`�K���p��"+�rUw�q����j�H6;�����,`����%�V���D_�`C�3ϞW'[m�>;?]/�����q�/ή�ң��eD��]�Vx?�^�3"����Q�@,G���-^�����;Ȓ�JaW>!N���\�F=�`32�z�F�5�l(i�$�u!��rb������h+��͟��C���k�#���3�'z����B�z�ĩ�$���-%�7�G7il`fek��Y}�+z0�����,����N�hWd[��!����&a��w�+8΋=5�=�3OTUCQϻ�\�WX�(�ì�LV9��WV�xʘ�3��������;�򔌩"j�Ȼ]�8o/�g!P�z?v�1(`��!N�Rt�?Cػ���+���|�֞�.ľ��:�/
$�e�����x��-��|W�5n�\ݝ]�>|1�u�T �-1}�s��,f��c��omo���/�y��e
N�a��}D�M���-�����d!������C�Ϻk���K�ngҨe9���ܜ}+��rxMD�r@�]�yƸ"҇��sYB�:ar"=H�X��\n�ώ�aQ�s��R�C�/@ڐj��n��캺H�(�f�E ��M��,�H<�O��?�F��Z��(&�˧�7��OR�i'h9��p&(��䛴�{��RB��)]WO��lVG�㥕��E �+��1�nȯ�;\;˕�Nb[����#mRDg�IV�j���_$���O�fԝ�c�.b���9����@����w綗�%e��6aF;�m�?[�U���^O�����E ��FW[�#�|�������:RA>)��'�;���)Q�$O,3� $)#��'8����Gq�k0Y�J��U�ė�J��Jү�}/?K����Xh�́]��^�!�_Z�DY��E�4Sޱ�0�P���3����ט�զ��,�8��R�S��p�n3~]���� �����]	$���Ȉau���ܚ�-H�>
)s8�l��Q]�:0��h�*��-�*U>���~9�n�Ӫ\�=�r�G`Y�C^�g6]񶡂�.ؿQ�d�w����"B�;Y�
�	�>�f���yۧ_؉%Ԫ�Qt�5A���e/C�~�vQ�����3-���J	ŒW���⛰�[֊>0IW����݉ah��&#sdi�[�(C��xI3���vw���o7K�J���j\��y,Si�(���*É���]ı�i	�Y�Qb� ��m-y����A+Y`=�Wh��<��z p*L ��t����u���z��9;{m_�L�֞7e�)�N��A$a%7��P�-��a�>䆯�R�ϊ�.��c�oհ��V�i���/$
Z�<�X�u_�6dc�dRBP�����*�<��K;����s��qOmCm�n�"��4<�V{�R"��թdM7I�¢�>�\�6��7g�r!�",Gk��\�����G|���EL��P\?�zT)q	ya�D��N�J����.Z9�ҫ&S�\(������1I2�^��BǮ��՘x���9/�����Fbi����Ţ�=���qYۧC�_�E������5��_�c"#�h{��z��2�AU�޴n�7��!���]����4a�w�Md�Vʹ4r�O�%R˗�jȚS�c)+�"e㈷�*���ͼ�C�>t�x%\U�����(�����1�L�N�{��%o��=6u��R-�i�D�P�ū���Ţ~T��)�m�/��f� N���7DѷRJOT�&]7��6Þ5�7C��-|� ��G��,V�}�0�F��X�K�C
j�T��[��O,{�)��Kv��G����2��q�%�}�{˰��yyܥ��a� �@��w7�`�@.����,Dq݈N K�Phȴ��&�y{3���Z��קHΜ~�AK�|U����_
�������Ts=It���M��u15�B��'f]�%o�>&�)�Ų�Ɇ�M����K)\V#�hN*���������ަЙ�.*�wn�J:�#1�}�{Ux`��yu�~'�y�T2�Z��&��k�f�2��ܶ���'��]�	}��n)�)�|Rf@+����`��E�_�����G���d�g��m ��*-ų�c[�DMu �q~zo�tqa'�"|=����{O䴝f����&i�e��G)���-V[f����r�1�����յ�`�A�l��m,מ��G��/�1k����Hi��ϟ,i�M	f����˂�R���/��c�;:V�d��6pz�J3f�6y�a��(p��j������p3���̷�t�I��pðu1�eX�����VO{����!b�� 2lMŝă�B� 0�X]R��6[G�!Zw��^ ��~:����g��{^�4����X|��q���P|�I���C�]jȶ�p��ӁG!���8��:e�c����XH�p�	��a!g��F�fq�n��#`_\��.#�~"o�:@S%k3��+��B�q�6Gz�nG?J�0�z�p��i}0Bp�)6�fjC�Ӷ�殐q� !��f��k��5��g��-�N��x����#}IW< ����.�w���S�Nϧr[��@�Êv�\��)Ǯ���|ˡA��=w����e�`�����*d���:�їc*e�9-qA.�mH-!�Z5^8 4��+?��N�*�C�^d�e��g���DΟF#_H�&�<�Ԩ�J=7���k�  -����%k�$J�%y�~>�,ڱ��R�I�j��َ������M]P�ז�� �ă a���,��m��t�)'��X�egv�����j�Z5�p�Ko��[;�w`�j���I�g��m����Nv:F}M5n,����:X�N������1�/���Բv�t{�F����ᷚ�����З���ё*�j��m��Z��k_�\���CD6yH|�?��8j(�,�W�ڸST�3�A�H��H @�E�Xr`QV
|�:0SGgY�,ډƍ��@�Y�,�x6�t�B\%�b�TzO����	 O�/G����(��;�g�l�zE��2��e2`T}`*AŬ.�X�mIb��~����L��/b{��2�m��tf����	��)���X͕��+�
�����~<��r�L�˦�5���_�6�	���U(s݀H��"�bO]a���m*%EP�S���n�s4�U��3�d\�ɼ�Bv����|�N�/Ӏ��#��?�k.� �/�#hiU��"���:ri;F"w$�H�O�Mp�_E.��f��<~^X�#��O�idC�O�[�~X��<��H�o"�X1�����"��O�q�Y1�7��h±�G���88`qZ~�c<^�myD܋�N����r�+��S�j�M���T��߈���L�Z�*%�\f5��24�Uyƀ���)A�����n5�(����p�gn
ix��ˢ�b��$��!�����1U]���ᜥ�s�"���N�ۧ�[o𐜾&��`�͛׼ȸ=�$.96c��J������GSA��snU��l)d�vP볊�{>!�<}5^�.��:����Ȋ��F�PG���.'��Hʚ��⺣1�����~ע�����Ag嶲PT$�����ɰd/���@���8:cxZ��).YI��D&�M佗��i��1R9АHbh���-�pxU�]�i�!��ԟ��RG�v4��xKr�}�|¬#p/� XWr�n��?����Q��$<�����?�@��Ě3�S�x��!j��R}Rd]M��Ne W����q��Pp�.�NX9�-���jh�����3� ��"���$�����1a#�Q����7���)��PzG��qT"��ڷ^�&?�?
F��(F7��v�?�uJ,P��3QЮo%_HKy#I�.����LS�Y,m�$������~�_�W��>3������ ���c!�d��Y֪yo�^����j&��_�lM�5����N]W��u��#���895�ԏy	*En�ǁ�Չ;�I��5li9S('�|h0;-X����.kr�UrP=����a9o��yD����v%��%���$�([('t%x�'����Ip>r� �.S��rae>�@��{ZQ�>���;��)�鬎�D�gs9���������O�ӓ�O����]�~��&_v!�Ѳ���#ž��גPm���wD�w�T��h���t�ݡ���1�"�L�)�u���q��y����j���/�Aّ�ȷ�t�[gƆ�y�qt�����R��鹌"9����$c�k�;J8�R���tB}[�c6t+�Vʪ���>C&��h�mI�3�%�ߑe�u="�?H3U]Ț�z|�A�{��/�[�QV��q���������,��k���j�t���JT'�� �'6ܠ�MJs*-�j��
��H���'V��U�4���i�V�
�a��R��y����0x�q@ܮ�=����	n\�r�Z����N�]���#��"���dE�T�[-���s�^4<0·��)QBU��B*WgÊ�,�a���:���&����F�C��0]���Gx�`�C����(�i�3��{�I��m�*�T���鎺;7�.sX��`����;&�׫5�!xR�����	�n��M��?� j�G嫜?���8���R)��d��2Y�)<���E��ũoSI��*����W4���{D�t�zxZ۪��M{F�ff���ـ����		�3��&���D��?&�S�	o���]�hC���VOs�(�	j��:
���S�ǌPO� ~q[)�����xeyN�8���jo�]5| �"N����f��R�!�<�v��XZ4��u�~�p�uŜD\�'�����q�1���u�Q�,�5�
}����1�<������b���n��o�����⪎�@���-U�����z��1�h��S��AZ�F�������6��Q8gi�p�`m��x7��K'Ox1zQjYAGFC5k�U�p�P�C6hπ9� $gb��O%�$�}���/2V0#��q�S�-�=X�<�b�6�Ψ<�)�
HL�U��ܢ�;�M2� :��:�$������^�S���{���q��+�5��u�g�V���!{z��p`��7��@�zA�U����q�����ȊJX��87�A��҃=�]7s����4���AO�.�ѿ`}�ݼ�.�_����s3�Q��}�Pų�W4z�2�L�&�S�W���%x���=��Ѱ3����M���J,,�9�K�6�����D�8҉&�R��{�jnw���팷U"��Q�^[�Pb@G�p�-�3k�;b���U<����d�V��[�+AX*��G ����ٴ��z�;Y���݇�So�~�Pq��,����r�Fѻ��������.Qq���4�6��#��_}i ���j�z ~״�7qd[���t5���+�h	��t:wo��~.�EM�Q���O9�oT~��sw�g�Y� ��S^5��b �]S69�l
].>��g�ԌM��#�qO�N�*��nȲ)�t*�@�~Qb�¿;�hX�;�$�5�5������F�e[8B��'ͼ�ڃޝ�0|�S��<q�=�q��T�J����?�x���~��W��s��O^���D,���)f��}
���b�m�Rr����b�gbx��nI��;O��Y�a��FC��l��
x7c�����	a�~��u�#�;����bv,�t\#䶁m�Jʢ
��}-���H\�$�.�glBe�L2b�I�b�B%C�)hg%�0��I��A_3J���a���>ksjN�1}��(�?�A��6��uI���|@�?uJ��<f�	���Ù>4x��1��1�=�Γ'Qyp��t%�"%5�1�fK!�t?�X �ޱ�I��0��b�M�(����% �Ԇ�/�N��3�e<��p���3<���X���'��'��`�79N޽<��bn]���-����7x�*]�\eEB6Q,�9L�b�L;��~
�E�0����Z��t6f��������<�a:��p��-V���󅗩�q��!g����N7��eq*�,!幗���9��y����%�C��S�������hN��ݭL�92�7"m�������	�E!te�5�Kb��N1~�`p=$&h��hB~Ct�4ʷ>��,����X�d�݂�9{l)�_ӓM�Zyz�U���V1�Hգ�a5[�&)������e�H[��,�Y�U�A,���/B3�0%�C�#g�A��$��������&�����#.u�@��G	Y^���t����6g�� ��f~�c�&�����2�Ʀ����q�#��VY��� 0���pt��<�t���"�r<0ϖ͘��8���'Р-{6��쨍T0�0�o-?O�zɁ���V����@�D��sYz^��%ʎϹr����� ��>[ݓ��W�ҌZSc��@/ �m�ʴw��r=A�5�?��Ӌ&��*��T���q���	�����@M' `}��:	�2 B��-`Qߔ��zt�A�^.�7�C=�t��a���r"������V�ᆟg̔|S.�0h0x`;�^�.��K!]!}�w#�̷�_�c1���x�쀺�DG�껽d�W�׷�~�Co���4_c��e��b�W���T����
=gA��3����r��+x�A�ie� ?�1Hk��I$A���uԒ��$(�cuj"zn��z��[�$ȱcȾ1u-1ؑ�����(��P`�f:d=`��Z5�O�`;�pW)���?�rHa�+�u���4*_���@�!P.�&UXNC���m��4X�����IM����ˏ���%]i;���>�t��qK]Ө�#�F���_kƞ��C�y�_�;�J���<����
�\{�t��N����i��uI����B/�ja#��ly֜D���T2;;}��z���b�&*֝��ב�,����]��yrEU�1��s 3������n���㜅�D��&}.#�\`�eA?���H��(�����b���� A�F��TeM�l-*�� �l@S���#c���pEk�a�n���E�ҲN����@F㥼�t}���]�0��󦗷�C�x�rY�1&�t����z�߷��Z��w��@�us�v.�r�/�p�z����~/J?Z�6�ǜ��kCsFW��cq+Cn�=B玥nJ���R��u&^Kl�̲��1nڻ���K���ώ9~���I�Z�/�� %_�Saj�W���Q�wF�'���:�p1���`��V��@v���`�5�
5�,v�&۟��w�<Pxn�R����N�G9��
��s1�(��5�{� ���y0���������3�b���<�3��g__�|�mE?�F���yjt�;���t3�����nwG�{��EP��쨅_��了e�-��3���k�] 380�D\Ы�	�4ԭ����=�{B�V�+� �c����92��pp�?'��#��pE`Tt����(��	늿j��e(k�#��@��3Z]L�? ���A&�	��B���9NIh9��������,���MWD���zߎGD��U����8C���U]n�޸=�o����|u˅��\��/L#=�>���v�u��M\?FG��b��[��O4���d�Q�@k_z��S,�P��{���O��,l[�$��<���O��w>����E��۫-�B6�~�D�%��-ݤ,��ɵ�2�R_�+�I+~�	����LaQ:�{�N_�or��|��X���Kju��q�`>.7��(B���s�(�HZ3ɚ�!�;�s7�?�?�;�r ���z���a�ȉso9�}(�<B�[�IPv#`��<kZ_Ծ�pn�Oτ��k����2����� v���]�oQ9v��S�y���R�s��~�q���̢���}3�n��[�p��-r��*�E��;����>�7��9Z��0S���n@��{����r#�Zt�21�`��0Ԑ�m=R�1��w)H���]s�X�P����VE�;��H^�����|������A���_""�V�1LxS�.Wv{�AD��0i�L|�ߙ4o�e�z�4#u��$�%�}�J�	��l�f|�̵@�{���!+���w��.XT�ձ�+��S�E>�ZZ���"�AZ�>��pwny��*ݲ�Q!>z���>B<��t�*]\	�Y����"���M����[aG��t�����1ul69�v&�`��#3�"�$����k�7\��
���7O����H�T����{�	t��S	w`X��(�(H�#w���'�CП]a�K����$�J*cϝ{Lt�a���E}5�X��g����\���xT����6t�zW�m`���X,�cϐ �JN���s�I?�O������ZB}�c�x-~��\؝���O�A���Ն���2`��.{��LH���:��r�>�R�MV�t36f��p��+��z<>�ˠ��g�/7Y�� 8��W�&)"c���i4>��QcٸĈ1Ļ�B>�]	8	YZ*Ά�q��}A���u��{��ruu9Ȼ� U�K��9�)4��kKD �B�0ww��}j U%e�tb���i�qy��g��i����ߠ�
mǣ�[��]�|ŒrB������E@"�8��T�?��&T͟��>R6}�:)gFP�v��ŗ��߷�ɷ{�!9<d8�ſ�i��(�L���aqʗcB�D�P1E<�D[la��q��".�sA ��\�̍��U� �K ®��@�u�Y��~}���AXд����"n���=�p��	����m�I�����K9b�
�U +燫BdH�U=h�%�0.�0�3����.����߸Rq&������a��Uz� EFQG�����fW):�F��s9���.�%15UdQF��fv#R�3(�~��Vq������{��T�q	���6��9ѿ3�`��%c~�˘9��f%],�U���2'�I�j�����t�*Q�I���F1���_yX��묶?�� %����Iy��f��]�����wW!'���n�s�\ޟɤ:��c�y�I}LP�`�ԑ7�9��7�朱=�}��vѢ���	���*v��ԍ�,�q]଴��]�Z����e�n7:(���i���|h�k���)�z�9��8��gV�N2ڭ�������CdR���a�U�x���K�XeJH'��������]�]��D�mg�E�,�>Cnl(�3���A��"�9�Z(�@a�O�d�Z�y[�B���Y��ݟ�N�$���/�I��L���W�zA<��G��&H)�B�U����X��w������¹2���3pZH~Y�L��ї��;�|>��=n��}Av��vߟx�O�&�V<Bh��S�NU 8V��A}DY�B�s�h�J-L��;	l���ҕ��ջ���j�H���1�*3E�}�Ը��[��[���^��;�LC�#)Ԟ������3ڰc=/@X$���`���5�$>���_�Ä�v�/4��I�@��&0j����.���L�2c#A���c�ȧh��������!�����ג}��7f��	^D�����������C��P��zK>]����ژv�� .[�?��*��>��z=��t��/|:�����R��+58X�SG"x��S�/V�*>�M�Jw"DQ<���8����Q"� ��9�h�RB3nyC#�Er��� x�*���f%ρF[j�p�zR��[��%���y�b;�/��=YE�ضݍ�����EI�HV�YH��O��]� M����ʱ�������)���
{�jҧ���5�)�	�/�#�B_sQ�Ά��?@�b�f��-�7 �_S:��c3�� �^��D{�?��b��g��K�8B�/����\PmD�x��.6�r_���ե�H�d�A�g�+-a����3P�#ےIY�X�pd��R�B�%��GSšG�M�E��!�*b��:g'�
ʮ��@"��G[%�$b�����/-	{�H(<cM�&���~9d[5t1V���� |�U�&Mv�i&�w[���!R�U8��*�Ϩh�("��CCf��m7�Mt�vYT��_���r���Bu�!iն�L8 
w^tZ���W;�~�T�����֔o�6�9���C<χvU�q���X�yu�`���ȟ���rܩr@��C��̹-�bf�X�P��u�A��B�`�U��o��ߨ�����*�`sX@)��G�L�l �)|4�ji�'�ʤN���:�k��{(L������7�G4�I�tϙ�B�a�:Ða��Z\�K�v�<q�z�N� ,����8`k�m�.H׹'��s��!�n��x����3��Y_i���o:`�ߘ� z�e��񺉌������I�q|�Kө(glԜ����V�jѾug'L�ݳ���Q��8FU2@�30.�?1��Һ����ڕ�0���k}�Ņ���3���<��_@8�� 95M��p�`���(��ͧ�HÇ1_�9VC���R@���*�$9$�$xD�d�K�@�.hR��"c�@T )o�6%�c_�z�B���W�e�{��[�*��Y�����+��فF뽺��a)�qr�8�G��!3p��3�jOM�"�������0e�Fk�RK�Ka�k}�^�������������X#k��SW=3��a@�8�H}�#�fʃӻ܅P��;���"�Óϊ{z9�aW�=(�H�5͖�dsUh��%o0��F�*�C�D%�S�џ`��ȟ8S���we�N��Go]V֍��R�����s>/w3Yu�:����S�:�=���~�}��  I��� 9�̑�M���Uy���H�p���򏕗�J��(�p��0�t���!��]�$ ��움�÷�vi�mF���4.��z~>Z�x��k��+6C�y��NΓ�M!�
,�pj��ny0D.���,~�}�E���^�~Dؓ�j�rˮ��k�}X�(�o�5H�%zR�Z��ohG,�&�����U�zIK`�Y�x�ɐD�����������Yv�k�y0�ó]2��+U�]�\ �oe'�$��:���A������yſ^�V�^lEn������ba��^�y�s��*U�fsC�Pe[sW|�U�1��!S���z���j���;��%��ҟr����ᶳ�,��li�?Q'���^���L�	ع7J��b���2g���a_�+�B��e���+�}�界H�a0B�Z��O7�b.ݘ*�b��RB��- �(����Hm|�����]�O�5y0���z�p_���I�h��z�9��h�'A���5�{�<�K_Z�F��Y,����p[7���KI/h*���x��i2��@�)q�4dh�4���Q����K�n}��`�k(��]�e*{��x
��+k��IFp�~�(J���$M��cL2����0(���T��"�1�W+n�c�(�}���Pr(���l���Z+�&�+��ő:���[�-�����ȡ��m�w9����o�����OtK��<a[g�#0Z��#C��Ӟ.�����Bm?�n��,��vA���#�x2�y���o��b�j�Q��3�]I��cgy���^h�R_͵����5���yI䡆`���'��i6I}Wl������ ��[�Ŋ�I�S�X۟���]�����'gĠ+����b���tͬW�|Da��z�Rٗe�8C�Q�R���zB镰<����i��g��H��3�`��:���!�2��)fegE��P>���o�В\��F,�8X�'к��j#H�*�#�Ơ��|�l�=j����p���
�.��ƌ∝��}�>��(|����y�#���\��*EΓ��/����J���,�7���`��i*���o���/�Ƈ�?۹vu�|ᨢ<dΠ����4��0?�ՍQA!+��H��>(�ٽe��y-й���]�d�
�����<��Z8Ӏ�4��*\�C@�c�G��h���P˫�K��2m�T�y��PZ�ض�[��O�3.
$�3 �,&o=���t�d֏\nB��D��S�zd�!�8-^�ɪїf�=:���x��s���@�%�r��o�u5>�+ߨ����H��m��×���;�2�+��L^����-�ב~6��f �aLl{1��w�w�bp�u���ҘC9�N=d��Q�n�ߪr.��C��
��#��Jl#;����/�F�"@���� sw�ɇ��f�/<Ś�XlS�O$��*U.�o}�^�r�\Ў�����pt�&G�ߥw�h�CD����b���c�yc Ӗf"��3��`��Pu�^�]l�m8���vq��ȇ\�+4fa$!�ӓ'�)��-���/\�F_'9��O��z��b@w\��^���J睸�j���;�|HQ�:�%�z��vKb[���z��c��|;�A�n��qU3"bwn�1���έO�(0��R�JԱ3��H5ء���(��ƕ	����+��.��Z(�׷���C��4�
r�6kR(�s��Oy3����L�(�,Ѽ�9܏HW�hE�V�Da�s0����JӆD�0�E�"z�bN	�{}�	p���W��G\�G%�����D<K��0�� �jX���랅��DԄ�H��f#���,^G��� s��s57�ur����fH�=�C�~�d䋲g��`t�T�j��D[�F�����ܭ�[�i���� Ev�S�Ǩ/�����@�L��ʥi�殃���o,��Q:a�j�Q���I}��b��`��0CX{h�;�'ɏ��`6�~2}���oQ�0����v�.N�U\5�O#�L�U�k�_���tb��!��UQͩ{�E�0��n�**��s��"�����&���kA�Rm���P!����G��|�Y�`Q����|�i5Ʈulu�F�7OeF9ν�V�w�����z��Y��J��%O�f�����(����ͪLjY�.qGeӧL��bW:��j=a���+��tC�_��$��~h���яd(*[��_�	�X��L ��@o?��C��Ii����|��?�.�B���(٠�Y�]�����&�0f��ݬbN67�%���p�|�٘k�\YAf��诅�3[�C��m�dp�	�WXk�V�璄���{~��e 7�����><�/k��z�U�A��|��ɾ�G~ǚ��� ������LJ5����߿��`��+�b�8m�L�����2u=��ɘ��N\{��}�z\�-[D�����8?��eN��<.6o��'s���� �Xr��g�y�; h���.NC��j�v�u$�Qà��	�1�+X��{rE�Xu��-ʝ��MW�Y(�^ҥ�l!��L�f��"[������Qɮպ�L��$�Md��}�������(pV4�=���0�3u�v>F����d�?���Kx(>�R'W�]w�t9N�q��'��u��@�|BD`�L��*CD���g4��['��D9�oa�.�M�����?�Q���d�@���Un�r��5%�t��Va� S�;F���@h�殏Q�K���`]����In4�N`%Kj����ch��q��'�nt�g��W�҃����F�p'�_6Q�J+�t�jETB�;\����,IE ��%�g=�{���%����-�Aj��Z��&4�+���;��ٰ��GB�?�[�J�r����.��������M���+��*k�b��i4��]>4dD�1m?e��2#=���h���a@37H�!��&D<ngIg>�F����M�wU~�)$țf��]Z��Βm�
D�;�9ZqI�jw����#�S�h��
X�M�;�҂�D�Jۗ���}+�h;�d�ꂬ���|��j��,�VU���Qk&�{��W����<���"��
�D�[xTv3`��2�,L9*p�q?؛~Z�|�W�gR�u�-��Шym���E��E�g�D{'hC�	z_�܌�MؒozX�r�,�n�ި���;3d���;�A�֒gd�'rtLY��rU��?�z��1lc~�	k��~4��O�WDֶ�eڞ�~�~�a�i�@�U�����\6)P޻��ui�U��I�g���[�$�D&��?{��,-}��X>��R������#�F4~��nE�;؊ƺ�R2^�1�/6���kGPK�[���w�Dc"�����"���CR]<y�K��-�ZQ����34���x�)���a6�A�jKxG;އb�h�F�i������{�xR/��x�7�����(��W#��wn�ʝ�r7)����Eг*��,;�W(}�~Ü�C�r�<;���6�����Y�	uo�̹B=��f:b(r�u�).-y	k��[�i�/P�J���&A��K���6����I����"*l��K�p�۾(�j*}E!o�p�4�L�y`�����1!��P6�^����P�Yc��z��au�5��!�i�jq�DvJv��W0Z�{�x�]O���'��)�}���2��WAG��X�a��[�NA+w�oOF�m���%m'�<��[_���&p��1y��qG�--�U��l��ݰ4��R�-��)�E�8&�UrŻZ����(�e��(�
�4�<׿c���m���hNe�L$����mBvW�{��ᙚ�I�h�M�g�N�C����Vv��f�=>wOzW͜��򋏊����� �������0��D���o)w��`̡C:���ax˦ռĠ�s����V�/��k�ĸ�N��/ׇw�|��YED�����/Y�v�S(m �>/�M`$[1�����h�~}4�������O9ME�����a��p�SN����|��2&�o��ԩ�>��g�g���[�}�Կ(����J_{YH$��0D��+}2 4Ȧ�jI�(S}o����-�]�4��`�nW/G�~2:�ßƥ�=��D���d�$�˾�6$Ѽc��tT�V��4�����0�CY��W>��43m��&�Z�̽��N�*[;V���N��9�dʼG��4�2���g�\*�~
l\?�#�F�F���[�T@i�����J9+g�nXAv�\�B�V]�m�2Z��G\sS�>�~�}1��� "xfZ�-630���������I�_c��p�ں��5ׂ|c�[H��JU}i�0$3Vv��~qp��J����j����\��U\���&�L����%�H�\�`��l�ݿ�@�����2ƵL�B"��.�"�0IS���&,�e���Z��#��1��L�u?�j<`���z״9*�J+���+&��I��l?
[���wQ�,'�}�m
Hy��{� ���}���h�\�T���h(���`8h/,Q�'� ?�ل�;�g�N��n:����t�좸�N,d����7�B7��h�������_,tmo>��=D�U�6V$7�aN�g쓅�FSȳ�`�!��[u��)HV�`��s��G;Z�|;���X��d]�mHO~�j�pR:�
�����
;�*P7�=�����0�M���3pݶ��oTg_�lܿx �i�7L ����i�n�D)e»w(��o3��pA�t�V;siؠ¤�W|x�a����1z�E �Ozy�roAG����Xx�����`4*�H��|y�.�L,�Wsm�tc���ѧ�Ů���d>_��y����㈧��0�#b�s�Y���H��L-E,�V�&1�Lԣ��R|T{Y�}A��Ze6UyczK�ʑ���',��9i���(.R�e)j��5��Z���8KQ��Mq���CU�]Pxb1T^������#R�6٪Z���B���
�R4���=ylr��t���Mf�G�T&�Q̄~(�2B1?�-���UAv�^0�w�\�����j�:����f��K_n�*�`/�¤�1�_ؓl�N�7��!fc룖�!��o����a3��ǀ�ԏԝF���-�9�g��xJ� ??t�zA�g��65�c����Li�H��J�+�����M�5Z�#��{����U�d���~z���qYo�_��'�U�����uG��0�5v�,�	H�(�C��ɔK���]��g�)HA�V
D;b���&"8e<� =��@5wܰ���KXl|p�(���C�9U��1Ճ���w)p)_�xM�`Ma0��G������I�_�mI2U�盡R�N�i�䩀� "_l҂#i�m�d`��_�&>���M%������xz����h�b��60�}�����^^2�q�s~b�������@�"��i�d�1t��$�����/n��9��j�%����kɽo}�V�!H�o\�t��8
n�N4���˝=2N���$ ��V�2<@�lAB�t����n�Ӥ���i��)�]��ՖK���>�l�g�]���EI����n�e�PԒw�����W�� �u|���j'b̹�"?��X~2��Dh}�i|������V��7��a���MG��0J#^�	ע�F\�,n������	v1[�I�$�2�-P/s��\�f��,�ܧ������C�w_�?�9�*�?Vs�#P|���Q�g��C,���R�����
�hh�e,��g��������HH�|�aIa�Pn3u	��Aa��TԵ�<˿�@/�i���.n�I���J��IP��v������)̅o�{S�D%X"޾_񌙺�-�]�Pj=�_��L��i˛^.:���71�B�*�#T�ս�r3����'������M��y[�wNi��>�a�J���Dz�i`�?�4Vn
�ބ~up����K�|�9R'�U�`�G�7T��q�CZ{���s�̋$%�?+8w؜,��r;7��S�(Dv���g�X4S	B�^)9� ���n!��H�Wn�$`�Ъ���������*sNg4�`pa.�3@��9�~�r���$�����4�g�7p��z���{�,z7A ��У�r�5b���W��*��W�Xm�I�J�].���`�hF-m*H!�%JD��du��seE_��-yz���
��m��L"�2�<�l�'d���$�SE�ŁE��H׿	�qv���IY����Ӽjާ4D��E�>�l^�O�A���f��^	�ސ�'�j�8�na�G��:���j�g�T	=�=m�2As����@�����d�v~�l��/�~�5A���-�4ėb�1�-(�y�WZ[TV��x�d9�	9J>�$�� E�D.YP���4�͟!i����c�g��{���w%q���M�(|m��2��vڛ	�}9�9����T��e\�\�l�bvH����c�ro�9<8�̥�Ѻ�$!0�DLnz�@�>�J<�[���`,Ԧ/�p
jc�GL�W��R�h��,<��)�L��!Ə73ӝ�Pl�RU#m9�B�k���sEj;� 	Q)�8�5W����)��W�[�sx�_+=�#������ .��/s�:�T[�JC%��/��u.�E���g��x^`�X�N��1����ϴ>�K�3Mt� �`�Ɖ�
��j~��u��g|�3�X�j&I*\�r��z�A�z������@��s���n�$7�,�|�&ݫ �3�V�4���j��G��<J�fF���GXڞ0q�����GP;��s.�ٔ�	<B�[0'��9�Nl_�:�������mm񁘏FH=M��x�mD�ٌY�j�׈@$�͢�MS��m����ٝ�p�^�<�O؞����p�+��}7�
���0b��m��-����vf�-��LnL�}�`��av�����0Z�Y7�$��p�Ky��@HRjݧ��,VϪ���HJ��o�S>�F�o!���(�8��-�tz�|ǝ��o ��Y�Tɾ����"�3�<��U�"$��m�y}�\YI�(A?/f�#0q���������k�#dՔ�ɗ1+�
|}��s7H;[��!Og��{������̲�<���l�m�}M ��H�Ds���W΄|�4@��{Ǵ�J�u��靳9�#�.��X�sܦ����y=%L��&��x�:�_�G7�>������2}"�?��J8$����V�[֏Z'�L2�����Y7׻`A}���������x:�ϔ�텤�����S��U#�b�)��c`������V��u�V��ѳ�� �RHQ)�젓���&CV�ɝ�����+e�� �����4L��q��C"Á�X��',Q�� �,�ґ�W/N��x.S�(D�X��6�Ra\Wᓾ�n����୔+������F���y�Ò]1b�xdt�"˯�$�����O�.����[^�c�����<�m�Y�����}�seV!��q����ԯ<�N�6���
r����`J�����}��)�cS����k����R�����#�~��������'�P�����l/&bxK{���n��H������E���i�FZ�k�Y���^�˵�Kr+|TBK���?S{�� ��	�g�Q�r��ZV��8R���^Tj�4�i�c$��ق�G��`���)�d��q���?좍xEwӶ��]%c'����4bK̃����������0���t�� ����y��:��k�k��Q��r�KU��+(N�:W�y'~�E�<hO�=2�%�b�`��(�����OR���[y�(|@[P?$z�.Z���I��<���6k˩����oV���T��� ᷻U��ǜo2C7�e�o�x�ӧ<��@� ��z�"�D���8��U��x�
�C��#�?,E9�7�?�?�}�������e��ŕ�B��Lx�	�D^���ƾ�փCz�Ә�IQ	lB��pw]��>���ͪ�P�b=�Rn'��w��M��6;ۜ��Ohq~3�W"S��N~X������q+���5ά���(8Laϛ�� /𕬽8��=���LE�݊��	�QB���}]h�{{���уh]xk� �	E����#�DiV?�R���g[� mz��Oؓ����2�ҵi<+	c��Yj��^,$Ҵݵ{N��T[�r�@���C̞��1�݌�j��~����fd��}�?�d��tiL����c+qp� 5`~*��m�
���;`���k��魴�����dR=�O��}\�7� H��c�1��W�!��_�"��,鋿t�:��e������ /3�}����d��'44g�i>�t��F�K����A���b���p��Y�)^"#�V!��*���6i�Mp�M���*����<c��ۖ���'�v�]�Q�0��^=:U�%/�Q<qp��̪�f��ЭRWV�̣�%�3�aa�>�P�>�噼6� (~_>>�����Z�*܂;����̌v�H!@>��5ÀL�L�#O3U� @��$���6?�ox����S����:O��9������]��T��:2	��{ �Y���ZǶ���R�(�k��JQ)=j��P����Y��\)Q���>���8�2LY-�OQ|%-�K�,{�h������C�<��1��wd�X�Y�����>K�JVgNܪ�C��\(+��{���< (r`?$%���Hy��Ю�A7zg	�Q/ӭs���QX�ce���Gei�Y��M>M[G�e�����x*�8�g�b뻏9:���@2��o^��O]?*NCY��?�� 5z�L��fh�Yw�|֛���X��)Z�|��æ��74��f�i��Nu���7d�l�Wi}\�������F�Jv������G'�/�*U�q(��%��:yҋ��r˸�I�gd���F��*q��L)�o�<��g���f����St���qE:r�j�v(�r�,Ə����+&�y�EdEѧ��ѿ�i��"���(�A��z� P?��,5�~��Zrm|B9v���sS�j!pt�U�L��@�D�|���f��S�n�����Y��JDB ߅��QDJ�pc���;{?�n�����k_������+�c�N����4�C!��~��M�U�*�w����������x����S�±�ԩu����S;�7όې���/T�$�:�_�2g�C��K��T��	Ɯ'hh~��)o~����[��[.��p�9��*�K~2dmw+��Z��>%Ts*T�o܎�l���w��]�E9g݌�ϡ�l�������G�6 {@�K���e[�6R p!硻�韴O7&J�7~x��l���� ���淑��P�Ǆ� {�����!��|̮J�Zr&��3$����9W�Q&KI@��M��)dxaC��t�w�3�(?Ҳ�{ȩ]��ǝ�w�k�x�D�j�_M��u���(�)��I�����6�mF�����{��P�@B6?����G\���?e���*��-�.mLq�EtJ=ه�I�j�Џ�n,C�[��;�_�P_�W�{����X�1&�A�ܰ�=<6�z��}���bt��:��?�{r�JO���-������_<�`���QD�����z6�|S{�ntޢ2������J���-���@ .�k:�B4����4G�_-A4��3hYɢ��MLLP�vs2��F@�S���sb)V��V�3p��G��_c�ѻ�e�x�)��o�9�ď'f���T�x��ޔ���p�� �f(,�RYd�q�:g3.��,��eH�K�?�0�C�V=��^q��S��0�ɹ*�yL��i�9��Q�^rr�ď�@/kmא����Z4�]��<��L���1yZ�P�(��3E�[K!g,��xъ&���8�$��n�d�C/�������P���B��=�ll�����4mn+w�����:I�'�>jɑ<�����(��1U[��IN#���ni*�ÍE;��>(���h�M��Q�r��ȟ���G�W�%��n6F�e�X#2y��{��n��4���~z^ྗ]���j^�1��ZJu�x���=�zFA�6��}��q޺߷M(��c����g�Н�5���e�����K!D����/�ƊK!�ˊta�3]` ׫�[���F�Y�vnƝ�M�j��oH�w�JW�(���܆����y�Q`I��_8���]����*+˳O`��<*,�VC?�VwX5�s�Ş�@�?��� ����4:ܾ� �m�����p�^�л�Xl;;��e A0y9B��d�`�ͪ����x�(:�Ə�Z�&l��oT.ݖP�%pҰ{���p���Nu�{��Y���n�����E�=�b�eY��qؗ�"j�݈&�x���k0��N��J^,Y<��[�{m	���y'� �Ք؜f�dU�53xൕ�)��l��> ������Ȁn�8�[+��#PY��i��zP�r5B�S�;^�U�m��59wT��C3]P~(��s2�<��j�4R4������� ���*SZ�*�2���� �3�OU�rWiZ�i���R2Y�.ðY�uo&B�%��⦰��F�r�]CN�eP�q��X
Fai �p"�c�`�޶R�ߡ�"G% O�i��������<��sV9 ��w��l4�{���H�F��Ύ`=e+X;S{�An��N-,�]=�N7fpήa���T��_J�*X��s!7V{ru�������5��]Ŧ��T�QomN�u,���^���VH��D�̭I�y>���+8��x �s��2T,F�Cl�dV:�^3���
pXGh��_m����C<R��Џ���~P;S]fy�Z㺯��5躣�4��ū�lQ<�?�2�Z2�������S6,�����B�����2���S��p�}z��� ��ކTƐ���g�P�>j?遶��v�������lV��k�Gw���h>z"��"^�-�U��<
{�Q}�m��H�JH�X���ؙ���O���ʭ��b��}������u�CGT�J��\=)Y���{;\���]����0NI�3��8��������>[���k?jXB,H$ȡ{�� 鋡十����a�ɏ�d��4�E^�7��s�:s���4!	Q����=kI�v���?!&A�K�z}J�'p���GS+[�N$x�(��R{;M�a�Sc����E˧�������C�I��>���~�A��%���*Y9��A�(�e6/�������
��oH�-w%���"Q����x�� �8C����۶/[�9��oT�j���=C)	B~m�Bt����>��d�D}����J���N 
�͊J��<�!�so�g��� �U��1�(/��؂��p�w��@���*a�Pl�m�̍�
|�i�0���0�ߊ6�r�P��"P	��AK�zn�\����<@���{d�mI����=f�L�r.�s �!���y�hf����t�B����v�w��m�����m������|$��-f$���u~v�l�B�,L�je-���b�2G�9w�O6w?�)���
ְ����O����]�����O����i<�6.�i�����q��{�Ė=�']C�Ѫ���N���(�����.���(!�/}�0Uu�Iy�G��R���}�I�v�,�1);��1��	�~�L��>�
�O�@�6'�<{��o�X�5�٘y@!RLwi�^*
�~Ģ.��}��F��.���7��0%���M�l�S�T�c�F��m0+M������ ��}7g*���Ӄ������a]:1D��Jl���#��z]ʒKd5eȩyUӹ�,Hw����U���I�\ �s��O�������H�Mu(y��h�$�;��o�����E� w��E]6R-	]��C�9�/���|�X�)<�D������w���+sA��v��D���f�G{�l����7u���V�d7c�9Iь��%\K*3BXmC�[y�L���i�KH������[T��C��R�ՠ�dN�0�B��Ѵ�2������I�������l�}��X��"��qf�g�X��"|�f�yzSǎPT��׃y��-
R�˹����4z����GȹM�gՄ���]�: a��`��K��~�ƭh��T�N�^ Cw�Y�v��*%�)�&��01��<*�Ο�x
ȍ�1���?-�N$�Qy|�Ob���B���к��,��]�����=�OMfW�n��ѧ�+��Y������)�y�(Ke�����l���2�ϐd+�*ƭNӑ��ȃ��V-�= scP�ëaK���A�,��8�F7W(���>��41X�{|S����(F��1�l��Ӏb/t����Z�'�͝[Ґ~*F=d]8M�E&5�y�����+3��rg�����_\������vY|�e��Ȕ�w�6NOHco�k��yC��8nϜ6q=����:KM�Bh��r��!FY��x���,e�/����_�� J�z�����/� �I+"��h��6�#]���` ��8}N}�X����t=�"�Eg#d���+���щ�?0��r�ָp��T��Odm�!ޘ�����DhG|���I�8tTj ���ʰΤ|IY��S�C�a SI[�����W|8����l��Q�v�9����զ�XSm��r冔�kQ���D-,w�+���r1g$@:��8�%e�|�lиS����Q�2RRp6���zfO\̿}��Eu�{͜���\�~U�$� _�	v2w�����+b�2]�t�8=yR釹�TL��M�~QC�s8;jXb�r���L�B��M��.�q3��Bx�\Ae�;���9�����'l�<?m�	���F/A����㻇X�����|S�$$��F �3���ɒ|�-��[���&����q�P4ضTc����0�����+?��a��Lj�#]{�%A�Bz�G1�3�T��q���{�r��{tL���x ��9N��k�O�r��R�ZL�A��>��@�?�DNv۾Q:m/~侅̅�C��
�NVVi���_��6Q� 4�aS�w�jj��H�`ML�h�l��py��n�Dh��w�\���g�E�D�Vz1� ��ld��B(�/��$Mc��I`�/l9�V�]��Q��69���~�:{A���"�#�:J1�7���@�@��\E�@|��	o�n��a�,K}�9%�M�\A��:%���W�L4���/k�7���Ա�g�ޮ� �hQr��C���@�b�{�1A�c$k.r6�"1�0h����}z3x���}�q��6I̡(��V�Rݥ�=�M5�������3��k=k�t�����6In�;����	A{Քi�^`썵��Bwb^���݌'ӷ��B�d��YuH��b�9�fi�^�B8�Q�m��-.!h�LV�|u�,x#�G�^	%�X��-ͺ#�h���Fj��s���&��%�E��A�ږ��h�S�O��`D���##/�Ds-1�[��dp-[S&���~#�Y�j�)�ZF�!��T�}���HS�#�LrTxg|?�1�|&�Ņ7.��Y��L����\Y!q9tf�ɗ�t�.g�t��AI��Bьk���~�D�M��� �O��/@aP��mWU������*筁��y��Y#�.�rE�����Wv�n
B!�*�\G�?�fF|KN�eڌΦ�l�hi�ܝ���@���iX����?�ź�������j�
.�Ծ��ȶ�vcV50��xӢ���2��<�������'�_���=6M��b��x��	�鈯O�4�4盁m���2��4��g!�#s9a���Y\���.8�)�
�b6XV��|Bg�q�MsA�~[�v�a��q��>���!^£<Af�D\�&i鶪���AAa�����t�N'=��י�hW��5ழ�
q�E�����������@G�9��ZT��%����M�R9P��eE�D���+��1RI����)2�-�&�d���7Cm0�9T�!�{�h`)��cRػJ�~��"��EۀιJ��R�/���Q�FTX�M��v���99�<I4��ژ�Xmh�d{���mcU�I_���g�)��>Qf(�h�
9�g[�W�Q�?�
�k��z�����MtM�c*�y����:B�v��u�X��
/J~4
p�� o,�n��˝x�}w���H�����M��Z�E�=���7�Ӈy`)g����m�E9l]Z��L��(t��f݂>���#�`(��u�h�`�6�h�0[4RAj�T�#�VH�����dzXZ
*��)�:]%�r&X#���"D���xt����s/G��e��~���a.��$Q�7�=�`D�Fڊ����ϓ��o��֩�kː��8`C��-$��B��Z��Ȏ��݅L�,���5_�k�A%FV6��*�����1��)E�%�X���6�	;��$����J�n�[�5 R5M�E�'S!�Q٢,�'��>�g�g�����m`t�l�#���w��I)p9I2)R�0�U�V�_��V8�>�C>J�QDf���K=B��択_�A5g��4���� 
4����{�o�3����'O��%��u��ϕ�=��T��ߊ�b�|KP�[g��|@�*ؽ�܃��Һ{�[��8C�@�u��m�z��e?�߲�k'e���<A�g����Vd�s���㨨'h<�}sqw�%:�K����,����C겑�3�3|Q����8X�s���]��������_���0�b�h�)ݯ�x�M��û"�E9>ֆ�,��e\��;^ClbV�/�^�� XF+PH�DІ(��n�L|)��<�|n&i��:��AV氅� �@@<Wc�0U���p(���vq!;�qS�t�:�}r�)u�B9���TYc��\�v�4	�
�,P�.�0+�=���R���~�
O�X�KL�q�B�].n���D������?��=T�n`�c�B��Ӊ��V�X�j��ЅP�����f��$��X��iD�V����0\���o��Z1������kE� ��!�
׆�a��J���)�=!����4�u�rM��̷] +[;`4�
���QNAt�4�Ĳy���xش������6e�U��ܾV�P:�n�#���P��:�v��D)�� �/.��e5w)WS�n+��O ��� �Uv�r9����pvo����h�j�,�8�A����(P���l��lH��0R��4���M�Q�5˸@��ċ�:`b�4�K�i�/�|�JM������q(���>S��9�;�X����?�HlS<�Y�3�� �'bl@c�X;�V��w����}�y�4�;%-�.A������;;R/�Si���S�� ���`u
{�1�x�� z�� 10e����d��溩X�5ڂ�|�<��W�|@1�\F��ʏ����v(�0�i����Q&��[�ꞁ�AJ�ƹ[����s��g6�)p�a�¨��4@�,L�3�AdC�Ґ��� Z�vM���}�x'�܋^�ExmMI�>��/�W�����S�r_%r��V�H�8F�@��Gl�q��:�	U�U�����qЁtNc���]�ё�R���
�UUS3�e|{ 6���T��y�(�1zzdm��Pfi�Եsf�g>���Yc�� 4^�2��^@wl�ܘ(ed�T7q���� 		T��Ǹ0u��UW*y�S18�m)��4&+��Wr�o�ͮ*}Wv���(�=F۰^�
���"�K�A�FX���V/�Ʈ+�uj𢡊�mRH�,S�\^
u��LUL\���q ��:sPz�M�Cu�^R]��>js>�nZM�1��.���sU�NͿ�u�d��<;<�DUq���P��i@îb�h����-ia}Sw?,��C�']�?��حA����9?��|P3�ߪ��m%�4�|������5ט�8�TEJ�ϯ��j�&��j�*�AoSS��l:�p׃�ҠŮeY�ׅ^iW��`�lR,r�A~�OA�nTTЦ�(do(%А\a�w�-��BA�I�c9pV�+�:R4�~}SM��Hj���<���4��'jEM�ޟ�}�zS������4؃/[TR������A��!Z��C(	Nc��뎶V+h��/��M�k��N�C5z���]r0.�s�y�a��� � �
�CE6��v����CΡ��~Y��[�|��ֵV�ds�Ɨ1���\ԀUѢ�|���Ý�48��H��\��	;F%A�ov��9���y�lҗD��忞!")�|��D�h���rbm�]g~/
�)t����mh�E��3�����^�*�ǌx�,�#�C�M^+�P�"���]+��o]��Yj!�J��[)���%3�g���n�g� Aכ�ޙ7��M�9�ɱq���ހ��i,�K�x�F�9gD�ߧļ�7+�*[�)(�,�[��$���!�-�N�Q�����ɫ�#v�J&���y#��P)���f�l[Q�'�ﾣ���P>)�֖��+���[�r8$&]��gV�6K0H"#sr�2zƹ,B��}��o����"K��_�U~�0hN���ov��T�yq�8�}��CC�㚼������z��e����h�+(0\�.Ϻ:r���o�V_Gjn��,A��&��cU���WPx��S�=�\:沮n{��
�ϭ���Omx5<+�τ.�����,�i�zI�7�9>�&���?`Q�H&Z m��
�0���6��iL��J5g�M혗�u`Mvj�Ff�Ⱛ8�fj֗���~�u>v�[V��Fۧ��
H�!k�t QC��+y�:�x>Ã=��oY�W�4�a�a�{?K��z։��S������P
��U> m}��k3��&�LxM-���h���	%���Ƭ��t�D��.�Zz�ϕ�L�p꫓��
D��7�nK��8�V����� <�̥j�sQh�	�;��2�2��p��!��kD��Cq��`Hz���q�-�,v5Z�K�zQ��3���_V�����e��7����*��Mk�̐�_���*RN���cSٝ�0} *-Ж�qG0Aaw/��D��3��UCe����pS�c]6�`�5����B�b��YX����RZ,u�S��j%�?��e��V:�Y�Q�������L�x�|P�������]c ��J{Rɟ�
�(��Y���� �<���yj����j�}E���2�XV������K0¸^�o�|D#We�0��l�U<Һ0�G��`�U˒B���2�ϣ�pŋ���@������-���+�b�tj�@ ��H$e����?�	�-:��ѷ��ߛNI��N�J�KǴ�w�T����p�1�Քp/l��ظ"�5fm}Qbܶ$�R��ڝU�9��[�y�z!w���e��ok�w�� =�@��r�A$���ˉ@���Y�!`�,�-���� I�9,���"%�����ӜSèÀl�j��aT&25Qj)0ll3Q��Q�����җ���R�H��Q�:W�:gBs��Wx�6ƪXi��l躟��oLA�܁[��br�(�������R'g�G��C܆��R���Q��X3���0~�^���o�kRw�-C].������y�HݮȞ��$��k�����o�Z#��]�ω�q���5��B�)`%� �[��Pv	(�ox$K1N5�d�K<W��
5^~EIَy`]�-B|ƚ=س��v��^n�#l�AHlh�p1�D�.7�[c#M�~]������Z'�-�٦���D��؟�� �$�Ԋ��q�X�Q�Ml��p�#��`�+��M(f�(��~<�
��0���d� �1_cZ����� ��g�!3B����kq7i�1PX�5ʗ���I*�XK�ZRG���;G֛�F�̸�������������~"5�X���Ǌ}�a� -��F��_t|��{�q����_������VZ��J��S5�)ϸݎJ�"(K|g�q(������h��v��q'g�e$צ:�I��r��;�GX���|;8�,��x����}#�Ꮻ��h���]���K/q?���~QZ�ixT�tV�I�x�X�൰����|�		~�y�����E\��.�bE�~=��
�D���ݿ�U3��)��k�{�TB�)&���!Qzx��1~^�%Q��.o�.$^�T�L/.C6Fn�� ���VgPH�Qw�Û}���P�)f��k,���K_��Ӈ^� "���P��O	���W~�\Sv�J��$ΜA��Wέ�]���Fd9����n!�.��aU���&l�pj�x����e�r��
�
9��-~�f��fQ������At����;̋���7��bоu�.an��'�W2P�M�7D��Q��s��/�_��9���N~���,��z�%�}�t3���T/�]W:����O-U� �� �\g�j�%;�(g2�E�=�I���M7f�VX��S���(:䧁�g�e	����|�8���
�����nñ�HU�p�:S�ul��I}�X���O�ޙ�)zwI�[��T��C���@	��c(��L�sa��H�i~�E���������a�����a�O��O#�;7b�a5����R��-Br������5p�=db��H#L.��A��C���RwU�k������cQ�8we��������G򍑸1�%Ԛ�f���j���F��%�X����P��ΐ�Xx��K� 2�ɩ��],�5N'T�!��b5]�<�X"i_�5Q9W~�uIj�k�<��^����� -N�d��gcIP�����o�G��z� �9��zX~�Ƅ��-���ξG
�&�`f||y�+#���C4���&���ϫ *uH�h~[�����rk�z�f&9>�����i�o�t �훜z�u&�ɼ����e�%�c����:ԇV���SJ}�u�[���Կ�%k��x���+�Y��`=P�3�.��.�F��D����������6��Khѳ�NP�W���p�VQZ�)x!?��0���z��o�BB؀I��mٯZ^]ॣ�;�i�ہG�4�uMz8��ӷ����&%�;C��Uб/H�Lc�Z}aoҴ+@�1����M�0�Z�ŵ`�
9��x��H)���V1���к[���m'�M���.���lq�F�*��9\*����+<�Mub�9	��;�l0���{�j蜨�!�E�����a��S$����"����-�Z��G���<+���)����,�����͉�}m���3t�L=��Li���=���o���f����
U6yJ�$�j+�D�����ٓ���{��I�<�����O]������x���N.��E�ԁH�����a�_�O-�v�v[ m3M@��u����I��;��V���)��I>`����8�_ߺv���2�]�ۨNԐw`m ��PO�7��M�5k`��l�Gj�(��Y%8 R�ClRw�p�X�oDj��7W����rkߐ�oks���z��D�
��o�?QL���S����.�1;d�z��hj�1S�'��
�Z�ܣRB� �_�k㌯�+<�G�V�� x�Jț����"/y� s�aws|,��â��+����t�����W���&�3�TyGfW���e A����O�qSE.�\?�����J�c����=䊉�/DrD��qd�ji$�o{2t�="o	�2�U� �[G?�'I���EJ�3[��.���Rx�,C��C+e�3A�b��(h�QKa.Z��Y�R�I�����	?̀�BNdzf�xHl�|��o�&�F�>��у���1��>dݻ#�(;��K�ߕ *O�J^n�j-����3HP}I��
U��^<=�`q�|�����5�J�U����?����K���oN� Gn���#�1WzE�
��"���t�h'͢$�&͋5*~#�Q�d�
4f�Vn��/5g��1�w����Lܶ+���Qj�v�������0R��� /y��hL��F�g����r%,�{���5�$�7o�I�"�2|�J�E�jIi@�� [�2-�����C�M]̷�.��קIpïN$*ǐ������ߛ����.:-#bҷ�ebȮ���[��V>�V�g�V=DxH�cIV�6@��G�[Aζ��˶��}�Z���7͈z�D���_����E�c� ���)�xU�����*?�����eA]����!�g'��a�����8(�$����r�k���߃T��	��O��G�IM�
g#�����r��+k�ѵ�W|�rB�;�[Lm����g��N��
ڇ���qdב���F�p
��43�� �i$��<���_����p�f���)��c�9�ʼ]aYw۱2��$K>t�|���^p(�@p
���j}+�O�`�B�2{�ݷ�1,��DQ�*�+���N�i�c���ҽA�{�+>+�!}r^7#�|��bI��$6:1�1W}�j��^�`�����(�V]``q?��h<���h�2�ǖߑ�A�SNFxO,����x�d��b4��"]li���-�s��P-���"�IZ�'��<ƻ(��,���x֊R�U�&��!OJp&B �޽��l!p�1�a���6o+U�����b8�&U��nF<���0ԼX��v��3����,`SN2�#\�\���u����ʗ�[�kY���ء��S�(Zފ>@XxҼܘ�lnA���rb�MJ�{�{z"��W�lr{X�u?3߃�A��gX?8݂�ώ#]a�R���q,@c�H��jfs^	�����)S���q�P����W>��BN�2�5����YI��.�E[`:3�<�G�1e~���,� �]� �\��y�KþF�,�&��[��*L�fdY���r��:�#M+�w-���-�w���_�O�(�Ev���:�]�[AQJxC�\��mہ����n�F���n���N)"�����%�+Zc!�;�D��<8F�\᣾+ap,�7�����-p+oi�Hl
�@���Sl��	b�HW^mfid��n%x��	
'=����.��J�ܕ�t&�=S�m�0#8���&
�U�q�^ɪ�z2�µ��t����h�$X%R��b�aUTv�����*�(��@�����K���a�|u�j�ԟ���-	DdS�-��PGd��7����ȼ��y�����M3U2�@*S|��A�~9�G�gƓ1x�n��y$�x�͓$�q�o��w�5X+8.��z�p<1l��C֭�^�����d�J)�ަ�D����B$jh�Ǚ�$\q�,��G����}k}�c�*PScY��O���D�F4_�!����;pg���Z��	J(a�OZ����״�Hַ^�[��}�I��R�VI��|qYzT��֞GP=֪6���vZ�1�<�В��kUh�աpl�����?]��ݥ�زmG�-����gE�'e���A��I��N�f���e���i�#�T��o�k�h��w�
g�	�Cq�Sf-#��a'_+�L����ŵ��i0�CV�X0KCh$0�7=	(VrcB���D_S�Gr���:.�Dg�Ϳ��������� �xI=g"N����T~�{�
a�����2�<T�PT{;��֐�{3Np΍�6�f���_��;}��
�����R���p�rβ,���s����KO/Lzy��|D��L��S(A��i��k�/��&�"�u�v�Q��It�@�ҫ*P##:aw~���$s>5k�ێ���xEW3'�YS����,C_#���'�-����P�.i4������A5u�� ��H�80�����J���	�~�� N��C��^vIy��sOFQzŋ�&�� x	{51�������C��vFy�I&�>Q#r&<��_��<mg�I8L��|��ȇXP �U�z��)ĉ�}�N�BҩQ��Tls^r�&�MU��WJ*��3�P�M��*�9�wW\�_���l���Negr̴�(�&]�2bsyK������V�
.�%�@�N�nhǜU�
�phT8ٸա���{�DN�V31�N���N�0���Bh �'��o���O�7�26_ �3>D�l�Lǆ��6:eެ���P��"�&63gKyT�i��D�-U�)�����v��Cb���~����'��6P
d)?���o�&��N��j�KU��vFɽVF���k����/��%�WhZ(J�v��Ty����j�Im�O�5-�^RC�If��<��q�����{��mp���R.泩������\�)�ҵ�y����s2��ѝ��?ao'�
�|�҉��o��^U�:'�s<$����L|���g�05���އ�_`'�.�����P��ɛ]�Z;��JS�IG�\�g�9d˿!j�I��5��D��$<���!��B�T��1�/-�;
��.k\xg.!�r�r�vW�OH�(3��2+b�~rn��G��+Uc�N���t�I��0��lls���!l
�	�J��= �p�pх�����/�)~��T�+���9�w���s�+��<t���7ⷫ;"<��D=��ɤ�?�'�#����*́(�+�3�_�o��A��f����o�>�A�;�(,�E;�n喩=���r����St��h?Q-��;�y����w��.�?��P�҄%���wӼ�["�{�z��D�-��5�Z�Y)]�*��mzY.?�/o1ABk���ּ,C����S��lQ��|ag;.�^���I�b�:z�~~���s/��@�Y|<�y��{R�_��'s0�G^���\ �f\oNH��K����j>��?����R�����z-�8f���(F���]s����:���<ec���FrR���	�AxM�߸����u$_gO�y=b��1�I˖��۝YEd����2Oq��Wn�.%&OB/k[Ei|qR%��5M��S��;�3(<Z��Ac�*w�Fea�7|6v2�~�V��p-�!f��� a.J-��2tf���3�3�T_[��=�Z�a�N�ǽ�#�91asܤto�И]B	³��e�]��&Ce"�a@������5�UZ��Jn�%��M6΢�����)��{9}?l��k�zj���k��X�!��H�GbЊ�Op �+���o=��:����ہ\�v\Z���:��P=+��,�6��s9�St�7�]�r��-[_��bK1.,��)=jk'��!|���:�A"%.��J�#P�ٸE��C�V��qd���(��L����Ľ݉������c�_��sE��L`*�|f�.���]d0c�#T���Q@�'5��h�Z[�b�6���s!���o��<� ����S�1�d��JV��>�*M���[�j��+����~'!��LI���1��U���� 31�D����`2�Q�}�ȼ>�S����ݰ)�	5L=õ������R�����L�M���0�X{r�|�KYVe0tg;l�������[y~���T�y��-4F|�j����YB]@���}�-�b�bt�oǏ��Š�L�+'���=��T��ҏU�`����U�u�%��{�&�D&&�!1�;�|�����6�����q8��N����R��j@�)�_+�������)��FÙ"r���-�gj�Z��1g�9�S�c�������09��p���Y�<��9Sl.,u�{�?�;�i!�:�j� ��.<
|ZaX�����;\V�/������e��B�2 �k� 
k��;�Г��w]����c����އ�Z�aQi����H����h�v��xTy�a���hd���}�M�Kb��}�Lw�6�C{�^UfxUS��G�'�Zc�q�c \��p��ų�i�g�d�)��4%���a^�QL�z��ԑ�6��6�]Y�B�m�	@/5E�e:ׇ�A@o�5�����@�I�?LԒ�������{�dǲS�3���{�Ӕ'!����MѬq��mj[��ۄ[���Q�
�J�7���ϭm��`8��9�n{{��[�+n��lY�Tqg�2��=�u�8�F2��_�`9j�K���ID���a�z���0Pd��p/��Ӛ�z�2R��P�S8�
�S�;Q����`4��K.�����8�!�b�5s����8p�i�޸�/_�w�_����mR��(�M	p9Q^�}�������yk���˶c
���_�����R�\i�<�R^K���Avr�M�֝�Dn�_�$�#�?�Rq���n:��� ��/�i��d�n=�>>�q�"��� �ī	ة��3wI�4���|L?a$���B�����ݮ���u�;�˱х�����_X/fv�d���?�[�e�t�b��{T�b�1��ZFQa�:d�*8�/�)���5b�v[��X*�f~z�c^f�I˖�rV�gi:D�4w6�]Ϥ|@Cj�$w"�YO9��&�(PyȒac}���J�I����C��U�f�Ȧ�������:���8�7�jW�fl����ńb%�;{�v�H\V=�Q'��3i�89m�9J�n�b{ӷº����	U_�c$<?ژ��ir8���B[F:�/$N%���ꮉ�T��d�'�➿X���[y�)�TvIK�(�'�v��4�m�f)�nj�ō��ť+�v�B�\�k�r�<u=~��:vhL-��#O;\���h΍�	�ţ�iv�5j|BY��E�{O:x=H� #C����X�m F�Y#��L�dnwD留%���v��}��FIFx$6TTYH��wM+'��ag�F���]�S=���<b��/7e֮Ew������1`'���͘l
�Tn�������0U:Q�(�])-����ع��*ţ��+j����o�2�}�,�j������6"1�H�你���?h}ksF�eh�fg,9�L���9u�p)��o`K!�B	�y�D�4	+�n�;�Qe�L��D�O%�`��H�w�-���2���E��Һ�<2�"㖗��rqP��?&��n6��K���i.�����(Q�V��Q���K���du>0�y+�VTÆ�o=	�+��9��=���eAi�εx��v��f�L-f]���L�Z�X^Sˆ;;/�P�;_>O��xJ5~?�����x�}ӳ�GHLA��!�����'�s����7�a����TI�ESga��c��[9��[�u #Ђ{
�VEE=�cRx-BG��0����3ǻXC�b�F_���7�>�!�Z�{����m�.��se�M>	A��� d����� �8;b�7I_��礫� �K�a�)7�D�"�ɻQX��P0��F+������ �m�7��Ŝ�m��1S l�]I|����� �0���n�|Ϝ���g�b��10S7=���s��&"����-#1�n���c�}Wi&��1(�Wޙ:�$�gauǽ���[�S��Γ=8�r�U�A�	k�dҽ����naS��,��6��%���a�w����_s^㓁 {)�a�aG!7�<��o�m�H�S�N�u� =d'd�N�1��҂�>���{��#����F�M�=_#�饖�����/�3�!+b�Ou��?��e]�0��톑�r��dk*x��O��.����2�0g�5c��ڴ/D8d�)<:���o��}[�@�21 0�z��#I�cq�f��aR�$�G�I�?��Fl��qJ|���U��Disy�t۝���ڊ��r!x<3���ө�&�G�h*;�tiL:=�c��~�ޑ]���'@ٔ�&���"4������B)�o��ř��R�dp���+)3��E_�g��M�t�� cv�[x�)qSr�vs��b!������FQY�3��kM��ͦ
4�f��a�����9��/$B���m�"�īCs^|�D�
�U���^Q�4�a��(2%yԝ���� ��@q�h�R!��$�BS"����g9��I9��_c�8M�-ЂGH������M`�D��
9�Q83��C#3 �"�����S\=8�OkbP�C��0�*a6�����!T�@�Z��]�U����w���SP#�=j���_Ͻ	ߎ�r�A��/]��&n_�D��4u���F��?��i�/�����3�|]�'{?օrJ�����i�����a���)�i��i�8�C��I��8��ex�W��"ٓ���N��I�#ߍ����D8_�T?I4d%�}s�q�f��]Ӻ,�Bc+�ĭSA?;���Q���_����I��)ͱ>��mtd�'8�v�ů�7��>���7��}��XiQ�a��:[��Ꮬ<G�R�:���i�=�y���m�Bc��w�Y{�j��E�:������n63��W�sd��qs�����J{R8#��$o8��/����nX�-4H�hUw���q"ZeW��e��Mn$����F�΂굇�k�F^3t3�5�W2��"@%%J�7��1lu��6y��{��~��3-�,�QpL�jIS�,�!�|���#e<(W	E��ƺ?���8%��0݂�킃Ԙ6Zz�\��ġ��)4����������Z�g�@��޿��Zޕ�c̘�hNp�-���]1��Sd#�&���*�fĿ�0�)���ذ�ns�pt��g�%����������+pS�@|i	I�)��mb��S�(}>.E%�X��8M[�]9����q�RʟZ�J����Y��`!\��3��j|�#T`��B�6�E�_"[� �u�v}�ɾ���K܁��K��	C4d��i��ݝ_��w�cR2GW��,ܸ�� _*���u��6��o�S|�	�N�_�]�Ņ�w���c'��k�J]�	=��BJ�48�-���ye��1�o�XN�3������mv+x��
��^����|���~��F���1�{�_w����Ζ�B���@(��X�1�!������O�:(��8j�mݒMH#�Z��<�
ğDy2��4v���w��{����:�g����W�y��F�CB�bCu'���9�W#YB��fD�S:����6�%�����H���#[M "4g&����&�������K�|y�<��'0�&�M��T�,��+���c�~��9��N�L�kH�	��z��������?��h%�4�����AY�$��u�c���(累k��r$PM��A8��̩�s@���ة�ei� �eo�=����#e�J�	��D�=��]Ж� �A��������4\�ʍ�ⓩ��ō�)�@3]Ca��Y�� *���p�b�7	���{P�.���$֔���U�<���a�ߍgO�:��G��C�Y	$z4*���.���I�o��:�Vb@�r׿�HNX>8Ѣ�J���S-B����]���$g�Nfpo�Nmd�9���}��K��%CP��x��t���Bo��
-�q��Ej#����7���U�"��O�_��� ?��g��bD�rߤU�K�������)�d�n<K݄ݴ�, �.*��!o�׉Hv	�s�K�kB2���3
��Et^�t���K�HAR N�7vW����)�Nt��bV =�:���vz����R���]\���Z��
,���͆����&��lK���O/���_�~a�S��4�
�f�0��j�dk�?h3�W���I�o��
��<>��ի����,�֫!yK�&:�DbY!����1M.�����i�+�(d�$����9"L���_=Uf=3�]�s�œw���}�8q�X��f_�j���`����l��E�u��&�$^/ȗ�Oy��r~�����j�#��j֨��ܡ/XZ��cS5��$l��BZ�}�wb,���F�{�#�����>� �@[���䂟CX�ϡ=�[1C���!K9��ZX�f{X˰r���oK���> � ��u`�%�6h��w���B�Â}6������Ԓ�r���@-�⤅�t=�x�3��C�����|R���e�i۝l銬���T ����	g�]M��I#�I	���6�[x��8��*��8�[c$>U"6�y$�E
�@T0�t�/�7G��g Xd�	I��NC��_�1J�XǙ���O�=��9��&��;���4�����/dS5�f\u( ��Q7��]I���3�ރX�	}Lf�͸Ѕ:5����:H�|���k�-�Y~��I���0�K�Ǧܬ���<�&�P��bv��#^��K��f.р8w'uP��[<�HR�Z�y�{�+U�U_�h�S�ٔRz�)�-)��E��}���81�a�m)�b�Z鐔���ǹ.�����On��q�U,G�u�z
�Ʀ_���Ә�S'f`w�'��R����~]VoHh�t�|h��'.��&�����F7u.|e��˯��E�f�^�Hi�g�(�V���D��˷��E2�jk5���B�MZ	���Y�&���i�?!��	���u�؂�w�*`��>[����$��\�"��L�Z�'3�D�U4�/ۧ�����d�
��в;�K~��TN1��֮cW�����dT���w���Pc�o�]�ٱI����>@�]T���+նHݘZBv�X�\��
Mz1�oD��ܩ�ny��sp��R��һ���<S$�g���!��h$�x�{��2���|� {�E�h�H�K]_����u�L������5����FQ��y&�XD�DwO�/��T�H�q�h#��؂u�m���#��O:���bVnJ1����tైF�Pq�V&^��]��%L� ���̶�^:"`�f̓���W^�1�m�KS$˦R��uo����@�KX�1�4E�����O%� m�,
ZD�D�7ZyL9�Ș�!�y�=�r�tQ�>ch�������o:_�5��M�����LsFe���1�I����*U�W鞩
s���ӡ�xy�'d���%����������k�b�Iu�P;�şZ)�P
��>�"�]��}��Cߢ��]��=�
�������y�gD����Ɯ���[����Cj��c�ho��ږ3�y��ht�Yْq�Е�^k=�YI��+y������G���/J�A��=ڲգڧ�^w��aR��t�e���A��ۇ��j��O��M�,��/�B�H����⋜fՍ.̻C��
ف���(��qÄO�'R�����u� ��C�ߖO�@C9��/]U
����l�<�K�r��%]
�n�6�Z��/~��r4���h�[�K�9m��ÔR�Q�����h�#L��g=��e��w6�Fj�`����`k� �r6{w_�
�zS|B��Zo���J�J �%' ǽ_[�x�ZF"�[�]��mk��;���ύ�x&!�h��݉��q�����W@��}��V�����ga+pE���M>�O�'^�VV;h�X�2ɷ]�	��:��n��~ɯ�L�D�e�",y���-]��k@��9K���*�?�ݟE=p&U�\��c���&Ʈ������k�N+�����4��������Nl�ѾO��/Ki����e���֤�kA5��O�
�aRPm񝜑Sc+Lpǟ�Z'��0ʒD��O:C�����Y�2QƜ86E_9��|Q���ˢ*�!!?�W��Ⱥ���w��~�P�M��j3\��b��<��2?W���wb,��چ�'a����X+��Qn*$�	;�(�`��ذ��<�;ο��?�ߎ�`�W�d�mmc9��[�p�\�o���bOv�D�)y[gڱ��(�ԬJ��w[(�{�֕�Op�Mh���Ά�5�2?1�sNl���d�\@��ÆpG$@oH��)b�o���p�I<����kb���}�� �����ǚ`}P�ހ#< oA����(�f��kb�v5cfI��8�k��``��'�v�u�賭�tĨ�w˧p0��W�cI���)=|�Ԥ���U��Ż��6|`�%�]Lg+Q=Y�lԑZh��Z)vW���k�h�\�ё����������Ii���}�э/}��R 12�$b�'}�,F��ʲ�p� ������;F7;�<�4�4��5�Ac�v�^P���v$ږ�d/��A�ąޥ_B�")�~�|�ͩ����Eϐ��I��s�H���l�*�8��0	�Ȉ��S�la���!A�JE�Q���iFZ����Uň���`"K�"	(l�~�J�)�����c���w��G�r���]gx(y� ��/��W>��ݼ擡�T(� j   wV�C�C,՗܇Yp^��,����&Ѩ�c1�(��V��K��͓�t�ɶ�*�K��tzd:A��C���1հk�шɜ���h����ᔊ��G��3���ya;ѾU[R����ع]ǳX���ϫdC�k�q̊<�<3�
!J�ݜ6����"@�!��̍p��_BUd�U�o7��L�B-����������Tn���-���;�ͅ��r&T�]���OH�A��
$�a�ը>�vH����L;0���|��<$V�PV��B��l4����1�.�ތ��Ԇ��P�GG�	��L�H8��S�I[v��OH��E{�MA3%[��۫�.�\#��%!-A��{�8U�� ��[���u����E�u����g��4 P*��!K^�3-!Z ˯�� �{��,�JI_E_h�w,lB`o����%�;�����f�[J��C�s�^]}H"n���b)�&4��x/%�pmXU����B#~:�r3y!��D̟�H�t�GS�uwl�����]�2��4mgL�r��[d�GC���D�w��#ӮqU-	�_�����g��O(�OZ��nsZ��=��ّ����u��:-`d��~} T䗠JC����� �A��(3@��^Ak^ԡ��l$���ŀ~,�>�M��H�壩*��6��U��7O�=��R�+�r�D�`ZpԦC�a�s�a�!��'�;�S>���������*��[J������E��Sy${Z_Ȃ��Fl����HI���o��&���HlAC徹Դ���[�<�����9Ob��5���� �8l���_�r,��X�Q��Þ�)��qW�X_g<���eN��O	ΓjY�*!؅w����\���ă��7L�.$ �����&n�� �=+�z��Q]Ї򖸜�;d9�jqi�:�ΰKr�G��n9�����v�R��ٓ�:��J��Q_0�v�v���R��Yv�V�&f�>
��,�O�I�W�V]o
�[j����̬���H�����	�̝�B�t���s#b��^`W���?�}�x�諞]�e|IB?�{n�P ����8��g�+���\��zU� ����f*"��E]��~>��ưsL��l�ٴ��Ո�!�g�ό�QA�2�a ��h0�5;IDg�K�E�,�V�Q�)��}�Od�|�|쯁��X�c���:Aw[�Pz�|Id�[;4��W:+�^3�T�o;���W��c����
8˫��J����M8Uar��>�w#�1�:4
%plmN�	����Mj�����? ��q������j���츓���>��z��:�2�3݀�Nw�pw��$u����j�DF����^2QҬ��>�b�L�+�"Ѝw�yĸ� �ӧl{n���g?� O �SK72�.��s��T��o�캹*�/w�>+���U�O_�:����7qB�*ә�������9���1^HR���@_GN��h��Q�P���jB�vxX�\È�ux4?>��͉W�B�YS�?s�0a�ǟ7���~��������Vl�ȭ5#M	���l߄��Z�fUj�K�]Z%�ˬ�X��W"�c�M�I�з΢P�����[���")�l�8�/��A~���c�Ӳ��d�?���2��	R���s�5�_�d��aO��+s�1��i�h�P��A��J����A��R�0������$]���"Y<�a��<p�b�PQB�@�E�D�"^�Z4���˿x�2H[6� wh9�)����`^�Ѧ�']��yc�E��R _��Q(&���n�KH{?J�X�b�
#@��,�@8͈���/0^�H�(Ro�`�݇0wf�QІ��]���\W�f0��_W�rW�+�E�g��x�vi�n�j*qg
$��g���}٧��1�E��C:��R��Y��p���1׽�w����������k�"��.�Cd�+�(/�D�RI�~W��j�z�m�f���Z��#R�W�&��j�*��w��SV��z�v(�dc���@��G[1��y����ql`���.����aX&���$L���YZc�	������d�z����c�)G��OG�3��	(�P�W
RK����R�Ńi���
+���0㚁������'#>��y�irPo^��r�̑�3xP�d��<G�f^}�|�S�~����S�
�N?q��s������(��3Q�߽	)��b�����΁>���t����&
v�%-�`x/q��Akf��Q���X"�7dѤj���(B�^1��ҹ5��d�L�������ƞߪϸ� h;�V�OH�l�������K�I��H��i"�Ol�F�`�l��Y�,fO�1Ozzb�Czac^e��~s��W�h"
F�N���:���g�����m]�
}d���/r�Π���S<�Sì޼���8ea�mC�m�����F�Y)RN�~3�3�#smh�]� �b�T�ĳ?�o��ӥAv�`��8b�݀ܫ�R��n}֏����X��%�J�	/�e��ő�ؖ��3;:���3�⻇aX����TQS.��k7I�ф�d)֤	T<k�(�����E�a{���S�D|�S�,o\�6>�P3�c���O�����5��+C�͟�6u�W;����ڂ��_5߯�����a����eW�zkhH=�$���З";��=�=�jJkzP
Л�󧆼�5\���ķ��۫�v�I�/̂<�M��ڙ��kL��.0�p6����r�E�i:�!a��`����$��R���0��/�%����.�T�#�ޖ��tA7O�V�����Ѫ~�/+��2�%P-�{��{����4t������f�]6R)�O���q�-���H��]A  �%\�`��^�!�d��)��rۿW���ᚨ��B�����J��3�*@��U	���g�z�J&x�=3<���A�0w��,�����O5�k��!e��jn�F�tͩ�H���?oUlP2L�F$���HX�g������^I�FE�q,��I�R#�h�.Ze�(&ɗN8��j�J�8�L�����>� 7�#��컪k��+/��;ʥ>����H���j�v^ܤ�P��b�S,,F0����& ŧ����?�u��Д}�v��+)ģ����u��C�3��)�t���YU6-�K%�h�+v�Ւ���W���mu�T�Sx��������5@S�Q&%H��4ho�	 ��J� �Q�yb����,|8+�Ib.���
�!���#G��]侦CQ���x��B/�:�xo�5h���Б�F���(k�ě�eŐ�<q�AQ��5%Gi|�����r������Z�X~)&d<��i�0��y#[��3@��hV��R��Xo��z�f�d_�A��u�D��z�q�������]�=��E3:�B� �1�i����8�m״�(3��63�yG�H�s.b����DS`�E�"3��� ��O��z��[�)�q�տ���U˽�׉9���לKO�G��b�|=M���_�R�K�H�Hu��D��5|�;�&���$�C¨����2,�qe�AC��*�Px���Yc�4!Pz��05�/���0�v��U�۪MDޝ���<͹H�t��>^��b��fWɊcߊiz�.� !v>T�Jz�bo�����;�RO*� ��8MOV�Z�����Bf���|���0���x'�ƨ`p�u���)��"a�^`��r��8����p۹Bj�h�tO��g#?��(=Ӹڣ�1�M��G� F.HG���4���hNʸ��������h�z �jgQ@��B^8lؚ89ҍ֋�� `N�<vk0d`&��&�C��ր��`�M��{�?��մk�'��=� @?o����AOO.c����TB�٫�M�N��$������ h���X)��]��A���v^���}O�@ZKϐu�C��.%�.���cm��FR3���*�BUDn�!��'$�TMw��Q#����D|��\͡��|�m���B�T��D��Q��V5ssB5{)�+�V��%��1�hKZV�hŀ̰C"��GRt�0�Q�|��,?�z5�I��"��� ��^�͋j��t$5g�վ������������A	'�����SB��y�+�娣[\��yp;� �-��u��g\&*m�ϑ�*J�Ђ�$���%�B��MV��e�,_��:�K:%�iL��+ @+'��#Ki��Xg��b{��-��Vn���%,��qw������_���ԏh����9�[v�.�ܰ�-*��)�mZP!�h�+k�F�h�$
ڭ6N���	�/?E��6�nQ���c����n*��ioб'�<7�.p�c��y���R��4r"�AG�v3&�[�l�.�O&��'�8�ӈ=�#b��߸P] ~U5]���ha6T����,�Dɂ��J�S S�A�P��OS"����A X(�g��!�{+�o�F�_��%�b�?���B�� ���A��6f�7p�O�@��|"��� |�\HE���f��0���x��a��5	� .|�R��՜c� ��Y$�!e�˕�$ˮL<�y",��_�N)��TJ�PB^^�bS�f��Ċ���l�����[hĻ����1�/��_�*io�t�s|�ֲ6��T�t�ˮ�l���T�#��X!�N��`������	a^�;#�d��M�C��a�ƲE�h ��g��Wٹ�?\���`�t�:�0�B�Ʃc�L���:�k)�#��4�HQ�Mn�ƷRWKE��[kICN{�e�����N���xlT�x(@�Ps���Xa*���|\��=�C�[h^>kC_s�4�x�kCw����9�ЈF�j(u^�C��027�̫e�I��B�u8�q{��G�.k�70d�%'�k�{H���� aJ�w�$QI>��۟��zi�sy
+�$}�N*����:�zYp�iQ1�wCkz�t����@Z��	�
��5��&X7�l29��J�U��˳�V�
�L�9�ŬFn�����0=�=h��P�1߄'�����8����ŀqW���곊�x���aN�A��+i����\�,�{U�H�}4��]�ә8�4�Ȣ1�UJI�K�.G<.�K��J�K�{E��˂���[�y�ί�yb���~������[�sG��qP#��T�@MyBq^%�&\�	�H��@hAř�����%�!V�HQ��b��[+��3>~C1>O,C!V���,TJ5�gy�RL��8�[���k��)0*���iM�Tc�:uVS��I��a��6����2�t�9�!���-�!�[g>�z��"i�ό�M8z��t��D[`�|��Af|Y�)��=("�������
�;%���u�#!�mg�{�xgj��.�!7�Ny��k4��چ�EK�l����+��(��������
�4�tV�x1���*�j]��R�M��p��6�r;� �W	>�텡�^�$&R��������֚l`)�.5D��d�8A�\�ţ��ť���?�oSɶ�M��c��j��Z���}�­@|�^�mp͋,ԇ�*[R+z#\L���[�M�z4���Ck^N�U��8�N�������~���W�DJ/?���[P��|��m��Q��E[�RΟ��Aj�ap����B6ϫ	����4�v(m[����)[�W\�89����Wb�����}��uE|�|a�F��B�x^�V"a�K��Pkb$;Y|u���'qH�="4���9�`��,�l�bQ0�c����I��Xc�I���d�=	fX��-�9�RFU%mä�����d���%�ڟ�v�g��s����_�e�����s��t.��Y5��y|��F$ڰ4�"��}5wϤ�#S�o����y���CwZ��k�"��M}�/������Hj!:����+��o;L�S%�V��B����t_�:�뾎ĝ�<��\�I[G2W}���dK}����������D�	���g_�i2��H��9���p�
G�Z+����s���s?v:�R[����3��J[1ͼ/zd�-o+Y�9b^2uKL�E��+q� u���3�ǿ���] l����VJ&7����^(�����Ǫ~��,�gM+F^i-����䖘�n��N5"�Ay��)��������'��E�<��������m��i~6
rC�s��QZi�"�D&�*,��*Q �E��`#Vxe�~���$Xa��xk��mrZUw
��8�2Oz�x��G��������vWziwd�'馡=��VcDb"MZn���K���Q��1G/v��2��᱐��_ĝS�>�5^�BW�1m����"�?�
��"-�����d��R0��>���I&F�� ̓I���J�Ƚ�y�����y��Wͱ\RI�[vP/�;��mIV!���Y5�������&�f�������&&�_�[�w��FPG�l��h;��g����d��O*�W6�\�����~���� �����f���6�2@��߭�=�p��X�AK�ϐ���ue~$�( �I�[繸�_������4b�g��bE��F���R�]���
ز�5�!'C���X9���Zֱ�F(q 9���L�A-�67�4�5'�L]g�d�k�� �1�����/��0�A �!��������N�:��Y����=Y'|w�G>lM>��t£l+�����+�Q�Հ��Tz��K����Q�6���L"p���J�Q$��1~b�-xU��s��3d�y�2����K�=���'���m]�S]�5=ƥ��P��!-�SbO�vr|c�Rgo��A�gp��P�k�`j�����:&�B=5*��te?G��m�R�+Koh���t%���i��LG��m�4o��V�'�����eK֚��b���PR��3�E	Y��K������j�S�r�qo�����E����t��?�.���Up��|�պ�耡E2={��'��
�}��V\��Dp��ew̃y@���uc���R�*DGY8�账�*��RagO�㭵w������G�:��E�)�{4�`�^���'S��8İsbsC�2�U}�ԟ���:�A��b�?7=�����\yS���u�h��:>��(1|;	#�sPx6!�2�#,�Ř| c]aT��i�����b"��������?+��@Pt�OdW�&�11cM�[;�-�r$�ז����l4����u�G=�'�j��a���MC�XXu"��	�;4-�C���m����]˔��}^��}��c�/M�Yk���nJ��,p])\� �ɺ5�*sƕ�8$��o��20,��v��%N���?�o�ޥ�!Y�B�UOI~�D���S�hʗ�:g"ōu�Dr���E73��ܟ�Z��ɚǏ�7���2뜅{��6S۠NGO�W	�P�Z�U��sF����uN��<*Cv�:�v�����J�ҿd�9J�Ɍ \�po\��џ!v��{�C��aQ��C-���#��l�-��[�ȘP��iEI�4�7[/ƘL��+����慜O�iV�?�����g8nSO����Y�<E�n�<�vO�Nڡ���_��*��\ƃ<3��,q��r�����1�����Y 2�������z�:��lr�����軜Sp
��Ao4!�;�U��cQ��'�.��
7�g��Q6��2x�6��08걘��eC�j]@l &�
*X�{6�v	JH/a��.�M�>���ۨ�8ҧ�㧊e_0��raI㘞ú'.hqA�m;+�� �q��A������r��?8Ɓ=��<�U�Cs�#P��|?T�X�S�Ul}�j8�F�n)5�^����շ>�ٙ�YBÄ%��&��.�焼�^(O��&e�̎^k�����V匚�8���7j>R��}f܊`6�a��i�B�
8�����)ܾO佘�i��@�~Յ6�-�Q�si7bM����
W*�������Y�ڪ{��CZ�=s�ftFW�JV/�q��ϸp)��:>laŞ��<��nd��o�G$�h����^�i������K�ҁO`Rd�o���X'*���_!�����]��wOr�?	di�u�Mv=�v�a��#ߟ����)iM��W�ae|
7x��Жx��J�9��ݾ%:W��q����KR�
���3P����$;H\�1_ǝb$�����K���7W��٪C�[�]�莙��z���/xC���8V���7�K�+�ޢi�F4�Y�ŭhY�W����!p*_DK�8C��2�o;x&6�LM�,�G�$/�� ����E��0�i��Tv:�T^���Y\��B��E��g��L�,�N�*�/��1�D7�����s�������e�_B��?�O_�����(-\���*t]kl���H-���T�H���u���c�w��/�r%��97!+b��clGN��|3����γ&�����yF�����.#���Dh?���B1�D���#O;bk&��m��v��d<\�2Ǽ�03��r]:���X�H�����r��Qw����>R��$�bl�v�El��m�'�n��L�J�ox_�h��'���ݨ��������l�,������G��ھ�Jr��u��7�$���ȳ �
v���#��ܡ�%Ȓ$
`�A8�E�g3ה�F�v2��a]�9���R�_3�Ɨd�J�������
�_��z��Bv��f��r���*$��`�u��cHR�)j$u~��F�%Aq6CXgV���oԍ;�k,��A��K{����3��Ԯ�	�i�����zV�ի؆� �s�n���_Ҳn������U�#L|t��)%�A{5��}m�o+:�w��FѮ�b���/�ʗ4u\sB������D�urvk{d��^�����,���a�j\F�e^��(��R'rrag���}��N#�N0��~t��(˳{��1 >zWb�����N�|*o^��'C,<��q�����?��o}�j����0�~U/�ޣM�g�gL�rjI$+�eX����\7�eCq���-�J�K`���Ʉ{��1�)'z��|{�u��R49[���`��e@ɾJX��yQ�T�p���M�d��`W�lj
	(񊔳�)ܫ��Kzډ�+���r]������<�#�b�q9��0#KΠ����q�r U��&��3"��1�U�WI?c���[Y�����?%u�}�?�k���_Sh��RX$E��������(�t�,z�2��d�kA�� �2�i�ENz�9kd#����^p�-��b+;J[�_ƪ&y��z�sGi2.��%kya&8��a�H�P��k��k�ۍ��K-�X�w���d�F�&�\��6�A��	2CTY�����U_PX�D-BLE����wX}�e�
�B����?� M��/<����/�)X�/�x�J��H�2?�@��f-b1���Pt��hۺ�ڂ���R �"J5��O0���D�5B�����@G)��34�˧�4�\Z��^�D������9
���`
愫:R�<�2��3�D���p&�Y࿮�&�?�-�M��3�m*�Q*���^"�����f���s�`	+�Q
C)��4j�4�� ��_�$�	U��*4S���2������헀��Ɛ��g��Mia�wK@c�e�d�*��AL���7���Q�"\B�iՔ��+2���+̠D%���t��V�-[���G:~��e���?�o��f?���8���������K�%�Ly��9�é2�VƱ.&
�����8	���g|X�d�T�'�f:n��+UL��҆خ�#+�k��Q& ��Qd��g��+�L�$�����C#���a/���bx �!@H��(��;�S'7Y�ˆϤ�F}Vr�	�٘/9�@�gyT�ܘ�i�1.Q�?C(�يf��pp7n�a���{��}��|����_���r�Z[J2F��D�&����.x�8���w�t�S�{^z�r����<�:8���!��,k�{u�(R0k������)�=�/��t�A���d���ں�ף����a;C�Bv	d�<BL���*�4���"�s���N��u�����P��'�I��JX�a�i)6�*V^[Ê)��]��Tf7��
�ŷ��B���y%ƣ�':��g<#i&3��o�W;�����ԩ���S_r��+Po��O2o7xHԘ���Y�i��I���1��GL/�A� ,t���>]J��L�Ӭ I��d^#�2�Q��)�K��h
|�*��>�T+�e��{�@��q��ow�yߎ�C��h�Ԕ3ֻ��� �ze�3f>}N�0�9�{ip�'�Vv�B��2=���#���s��%����K���~�;��3�
_��=r	{�m ��Y�#h�ŗ�x�s$%@|Nfʩ��l�ƥs}�%�}6.Q��m�-uof�_�8����'O(��m��u��&���[��Ar�
!B�gXӐu�)9�>�Q���qwZ��2�N�b�9\&��o�S��nM��1�{ݷ� ����'��,��@s0d	2�[��Z��<S�V�j)��l��(Ƙn�?�T,.1�]�5���ԯ&\EW�_yc����ݢ }6g/��Rٛ���B9(�|de��(䟢���&)a����JD��i�Go��N"6�����<���ћ���ۇb��ܑ�Gåq�R%�ћ�Kǌrz�5 "A���b|� ���SC�����Θ5KS��� F]�6+ v�@�gW�z�Kw��v��|�d�)�!���u�EP%f^b�m�'G������Ô}`_�{QŁ�n���R�ny�0�=�Vw��	�^�b��a��7Q]���2���IZw��$�DN�j� n��N��E��Ioe�s�7�,�)'��|��Ċ�}Ӽ�u��\�n��5�=c` �+�����ȸǥϨk�f;��L�D��;?i�˳"��
�r;�3���d��PT�����(��.. �A�{`jK0;C�n��rS���*�p]v�l]0��@���?�4��\ozK�#��] ����R���3����k��M�����95N^�>�۝j�PC��q[IH���(�wC���wT,?tZO�l��i�#kL*�h����ҙۯ���2C��|��#��P���O�ǉ�G�tO�Bo��n��]�F����=�H,�c�ֳ,��[�&�<�l��;r|s�����gq��`Z�إ.���?d,g��!��Z�M2��v��K�\V�W왥�)
yrL�����b� ����K#n͜����l���eA�ԓ;;e����-&(w�
��J�/��]�y���?n��F$�Y��Y硦e�E��p:J�+X����0�B�v���^�;M�'�L�c��Yyz-����� ����'ّDIUY��^:z�'��J���Ϊ��M#y�ǐH����<��e�g�a� �,cl	l])F@RqS(�ew{���=�� 0	h4���4�^�|�V�n.QS��ndRza+R��n�(�ШT�U!7�)Ǭe��E����y���Og�1Se��-�^m���7���rvH����Âߡ��X���{˞l� �����Li�\���{�i�/z2ߗF��cEw�e�/Fj`�Ԡ�������p�d�ܙ�˩� 7�Wwt�t�"� �Ǣ�D0uBĤ���XY�{�40���c�̬>�e�G7�}���e��m-�v`1w1�ÌG#ׯ�C�4��O=os3���j�몀�{�h��H�?f��-�^�v/zL�[������`�?"O��c�J���C��Cg�\�藟ۦ�V�[ǔ�4���%�oU����	TX�͵��Z�F������}��MM���������@���(���i7�Z���E�%�L�?ج�v��&����+���(�t����3�R�yiEH\��K�}A�G�xkur�g�p]t�H���X~(����@�7�ʷL&�J��mnI����	�q���n�c��şWi@�r�l\��nZe*VR8y������s�l�>�P��W��f�u#��Z!6���Mp}t�c<�I�"C��z�?Ǳ�!��l��4� �������~�Zv���S%���-
@�pI��p�a_kj2�xZ��v|�>m:k�v浶_S=�R/��z��H��:��?l3~'{�{�Jd��\:���a¡���-g��u�oWB���J����������2�kX*`z��"܏��vZ�t_��Qoob����"Fz���ƶ���dQ���(�q 㻈�k����9h���Ҩ� ���|@I�|B�Y�����w2��֊/}JƟ�2_�z��;K<��E_�	��;g�`��u絏H��c��Hkk�RM�\�W؟�Í�j}��ǘ�PWx�����u�S.�*^�+\+��#���"i�,���3��Q�d�ٺ�bz$��Zʕ����y����&��R�U����R����=;�k�/�$?,����i�sy
���z����:��b���uں�f��:��� ���+j?�G_V��g8��p��2M}��
n��|�[}�����֠���-1��u�}TR��c����F�7�)��y�k�\�l�%�'�!`�Z��%37��9���Z�o\�M����s�;)��ڲ�#����8<�!_��̖���d�=�D�K�
ӫ ʜ�Pɻ���g���O��ȊY�Q x�Z����{T�)>l��7��wz��ِ;g+�ռ8ޔ���ˠ���|��U�g��m:�� �m�C�$���h"]}Ϥ3��=�c�6�߾H�.�k�V� �h %�zUq�o��p0���C 8��l7�'*�6g��a����ee��%GNl��#nc�q����u�5�$d��i3}�d��\8�t���^�)�TuK(���Xo�`������G��j��Q������;/����}�!���ưu�����t3�O����1�����t��؜pI���J�xo䢒>�$c�R�U�l�^wX�ߵt�g�8������ɇ5!���BMc��ɽC����O�nإi��!G�׊j�)��5�p��4��ؐ�J��T=U9���~�R���n!�2�O�A��B%$�q!��әw��F��6i��+�8>����|m����0��CNL��w��)��S���_���NY����U5��l}R���C��+û�N�ݚǉ���?:���>�r<"{�<�?��R�[�����F�=A�dP*��	��L���Z�t7(#�wܣ�q��c�.�;劰��Q�oLA�(d&���\X�Կ�7x��Os��B�(N��+���ء&�NA#D�Y�Z2lք�݉J�
���9��Fn�K �>�w��~��԰��2J������s*�R�`�J�L�z��W�|a��R�l�3"�'�8_	.��D��1�!u� ��֭�ѐ��k�M���㽹��P���+�BF�k���9��`��4d�j��ׅ	X&�g���8��& ��v!I�&CF�^�4XC3��1K���%O�0�Ub�lG�oR���� G0���j�%���_������������gI��p�}Yi
�@��n)%��;�X��^c�h�iV��X�E��'�!0�;@X�UZP�����}�y���&Ϳ7i�;���sb���T]�01�T��%Ze����YD����9d��Ȕ�k�s�Q;@R4�Dg��7�.��-L�[�O�*��인���?����!C*��o0ܑ��.v �}���xm;�|X�Un'�[�����S,W#39f�7�G��xK�D�,��I����a�sOD��0d'�����G	Yj�
Р�G��9o�c]�N��Hs�� �/�4<Ĥ�~IH���Q[�t  uuxd -���c�k鵆F���)h�4�9�hC����|?�T%fuM�L{<!�_?1��mWR*7�kY=d���ybTɔ�F_b������p���j�
ݲ.O�/�a���������Դ̚�i�gzV��Hs���it��@��<1��y�UsO����o��Þ��Zh�K�y��V��/�-�MC�S��v	�-4���� ���SY���_/�W���2��3o�5��*:�SG~�Ě�SPq�C=WV�b�m?����qza떵餯+V��͹�Z0c`2C=?G
��=�0� &;�S�l�25M -����G�����(��)�/�I���H{����u���*\�-Zo�}�^.^�"+EQ'[oܾ�?_`d�^J�渝�')z�K[���]`B��'���;����pX�qZيg�z��n`?��FxW�p������%I����O
_K�+;�~!E))5����18��X�!��S�d�k��` �:\e�"��
OO�Msb�j=�2�6�y�m��f�mtJ��?s[�[���١���H>��>Iuf�qu��C�O����`�e�js�Rp]u��8�3�s%�|��!w��]�o��
F��E��8*m�@��d?~~N�Za�Q�'Y�iLp���Uy���xg���6J�RH9X�rA���(1w42�4���*׀�i��J��FJֆa�ʞ�7GQy=������]��n����M��aM,�RY�h�e��G�qKwx@'��J%�b�@yQ��n�6%�^ALa��/��ԥ�_"���ψ�`Q��{�4��S6��L�+�A[P��W�er�f�����r�W_�#�nf?�H��Jvq�AvV�Z�G5վ��~��%

濴�\*�[���5 ��
+RM����*߳CY
�� ��ٵ1/�Z���~�L��2�ӹ��H:(_YN�XXF6�;Z��[�6����9g���щj��.��j3]3�}���o��>v�x�~K5�RlF ʊ8���B@n��k,5!�Ic�ժ@GY*[��Ղ����3KA���<�����Zt�l7�&���:HՔRɉ�E�5���G�?h�|�����u5�p/��ծ_�C�v{��SԠh�悇wK�Y��}��<�ݾϩeYOl���ܢm���;0� �Ш���r�����nQ���W���J��cJ�G_YF2�x
�W6v�m]Jf�
I�1����>]8�q�Xd��	���팻T(���0�X=�z�djX7�e�����i[��m2JDW�ϊ��'@���D��{�&�����t���$[۴�n��9)B$؛�
��<�V���:9!T�C���t��^�ufl׿$��݋��oX�����	�a�Z�F��Ӂ!�����7�h��U颐�ʔD{�(.����1�+y%$ � �ݫ�:&�a	X���ρB��SV�i�J��s�
:%�ήN�4��b�}{�(���t�M�GyLK�G�Ɯh�������������<$�X|���ךM�x�͜T��Qm�S������^�_e��K����{��URa�%�3�Х�m�h+�CR��L�{E���Xґ�Y���j�dj�e���p)�]���[�j���e�� ּ���г�7�u�0�=�Wa�<���[[�z?�mݰ��� "4B7���(��"D���[��n4��\���g�CXxE�Y�k5a���"oם�����4����7�Z��r@?cD�ҕn�Q��K�L�s�lq�H�}߹�[��x������-̹=��|^ oW��Ȋ���j���}]�$y(�L�ӆ���p,����bb�m)o����MY�Ƈ�oٝ��)j�Q�H��٫,*����L~
�B���A�bF��m�l��.�.rX�j��W�\�����Ȗ���!�����BV�ҮC#���9���ܙ�k� @��"2\v_��cy[7������@NUX�����u�p�sg�-K}k���aIԪ�7�Ք,�]R"_rE�2�uBD�3uq�a5�����M&�$�T��Dk�Ȟq�V�N���y�p\c�A@G�9�V�	�T�_#�N��RQ9���@W|6A�<����m�v
��-G!�m�w<D&?"��4xҡ8
x������m��H�Y�X�5�x趺lKp�~8:��#T]Y6v��Ϝ��ɴ$.�pݐV�]9��%����D���w�7bD�\��w+ �L���al�5����h
��T�}���ⴖ;;� �%I'dS?51'����\�?Q�Sm���c~�IGJ�g�0ߋ�Q-�?��'Nl��O�j���|�]*Z�r����P�Ő��ˤ����(���gV*��reF�v>	���s��<�r%�=(�"tv�� j�-]��J�b�_��<�x��'�����e8����ٚ9���?U�L��bC4#�$��CË�C�os,�p��U�T����F�A4+���c!��
8���^\�e�I���ǃ3�8���b�GPFU�:�g(��U���=L]�-GE�r�6��57[��|�d9�Ѽsm��!��T�]3�ؔ���r6`?���D>L�u;B:��8~��'��s���B��a�!�� "]��y�P��H��)ռ��D�0`\	�4ʵ��b���<�\c�~�� ��/r�R�@ӜA�T�����pD�vw����y���:�		�Fa�����:�6l��r#��@8{�r�;�LW�_4��lj��ꢨx��?Go^��E*8e�d�[�<?�v�M���M��}|��?W��&%�O��R��U&�5���8���Q4y�y�`�N�7�� �c)��r*�} �#ج6SW%��l$�s�4J��p�U[������Y.�� ���~�39IU"O<�ԉ�� �r)E�7!Z�jsr�g������]�eBZ��T�{{)�s�P�c�ߘް4��M����*$T��Ǩ�2�	u�WP�o�.�݌��]�T��fEz�%%ˆ�G���%�N�:�d^c��91����T ��N�������9�)���nk��º>�$r�Q���?�H�ґ��܆+������P�Z^��V�/��8�Pd�*1�_�ls5�OM�ζ�(-Ľ����~�3�Jl?�5$��=ϙ!��w����G��Ɓ��7��YE �j���e�m�dO"�ȃ��:�F�]��oh.�H��6V�V��+tb��Ӄ����Ia�L K)b��9Y2�Jb����S��9.'���/��6�������>$�u7'N���%H��{�ם��[pz���@�}8��s�z=<�*\�Q�������	�X4�: ����Yg+��F���%R�zkIz(���@,��{�Ͼn*��Þ63M�EG�2��~��X���Jy��G��${���|w5�a��S��r����s^��O�֥�nP�l)gK�V�Q���5s%r)�9=%�u�Ψ,��KW��1�*=�$r�cH�I�}x�^
�E!�޾�<�h��7��z������;�hA<�v�����2Z��|������ꦏ�E�ȡ�EJ��@�}B]�/�O���e\J ���w�\����\#�kY�,b�k�kQ�bܔK��Ջ+�:��W�c�ߑ����w��Dť҈^y�U��85��G7@��5��k8�e@�.@�G�"��J:uB��XҤ1���=	B��y̛Y�����z����t1��В��mR�Q��'&��c?0�F�{*�ξภ,l�a�DR��9Ŗ���(B�_?jq_тE����H���.K����U�~c�voH�0[�lh).&�N���^� �CF�߷s{ք�Bh�kQbm�m����5c�I�cL�_y��sN������V\=�K��W��q�NW-��@�Y!���M�/�?��fTт�d���@�vc��uB�s�T�V��%'��xH �Y�.�59�q��5ү�GT��o\]s:q^O�Sc{3����`B�"��S�z͗=���VjƜ�􈎓X��Gb�Θұ��	6��N5T5e���:<� ]�1΅�e;�pv&���&4��.&iL����Y�w���\�2��}&�*@��l�}��}�����r���0��}��w���ͺP�!�c2OCפ�ȾKh�GLz�s/
�����$P�5�Gb����0[�
D�M��=�f8�Ԗ��J%�Rv_��1�`2���	=1#}��W:�D��>�7g�f^B�+��3����������a�������٨���TABܘ�%�M+�M�*�RL�k��l=\cK�1�s�-1��xH�$���=���!9�螧�Lj0�J��$���>�q����"NoP�m&e�  m8�%�:������W4a�Gj�P%��a��ⶔ��C�xQ �c�o���/\����QlN)p���_( +?�6� �h!����
~�mh�:��TRz�\``����c�U��֞�xg�^�$���<i?�jB��(���׻5S�"̹���X6@�/��9��� }�b�s�r@'	���hrh%��X٢�V�9�Q�J%��Pf�,��p�N���o# hZ�F<�&PC�z%6P���l+����S��]�)���Ƙ�zl�l�^�I�n�m�&!��R�[d��Ɖr�S�[��>���]O�I�
Պ������u���y��.}���=꟠�ĨJ����|�i�~re���n�f�i�h�}6E���H���+��x�p�uB93e�!�.�)\Nn�o�H�BaOJf{6�Ce!t�D�)J�;bv���������HGG�(�s��F�*upmN�PjQRn
`�l��=�0B�F�*pt�ςa4�@�qeܽ���:�=�����0��"L������Z�!N�FDgR�#Y�xK� -��MK<�|#M�]��_�+Q;[ڂx��zZ��bά�����v�����&���2�j���;`�[�L֛�Dj$��u�!��1ܐPv��ç`v��5E��9�_9U?�:�45.�|�\zf<UA�˰]kꞑ�<^�҄Ox���K5�ҝ�#(��T���w̧4�2�N�6b����Z���e��k��Q��<i�w��mdr�G"���L��~ס��Nyy[�_�1\(x���W���6�o�1�����n6@Fo�$�t��؏N�a�E�ρr�~%�1!j7���+~3�CU��en�(#�n���7v�� q�7�����0�S��w.�j�mς�'e���anc�0YL����!MC`]�8h����5������y�h&�w�˓�������bO~�e^=���d�5���o@[�-P�!3�د���`��Ex)ϰ�?�t��{���5��خSL�)�q��sf�I��3�������B���[Ū@�
!���Gy�$YV7S`�&��q�*&R� ���y���/֯P	Y>x�A��3>aQBI��e։fo/حm�5�L^�(������rR�ω��24�(����tE���6]���T��N��Ꞇ����P�5�x/%�6p���C:��Q�	Vi�x?9�)b����d����M%W~�(�Ϲ�[3�,X�����Le[rʠJ��b6��Z��Of _q�6.>�e�o���m�1"hL����G�t�.SY���[�9z�
���n��-��.;����C�.�f)̀�������.,d�p�6�C��KI�}�uY�����u�(ԏ�i\54�=��������jK:��75��mT�X�!1(��<H����2�=��x��k��΁��a,��Ѧ"j��	`9��G�ot.���w"�c<:͒��-9�JlHFb?
3�������*�.��W�,y^i�,3Z.��`땕!�O疕��P2��r��t�t�G�%��~�
M��]�S|�԰=H����7m&�@��y o9�ЂR![x!��5�C��r�i~?��#��3�c�/_��S�.��d��yt��$��Ɠ>J�)�hiҔ�N���~SҚ`�g�
�����G\A��c� �v)�d	*L�qPj����x���&H:�YŤN��=����!�{X��U*o}��Q��Z5�K�ʅ��"��:D�!���P���t�R���3��Pϟp}��`l�����a7�z�8���r��!#�)��Zwv;�m��[ۡ�~��<Z�a,��ya8���X�/Bxd[�!.52�FK��s���8CX|]��Y��N�ju�[eg1�z��!�I�_�W��v��#PTS	0��r�,d�	������V:�h��P����K�*%w���m<=M��hkV-Ð��a�rI$S�U�Njo��t�+U�D�.$^)?��Ʊ ��a���p�zKR~�K<f��.�P8�@|U[�/7��� ���\M��Yq�������ܘ^�p`�e����H�bN�Q]�k�����Щ2�Jz)8��_�!ɫ�����fg�>�Nri�.HH��wb�aur�'/�/��� \c��3�k����,\�y
�f��vs��~�EKZR��	]�k�S;��W�ߓ/Z���u�R1H/m�.U�I��?�n@�%���& �t��d�ש}^��s�Ѹ((�m�ۦ��N�!O@�����
^bQ� Q���Mip�Uy!�DYI�Gp#CDXrx"u�n�\L0|�d � ��
OWo��4�!ͮ���r�������D0� u��f��A�n�hj����������K�̈�ZT��b��v˘Q���3���W`��JA��i����"qDj2�E#���gF��j��B��A��0`LÍH�� �idX�������2X6xW�I��R}s~,l�q�,�&8d�V<�7��������9�;�@�!-��K#q0�L�܃��`H=\�V�h)7ߨ�_s��Q��;�+��M�������e�Z���hi_��*L�{)ؘ͞�?&��P�PU~'!GZ�!�e S��/������g$���],���t��c����W��,�`�7.Bm�������z�9h��x��a�2B��u�Vw�=L��a�A�s�pB��sr�����A����ؑ�5xYa3�f��@n�NJB��Zxw�֊}���9M��D66,�^���Iӭ"x��
*�p��(� &���$�uT�����HV�)��@s:Q<ͱx��Ulx�7�'�.�2��u������c�TY��,r%I���r��k��k.�v�t�B46-
|Y��b��7�T�j��l�>��0x���QR�C����P+bi���
�e�!	�Iv���J4t���z���0��L/jX��G��XP�\v��E���r�_�9�'[�������PZ!�`zI-��q��R�G	fi�%�#~=;�Ic\+e뷘B����m� =���@%��Ā�^k-�Ɩ��݇FC�(�;���=r�F_	p��_m�*r�WW��Ջm
B|X|�Q�F&]�:Y� F�Gȸ�l��g�.��j�w�Of0�"#l_rD8W�e�����7�m����)f��.5\_�|lJ��ͨd�����
���n:|��ۦ�G(4�ن
|>&��H[I��b��(x�ʥ5�viR�6�n,�rub;�Q��A�E�\J6�q�gN�G����z(��ԁ^�E-p�ƣ��K9�����S�s%	�n���cf���rZ�Ё(�7�����\���?��^�&�n5�ԡ �>g�E?3��M���ҕu�tC�<G¢%"�H{Dg����̋=�����\p�3�>=�;?\��gDj��m-liA�ȒWd��sIW@f���KD�����Od���#��(ߤlQ�ތ�+�{��{�a��a�64���+,#�}8 �p��XiÔ4[����� /5	>d��T^Ƹ�
��.�K���ƅ|�8&�Þ�)d��'�"��������n���\�����V-��r5įO��@�i����	�Ho�s�|��vW[$��v�Eۃ��*��,p^�U�#p��S�.U�X����%>���[bb��'
_�4g�v!��Yz̳�qlC[/ ��ˣ�o�y�;��a��G�x�U�����l-i.cV�o�5�.�⩨�D
�(��
f�^t��ya�р%5�S s~�9j��1��*_g��^�X������{{����3��9ϭ��*~����Ql�����|Ӝ�h�NYA�ί��<S�Z�Z��}R����دG"W���C��-p��p^ռP�~g7�4%���P`�{|�w%e��)T�5�����k!Z���}�;\�����C�ه���Ei\Bl�c�Nƥ;����,"���є7brXң�}��z[���}n���R�؛��?�B�� L�f
�W��?�?�����ط�۔�(ZF��,�׋l�Y[`xm
m7�ðG#��� d�{�d�+�dEe�Lxt��9��?�������릛=D~<��8�ׇ����;m�_x@BU��7Pf$+��rA�ß:�05���(H��w��1u�,���6!|��S�`D�h��u�˶qKm{���"|O�[� �S�3t<j=QV`6���)�a0jY��a����Y�oR<x�b��4g{v��@��:�ΔJ�W�1;���&t�ޣ�Dz�j�&�0�H~���(u5K�H9�|�3Y/�������z����Pe|F��騷@�5/j�ˮ��>X�	>@��/����(��Qb�4�l.J�
����y����g�P�ժ��VzW�8O�e@:2�zG�����;��6�*!6 �K#���'4R	�=|�`{����.~�TQq7�FG,6�������g�N��ݙW�j2-5�T�%l��qK9>���=>�&�tWLvC0Q�8���Y� &/�2�F���P�:_9@T#S���%w�ۻ��j�i��:�G֥�Q��e�C���N'�o�Lj��R�����e�N ���"�ĠN�5>B��<=�$~������!y\<��~�����I;+#�S w��P�TՃ|�Y�a|VEI�V��bjp.ʓQ�:����4$U��Z���$'�m"L#X3Ȯ��'@�+�̼�Cm7�]4�+M!���!����8��90}ݹQ5i`U�����
��݁j�f�|��dS�M,�;={���EJnJ�4}I+M�T�Pz*ۜ�L�G�i�
�:2�>���0���R4��\�z��n�9�oQ�n�Ȱ@���Q1b�{;�q5�����0�{=��|���	M���o�x�(�@��:���_�ǏZ�w!�*��gj�R�_w�r񿈲���F_��w�ɍI*2����:2FM�\z+)t���-��o���ĩ�YG�4X^C��5���`����͸����<�;��׀��>ƶf�1V]E��*4[�I��:�À`�T�>�G��F�����VH�	ƍY�1RP1�:�L�֑`؉<����̔��{Ǹ4V��)�g2�o��-��:>`�K��Y�u|�@!=9A��c���mw@m���D�R���P�l�B������s���%;$��P5j��\a�<�Ҫ=U]�s��5��rխzt` �_�_ �_:�U&4��7�J��dg�S�MO 5{�oH��Q*|�M���}��S9*5䤲�2"�)�C�1���P��Ϝ1$���+��OP.���9�v�W��wjh|�ۖ7���H=��+��V�Ŕ��&M���q2���m\%��.��F�T�M��H{�9�Ԋ���ph(���&����{!M.�s(u�&ni��0bJK����BEk����I�w,���ĜM�黔a�s�/f&RDjDI,O�G�2Ymu8�������<�~�#�g��1�r�<�@�أ7� ęLm��R�д+)r��o���PLN�t�<l{�ǘ:��q�¬i t�C��+��6 7��K��Fk���K�hg��V�{����)������6�x�anJ	�O����GX�ȦV�����d���/��8
$s����i2��H/ރ�7����!�%k�CJ(�ݻ!8�p�K�Ľ<�z�f�ƾ�}X
@������U75��3�*(��	8���OU�@߁�r���Qc�YKE���c� W7驥�D��C���R&�t�8/�H���H�Xֶw�"O�t���K��W�R��̹&)��,�Xl.o/�2FzH@�>Ú��!��]B~�,�jj� ���N>c��4z�6�6��I��l���f���>���6��sf!��򇣞�9v���"L���7���ț 曞6����$>�3���Ր�p�W�NW@�����quG����Z1�×:�L��b� �2ʖY���1��&$<4Z�x��<��38jQ��*���iᙾ��[�L�c%���}�`+y�- �`�:�+ �LKp_�0s.�����3��X��Q|NBi��[~����Z^st�G,����|��z�7"siSw�$w&��$)l�|��ۚ:�`CVv�"�t)��f�2��w�NZЈQ~�+j���Z��)T��Ƕ��P�Z4^�\ʠe2�S�/��M�֯�i���،�T=:��3��=X�AY�\b�P���mփOm��?�V��"A�#��EO�a��ӋdX��0�f?��=�HL~\5�r�����/����w|�Rqh,�1�%�H}WSZR|����P_NK�p�o�q*�W`N�K�D���$;���O]7�,�Њ[��������<�!��EO'Z:��t#�����	4k}mT+ ]����Z�u�J=�� �S��M��Y/�C{��ÄvK�:�k��M=��|SNv^��o�D���s�b�	(�h�.�<����FɆ��Z��<�4��d��Hf��TŸޙz$�n����C$�f�������#��:��	�n��sA$x��Ȍs!�R_dY�_��qB��\�y+��'��'�΁���Y�:E��q��$n�X�WX����f�����"P�ʲ����e !ha����+U���W~�%d�:�92M2���mj��L����P��~�t�<h�GM@��5�[|G,�X���v�͇ˮ�����b:r �
�@�9zD L"�f3M|k��ń������c�Xc�^��)�
e��]��c\��C(M3J>�0�ou��~��C0��p�`{d�k1�7`C{�%��2�^l���L�@�� ��z��Q���eNlir�5<I�784I���K!�&wp� �Y,��Cm��L��,��o�-W���.�߯D_��Y�q�L��EM�7��e<F�o4��7 �P��1�:��+���A�&Fh���f���$��9�L�3�@Uh���EݚhN����[7��ª~v���i�FҜ���6}y����e^���\�X�"��(Bb�[���*�{ <`�Z�E7��P0��-�{�y~*p�j�H�I�Zc�j�Nq���zJ�}�[9��8X:�L�4��2��3=ٔ7�U9)l�.|���y��	T�x�V�C��q镪����
���%��=�N���� ��K2�N���!��Wq~p���~�]���`���
��v��2y���Ý��zR�u4ç%����'D^��Ĕ"]ϵ�"c����;+7���a�>+�������_�ᣃ��/�����A����Z�
8���+�3��mg�L�v����%��Q�/d\�#�yU����UUg(Kq���^d� $>n;�Ӎϐ�@/�"��Ik+^�l��2]rЯ�~�,��<ρwq�,?�W��	�b�.��f�V��F���o�~'�4�^��z�����2���oE�H��_��ʈ�t�j</M��r�iT4�94�1뻶���|��M��@�v��/H�/����<:#4�h�'\��� ��,�D$!��;�?���A�euf��g��w�:�#�|Q�l$�#*<J�cb�]T��JT5#FaD6��"�}�׷�Ř��#9Mg��tB�4?'�����]�V|=�F�FUE�u���:�;Ӌf�-Lf�&ѡ!CN�X�Xjl������y��e"㾫��{e����tfx�k�V>YR���uy����yT��!0����¸���V�^UW��5u�20�=Ӓ� �Ű(^W�oz��)�]{ҷ�Z����D�k���tV���TCpV�L.XE6p�,Y��h��C�-���� EsN� `1��A��롰0��w�-a�-k��2���q�n@pP���|�SG^�p��>9��Y����F3P&��PG�لƀ�Klma�P"��@RL��":-21Q�V�b��4����D��Y-S�̸��=�8f�𺔀R}^�s#���$��h*&0�Eګ�����z-�H%��j2[�8\,ȍ��w�D��_���Yc#/�3�����9O��eꏶ�lhW�m�Ә�4�[e�Ӄz'od��!Y}�3]��t:��{=��B��;43�?N�*U�8b�He�-���L��<�LR燠����IEd�kH�d�����ߞ���8N�#�{�}Ù_��'H �(��A[t~~�������(@���Gc�����u�/�~�\�[Y]:fd	2�$�n� ���3f ��9�_�_�}bļ�Fjk&=7�~��b��c�gN��w�3ף%Zh��p����*~ڄ�D��8m��[�?�
�8�y�_?��MG�*E53~��ж˧e������^��+����(��O�_a0\�㟙q��?��7nQ=���a �����ٹz��y75���\��)��P���&�4=bݺ���+Wl�s���,���Զb�'8�j���:��N��F�;���Z�՟����ﶝ}2�]E������c�M��<����v�l�!O�[B�w�$k$U�b�Z3@��|���H�7�bև���(��j2�dw�XmCa�˒s����=�����!���J�`#U�R��l��r tƏ�.�����'A��h�0��xFS��`[�h1;O��H,��s� o�P�
A�ok���h$�U�{* H��mh�r��.�;H)eel'8r��`з�m�e�3��=nd�Vɍ�k�3lZ�='�^���ZN�J�YZ%�ڤzX�8Ơ��Sޔk����+�%=�(�k3f�Π������-K	k�e?�g:g�}72��}�ԍI,1(X���9�4�2޵�е;�InPT�,@ ���	��{����CC�ݳ�bͨM��^�?}q�O��PL]i�����P#�������I)��#�qM,{ H��d��HR_��2���H���D ���/��uzG����	9cS����&�YY���[��M@��]F.���1����Ȅ*�~-��m���"�R�,@�Vh�W��R����]��1�!�z�c-�%������� !e�̶K��*ɰ@���Iج��p�}ǨK���w^��X�qh$W�� ���8�[�"h�gq#d�1ºe���|�p��ij�J�W��?���*A VDa�M|�m05����f?Yak�H�p��7�n0�e�I�J��i���g{�d� �!�[X�n�5&5´x�		��|�N}tU�O�(�P 4�x������1�3;-j˺�^�i��9H}M�ҋ�=��X��
$-c�׹�7��h�M@I�*M�4\VRgj��ߗ"�>���������=/dW�qd�����e�Cݰ�O�@,2��p�|+�`$/]c/�/�����({����=���d{��Do�4$+[Il��%��䲱" �k,c[���b���50O��%O]�>�������Xs�qҟ�	Njj'U64���O �f�R����9Q2��n�C���k1�4=�O鵽�Z=���69ο�	OIS���Ɏ�j�?.�a�faS�\�K:�C)֑��@�(`�⡀�6m��������䅨�[4�f�|ɩ���Uua0�RT*�o����d"�{�#&׼�v/� �H;<��!�2����Ku��qk��1.�E�/g����#C����,Y�I #J\�B���rS=C�6kə_��N"��+	���`���4_�0��Im�i�_���e�L%��v�@�
���2��R�Ɩ�ɩ:E"d�Q�pf`�/�[d���G�CO|��X���J�����o+J�ʾ%���l��d���a��W>L�V���T���D4�o�D*^5=����e����A�8�w�y% $lg�^�̛ږ
���K���]
� �����)�U;4|7��b���Ϝͩ~�FS��'^*d�m,p�lA��.���5������Nh�G��;gʀ�I�� �{�!��'N��G���|^��� ��b��4<�%Ư0{T��%�&�?	�%���7V<�>'������f˓;���%�)��m��f��̔��v����<�s����i����S+��/B<����k���3�CE1e�!���J�h�������0��)9mE2U	�D/&w>fWc��Ә>����?,M�J ��?	����x,|�`ixx>ي*U�3�;�`41���S�*���vxk��}/�3K`��.�V�yr��/#�i��E|���M��@gΥ��%<c5��G�-a�������Օ�X���-Oy��Y3^�����D9�e��@n�'O_��Π]M)��	: �0���3|fc�U���v��WL�'l�X� y��|F�sSed?�ːC�����)��N�Q��hYI�����A�_y@���D��T��
���Ҕ�b�k�JC{vjڒ��ϤT}�Z�|`�=�����[��`�;�-�"
��WP��c�*1Fk�Y��|�����&|�~�}z]<��XvxE��}�n��(���`�=�ҧ�qW�<fׇ��z�v��!�U�áC�@��.���l�MgF����&�R��x�l�{=������ict摦80s�C>��w�`���ή���bZ���&�K�6�w��Q7]�4��b��o݉�]��i��S�B�u:��shsT��銟ՙ,@p�67j�-l��o~I|�yB8s������@��X�Y�+IMǔ��
F�,bZ�Lq��Ϗ]2`��]��j8�V�O�r	�U�VP~Z*Ɂ��z��z�&���*�/�b���*�L>�9{h�QآL|�l_9��l�y�o�b����G�hR^[ڠ:w�י�S�l�@�R����#H�����bR�[�ƕ.9y-�E��ٞ���R}c�Ҟ�.Ҵb䝈��;�;�&
4��c��(kA��-��F}۷��o��+Z鰈�<���C��s���{���oN�*Y+)��<�P��=h����S�2�����jcU��sa�޸�QG�R��B���8�;V#������
|��<5@z�[�a��8��b`��YSx�om�\�)�V4oZ�Z���)G�N��+�h��Fk�g�y�^�l"A�݄T/��\�R
�4q*ONoLT���@��B.g�L�8�K�
�N7kxa��2�7�a�X���9zO(V��h���7@#�[.͍�=d�}v�y�r�g��𪕺�_J�X
�9�"��}/p�#ʒ�H���̃��=�妖.Y���|��Q���o�����pP�9=�l���N�3W� ��^�!|9I�NssYOD�|a�/MPX��ZC�߁\s�����׹cښ���-Ld��jy�J|UCch�>{K��4]��8��me-�,�,�Б���!�o��@BHPZ-�yc�4,L?s��D��t�K��u���LC1����ufm�b���Q�<�"�����F�y�6�M�s�k�E�q�u8��$���l�%X�z$9���W�w��I��y�$�a�-�CY��2�ZQH*	ً�NX�t��.;��6�ojI�2㸨 ��.*�84l��Vf����zE<v@�n�~��G�6�p��`�ݻ0q@olԼ�A���v7�+R~�����J%������0: <�1����&�@7�u���}�[x��ҐY�C��uX��u���)���X�5-u�(���"N�%_ 
�0��᯿�������B�[������ �� )�" $�5uI�b�t�e�AK�������CK�Nk;�'PԹ�OV9�f��n�k;^IS���<��Lw�yF�Ȕ4{�Ӗa���]�i�^t3y�N.���/ќ�n6gzB��/��R�L���@�y��|Z��.#p���Uz��B��"c7��ʡ*��&��F��d�-Ĕ'h��nqi��U�uQ�D��4���T��yD]
����U�$��k�þ�F�5�r[���?�N�ֱ��3{���(3:�� ��Pt��"�����d�-B{*r���ї�vg�=�Bm��8|�E��R�.yØl�f�p���{����"ێ?�U����J��#�fs��b��v�W#�5W>3j�2�.����ʰ��):j̽h̓��T6��
�6��ޖ6-M�AҎ��һ���Nf�
�c�/Q���#8��m��0�#��h���/2�N.-\y9�����X��=����= _��b�a��V���� JH��+�r�0��9 �}�J!|�t�K>mW1Ǆ�"ڼ��"M>6<{��f�'o��E�}WtV�#����&�֔a�o5j?4���;�'�i|�O���1�-VY��ẶJJ�	@lT(�u�����!�ZF��3j�\�ԽF-S8� �U/�w���ֶОƘ����}�E���͂aI�����@PR_�����|����6��~7N����<�)�tK��(��I�3��ISn0d�D�����IC���!�z�3+J]���uz�z����iR�ܙN�y{���Rio����Z}d����>�%�,?|^��ȮJ&oT���k���~O���qx�/{�HE8�yN �5���z�L:N�V0ᢴ+Gx0�o���2�~�/�L�w��|��թ���s�:<Ձ3�sT�G�^�w�+��Pt��;���������-*1�NU��S�]Vg](���8��mj��T^�a�">k�}��Jz�+������/�LL#�$�~�0��j�B����;q��Gu�c�['�2,.qk����R����I�9�F{��7�sQ���e$h���1u��F����=�Ƒe|Ro��8gj]��0;�i�����WTMl�>lQ�z�����X�b��]a0V����B�,��7����a��4Oӱ��,�eZH�"�n�٤n�2\[��)�hF�GM�<��,�R����&�>K�u��~�k����?�	4�k�l��I��V&y�E-\��vY���Ʀ��m�NPu8�cO�5$�Q�k��L��dId����)�%nXɰ� !��1K�q�s~Aޑ?2�H)�b@+Q�D���]nC�`��#������<&>�C{�
��Cz W�!b��y��p��"���L�7�y�k��g���2y@�o��I����rF��˞�)�k�#ұݟ��ܔ��l�j�,�aj/�`�h#�xg�����6��>����m#��n�56�#�XO�3B��� ޯ4��iw�i�ʧ�XR��o���M�3��v���<����r�W����-��yT����  TL<-�����\������
R��w��l���g����ؘ�>��Ŗ�э�����-)�0�H�|��V��Y��x�R�m@���?�e�ًv_�_�\��@^]6���>A;DWE�+�(���vV����y�v������i���]�cU�A� #M��wKeݏ䪗Wo7�ɯ���|�ʼ0���qΉ�Sd��$�@?����S��_��o�� K��:�I�8��C1b�?:N�Ǩ�wKo�e-gܩ���
Ds���up� ���'�ӎ��6֌8��1�3�9%tr4��!���l=��ہO���1Tm�c&"��։�[,i��F��w8�p��fR3*�᥄��J_����fg�)�!�/�ۓ2�~2��ڤ��s^ ���rsΏ��h&?�=7S����F�RS3:��<o��#σK�U�@�i�&x"����Yff��^b}~ol=6�=�3�AI�R�5��v��24�W	�J������a_�{��{O�W]�&�㩿C�_��U4#�1�@��D��o``���3t����w�7#DZ���r}w�,��d�9	g)�<�[���M��$=)�;��,�P<��KyT����'�L�/{!� ��dѳ�k�)dMTs1���{�`?��|& ��q*ڋ��AF���$b�C��o��:t�M{���.�ߎ�v������,L�H��=ti)pT՜1���s�ղO]���Ѐ\���B��g�H�>����r��C�֫5ȳ��e���h �޽��_�¿1/����j�U�!w��Y)�h�r��8o\���` �NP0�'�^����-
��\����L[�B͖��E7ޣ��e���-yCx;*g���8����qބ%���yV��I�����ꐔ����ݶwz�,����r��n�u�&q���/M}�$�1�-p�k��O�wo�PV[&ѕ�����0�V\���ڭ���SD��|1"T�u�Z���j�C�����ic�|�EL��	�@�l!B�O�?�ͽ}�Ÿz��������O.�=e�7 +Qg���G�n�А�_+��q�g�Ҁ328��&­�g�\t0�^�9� �3��LH'y�V�+Q<I��۹q�c��6f���t|�
��j>�-Ρ{�0m7C猊�u���e�e��ڴ�����2Ū>��}����e�n��%Z�@�u{���٫p���Z�b�r����s��uB
8Ɲ��U\�N����L�B�����ѭС��y{����d�r�����p�O����=�>�{�^7[44
;"�2Bb6��>c3�l�_�U� ϧ�IU�{�qW�8�*�1^�%8
N�^,�:�@�P���:<�I�ÿ��x�Vʇf�,�5��M`A�N��B)�vB�5Z��Ŭz)'ه\�,M���q}k��f�i�t�T,x B�E��$}�f
p�	�fkఋ�>�V=U��9�T ��6����m��f�#sp�i��\�� `�i��������;���n�p@����So�P�gy�q�˕ h]0-!���M�`�O鳟"�KC�h�V��!0�:�g;��R%����<qe#*@1J�|_��,��=�.�������4�D8sv�m6#��[�j|�gi���"E1Zφ�� u�D�����9^��8��g��7���/"]8�w�>.֠�kj���5c��ֺT�5n�)��t�L0j9�|^f!!��Q��;q�w}�м����d7]�<�'�Jal2�ө_�y�v-�X,1�ҁ��$ �n�����.V[��vS,�Q��+MX��G�B������n���Xo�iM�X�v!��!�e�v�쪳
1ƼÆ��KV���ʘ�w��n�^*�g���}�Z�x~�N��-+��Ow�БRp�;�J�"Lڟ_^x����p;>��N�%����n��|�<���*=��G��}iaaBc.u����bT�h�Z'O��x���"г�84�$5QY�j�\�W��4��J�tg
�����o)H�/���7U���}M�,M���s��.̢���VɦcU�"E*2��@�_�����r:�m�J*O��QM�I�M�ȫ#�l�eZ����<���	OrʱohbcIԐQa"K]P����{�ِqeo�:�4��)��F1e���poԻ1|��,�������:'�.��(��������aVDEc��"�74�A� ny!�KTJH�d�~�	`�(v�e�q�B���TJ����u��<�rp���"�S��c���i����N#v�R8K{Ŋ���,��(W+��ܢQբi�x��>#9'��C�oю��o쬎"AE���"��h��[�Xx����9��=���sU�������߃��7�!��a�t,�)`^
v��e�h9�+=ܵ�A3���y,}�H"�Y����&@��z0�2��)�`|(
�N���$kj>���0܀d���K�(JiY�T8�|ۿ��*ډq��MąF=���qbP�Ɏg?�{8擭OގP�-��NH���]V�0�/�0Xͼ�k��'�,J�=4*1̰�;�P�Fyr�s��p<|�T�@ŠDlo����w� <�d/XA��	S�u�_%l�K�u#���S����ޠ��T(�� [ɼ�jr- ǘ[�6��BjM���&x:�(E�NwR�i�؞)�W�i)���b����絵O3����j�n��|��B��m�ԝ�ěK&��N����B��t�Ŕg��-{NE�7�?���:�`�"�~�Һ��ܽ3�Y�g�D!GN)rZ-\���f�N4I�+,!�B�+6�'
��=H�A5�Mv�3T�YS'R
�5q[��M�y	��7<D+y_����Ze�E��/F^�#�x���k�8��E�3;�jϮ�}����p�[�W]���ח�Ћ�'"���.�)0~f�R���6L��rk��v�&�X�g�;�M��p�������X](���A��_�Ec��Cy%�%���P8耞��H��#\����*-�8�����~��6NTm�����2��g������ Am��eG�.SUSu{�F�㚦e���6��H&�ٍ��<����M� �RW�n�}����qL��d#0�v�����1��3f7�u����xn�k?�$!d
c',���,p��`ևE,�Ί��'�OѮ��<�JJ��=Fb�uL���9�.��)d%��'��Tc��H��Ɯ,b��|n�/��9���+I�@^w�a�·?n�z���d|�9�J���>{����u}?��@G�ڽ���A������YY�g9��GT��b7�w9�i�ti�|b�qwr{�n�3_�_��y��j�;v:
���B����)���f%�@���'��٢��]>I�u�?I��4d����Fp��W�q/sS��CX��d��ݔn�w�M�=�R�(;޾΢�˫"^6�m� ���Q�\�f���WFv�)s�^���6i�ԡ6�E��1q]�
k�����u.DX�k�`�U��1�����uT����;�kPr��F)��8vz�e��l{�0FS��� y�.zw�x�p	��i̟���r�#������{'��?U�/�/�Y�����f��<��Q�>��[T?��c���7Z"�=ϒ�J��Ioi`�����j둱�
'�Gڧ���fN(�;d�q�{��X���׺Z�ƌ]�5�Y��.Y����8}rU��ܶ�����t��C����oL����C6*��R��#�RL�N��x)��b��<�TJ ���d�+>ы��q�|%�v}�\Jt��ΰv�W���5��gM}\�Iovy���6��T�w�r��Ϯ�#��g��js�!��[�="kb8�|>�#kd���Z��.,?��s��JY���[�+�{qY*�2����e�1.���=�\Kp���5MO�hh�PO����!��t£��52�C�B�d�	��1r�	���?�ލ�u��5��~�V�.`h�/�(��ǹ��G����W�����i�{bwo�Zљ.� <�r>ш�R��$[�Q������f�H�������q������4�H#��7�rA�����#ܿ��}
���+S�;5*z��ҨN}��Ä��ƌ�w�l����+.���Z�{�9,_b��R)���g�T�2j!O�y��mopP
�����n��ֆ���
~�b��V:��=��0G�k��G�AEx�Ɍ%1�qͽ��fg�AD� ���/�>�SZ������3c��~]K5��<���cB�D������&�+�'h��|�.���"�h�Ͻ�@��t̀T������KI2)�H>��Tj�4W=�k�;���K�'/��a��E�>)C���k½$V1BI�o<������=WYk��Xq�0��w�圄�%�|8T�;Q�����"iH8+`�oj�4�*�;�BR�U�i��^@B��5�Ř�0��U�<ʄ���'�mG����a�_����QB߷p��(&kn��ڲ�|�A�z'jƝ�A��7�p��I����<����U���`pL��QMe[�HA���E�R�e��H[�������������:v�drJ�o?�"�w�dAI-WWŽ]|���Y�щ����^�SH�_;�3��wQ��O�`L��F�٪*o�봣 �j�!lW��A� M^vk$5�D5!��X(��W���e���SM���[M]mZ��c+<��T���R�hDb�~շ�!��M��x�'Y;nP3�7�ܾ�P�'���dcN�i�ww�ׅڙ���,�+� ��u\�?b8��s@��guU�3�c�js��ˢrr#X%Q��&ʴ5:ѷ���Kxpo�&#
�D���r�D����͚�{�4�"zv��YD˂~�-�l㇍��0"ÿ�:
��*���#_Â� ��ݫ�˽<q�t}V�.
c�1��W�@/Io ���;,^�A!<k^������*��v�xЎ� ������U�	-8AL������U�ʫ�l�p�����򭈑"����+8�I��Ў�b���F:��sy��^��oZq
/���9I����遲���#o���Z:Rl>և%B\�a%����H��f[@�N���Y*����]dPPvjK�"�md)q�?��9�8j��Zn{�Mt�>���O�#"9��/Ǵ=��W� Mٴfw�]��M�8���S.�-Y;��B����YG#j�Nߋ:h���a�Xt�x��4��f�c�zO�@��ּ���Ts^��tEp�fx����3�+�\Z��s��`Q�&��$p��<c�}��	��6PM�m?�*�o��@����T7�'(���e�s��콖d{�)���=��:Q�	�Ζ���q�w�	`��-�D�H�.F+�$+��ߴ��Q���h�t�k��e�p�$���s��n!��ʰ��.=����U�� �Wֻ� �Y�d
CT�W��)���u�)�?A�;���I/|L��A�����n�}�Q����1V�H+��^n���tS�]�W��G��$����t�bj�{�6��dB����/���LeEL9��v���%��w�ȏ���vn2tד���I��#���@�:�$]�=�	f;w�u���e�Z���D�N`(����l	!eن�u�v����uSBG{2�C�/,{�i�Eȅ1P���;�h
���~�e�F[ �:��S��VGw5U7�L��#Ȯ��}�]���'i�E�����%ה��:I�K��
�����)����{����+�z��d-$
�Ԙ��z�A�z�|��V��9T���䋈�*c�J4娎h[X�S����mIE���脺�P�����*�:�_K�����p'z5����=�7W�Ǝ]�e���w���Λ5\.	m����b�r��g�f�Hx%�g�w����<s5Tp�vL����<���;*}�E�78���:�9��݁Yيdsc��Tc�Cǭ	
�ۋ>�}H\}-����U���M��zG�{�[���1�ܡa�Ee5�jt�u��<H�Y�<��,fW	� � ���s�U�;�O1�1y�t�kZ�����1n����p'A�ʁ�Xg���.oܦ�R�� ��1����':,�������֌��*�y��me��!�|g'Mo��Z �e}�PĚׯ��T%	X����k��CV�M�\|�<�� �3��u݅A � �����-  ���46 (�h3�W�D���_N��0#jy��`ak�r��Z-���NA�4Ç��/�6�h���`�m�.�T��Dr|ǚ},'~";8����F��8!�x�c�x��MĞ�q��ڟ1$�(���Tꍆo@J�2�4�c�y����ZS�<����PoOx��)�M?7n�'�;��g��=�b�tVcH$��q4���4O�W ����wF�n�u�팿rt���D��x��O��#xA��8g�e9��i�w"y��飲1��(
��c�ݱ(��H�Ռq<"@�+�р�&A���S^?!�J��{D�^&v���1�yxŧ�U��m��ס�?��|Y`^�T�F*ff��y�g�32-ߧ������I�c��
c;m�"Ӆ�P�{�P����& SI�/�<Z!b�&2Ɯ@ +^I-p����߇��@�"��=gۛF~��2�q��iֈW�С9�  �G�A1� J.�>54��ú��Nq�~֢���*`�V¬_��ȃ��c��6��6�)��/�7�,[��!kMѓ��Q���$ �v�+�ǛY�V��'%�q��U:�li�ыKƆ���J<�2��sHx��:wW2���:J�t��N�z/�ᩜ�!O^��9���5�[��,�%���p�����DZ"�����,�����E��3)�`
�ő�}�6�P�>�Hl���o��c���[�.	C�Z��^q>l��Q�h�_x�i��������^Ҕ4n	�4�e�+�h��s��㘳�Ndh�J[�.��t������ �ܧ��x���~�
��y:���3y�ÿ���^�Nc{2T�����>�*��P�{I_�1�ڥ�'/�Vb���z��Ք*��kp��l���X=㢳ꐥ���H�:�'o�/�Ax���U%�=�9�F���R}yԵä�؄�Z��-�����8,00nI�[t�8�Ѣ���V#:Yu����j�?��B�~R�p5�2r�ccrz�#ZCi��툠��n�nɈL��ͨ�zf]�y9u����"�W�=j����T��>��(�
僯4�G��\G=˶W��6� �u�R9_�b�-g������H7�g���#)d*���$𺞳�	����S�t<**��
l%H��_Dm=E�KX��O>�v��0����z,m/�j�ͥt�i�ms	\�g����D0�蹲��Z���T��/^C�	U5^��)5��.0uy�m���� ub��ڣA���}�e��ۦӇ�ӛ9d� 1*A�A�ܷ����Fm�W�%�G[}݆ǉ���A U!W�&��Ñ�/��{��P���9CF�a� ���/�V�+�%��x��
Z	I�D�ѷXr��qej���54�ʫQL���$�UkF��Z]��Qgs��?���`����ג�V~cc��T���i�Ǽ�K�R<.�	��9{i���#+̊���ʎk�%�F"MGLa���HT`>�ZR�+�5X�,rb�86���Ch�0!�b��)������L!H6\����E�>�?_f���T.�4 �H�7x́Ϡ6�@B�#�~8�v*��2�?���/��bA�hG�5��H�x8@W�)�L"c>�5N�$�d�j:��t��ĄT�s��C��ѻ���5������z�¦�1�aFs�����(
q���eb"����n̜�["s�(+�o��p�j���֯΍�J�_�$���(`�e�Z�Y��<�x�欺L�)�I0T+r�s���a���.*L폻d8��fw<8�`&�������,�wb�=i`M�kh�(���c��#���/U��T��a �����娮�	��ݺ�=��%qx�dU���'����`�����I��S�E��_��Cf�+�b=/�%K���cw4&����5��zC�O�Yi^�|��iN�.�x�|1!��q+�uz�w%��@�ċG�c 8��I�@�TU�w�oi� �͢Ql����uЛ���:���-��Ѿ�v3�-����B��Ee���
;]L#w��N�1`�+�[3���ox�8�?��kw�����!��J|̬����<�
G+�Dm��\�.Pq|�� �l�TM�P�jg����tj+�3B��O��wk/�mmU�ؑuC���=�v��B��h�U�#�9Y�:���X�^�O���c<&$b�b�޻��z�]��}��v�ߠ�c�T�ꢇ�x���������0l<���(HXV���L^��D����u/:�5 �x�7Wu�����d)R3#��f���ؑ���v}-�R���k��	󣷔�.ݬ�q&�  V�Q9��&�bP}�ծ6��G�Υ�r��Gd�<o�h]�� �˜X�(^75�zR����H_���#GˁW%�CE�"����x�oh�Uzo��
`r���G��"��u�<�a(k���h^�YH	�5�f+ Ɍ��X��kO@����4؂�ѳ�D�Ĵ^m�k����(�\b�w�E��m`/A�?z����S���Py�x:8��2`�4�$��n��91.�,K�be!L\Y*^V���^M����2"͡KyHe_zm%�uƤ[4sE���5)z�n��D�
�P焥���+1r*0����C�\�@��OC
A@d/�qB��C�ex�	|:JSʞ���/��*Tǟ�Ú��X����Dx<�/rm����,�<��L����;���Z�Ҵ��G�GB��r��6_=�j��rZ���P��]��ZX�߃:�M�X����(J�C���c?�x�൲`��8b	�x�y'�� ^]&�E���9����5qZ�mD3�'�]݁�EH�U�2��A.r���3��G-�^��pM��ɈC�tEYƭ;�$ ��p�U5��>Tx�17 ����I1:�s����J�)|if`6�Z�NuQ���6}I�b�mTJ9��qԬsqMK�I���Yh=x�s��2����a�'��S��>a�q6r:I��5�9�CQQ=�v����n�F�C�6C(���6�OG��NҠ[��d���-^�2�ݍ�=W������-��������-�z=9��������+i��&B%��ѐ�M�_��+�#a��uC�(˛Cl_L�_2��t�=��_�O�3�W�эp95liO�g�[�����?�1��� f���R��5����C����B����j�T(��#PŃۇ�qݱ&�0�%�����"�;�Z�Q��������L}�az{3ۘ���"�4���7֎�-�?+�ю�����Yi��>P��Et�AL%;7'�K��t��|�AfwV^���E���N�V 6�O��. �qZ%.l��,r�@��!�V�o�X�/�G�����%c'������"Vbo-��I[`
�σ�����罣�M�`��{(o_�.��+���ΡR�Oy{�8\�n0ޖjF]�uK���������tNƷ��m�dn����LUW��g����E7�M��[f���PU%�\\��#�x'��dU�1+;h)�®�[!�A��c?����xɺ�M���}vU�3�c]Z�o�����K�?p���^������$oɠC��4��lw}(�3Ԫ{D���Q����ÕZ�s{�n��>d��䭠��x����]ɔŶG?�-^��E
�т��aڹnkN@�9��{u{���Uz���J6ȹX��i�W�9��6˄B�Lt�Hy��K4{ ���D*noF����~�!�.�]t�)�TA��$a��z�3��8�(Q����^�PuSH�${Ò����G��&�-��2>S�$��+�:J7Ȍ �g�>[1�e�nC]��/d˲��?B21�kRY�նE�-}B��4���7���:dɹ_�tZ {D��J��A��c�z�P8�Z��~3�,��(��ӎ�WZ�̼*��<C�&Fr�UQ"���"j�K}n��5�^#5�	��d�].�m��\Ĳ.N�uH�X:g�k����>��
j�j�1<?�I�|���O��8p���Qo�Y\G}�0�&�׭�F��!�;�=�����8��(���l��\&���y�p�?q]�a�/��tӎ����6m��J(������m����*���²a� @/8��o�����2�-k���3�6����5s�T�����4��y@I�v�Ja�/-�����K��+�s�3�Yll��h�؊��s��.�g���]������%f#(.��(G���-+�����U�7W6�o��2:̶�.t�^��#nō���ʩ�lw�^n�H��At_��nc~��ȤO�b_�e�14&�?���s�a�=����	�h�ܩ/Z: �O��c�ŭ�x���0�)��uT��Y��&��m�e:y�ft%Gۖ8~a�I�´��(G�+ۍ4�$� �,���6�v5KS�Y���w��1<6U�v����q+��j��ed[rF�{7�2���f�N���(���U���뱾�Z<��{��ΰ�vjwCC�@�T����j6�IM�<X�����H��|�~6�R����~�R�'}�������{��Hz�r^iT�y|���.�_�,�n|wۉ�d���W�U�Cr���f�]|\I
I��]=֮�q�!<�$&�r�i�i;�����.��7�ȗd� ���Z�I��(Ǜ�Q��æQ�Ϊ�Q�zs��1�|� �t����֨�5��i�$�\ ^ָ��jb����ڀр�Tjvt�?s%��A{���ԯ��H���Et*z^�~.x�ks���� �_!v�u����!H��g�T�k��#����8�ԽN�?H���&��90��Q��j|��Nb��������H�p&-������f&���/�3d�ϟ�A�fo�"HX<��<t�8 Wp�[|�ռ]0̳	�qaPU�E����9�BH��!{�<+�������d7�a92S-�	6kM�콴�����0�ȱڗ�+���6O]�jH��Ѿ�f�1#�B ��3ku7����֖Vέ���R��klq_*�M�hC&LPS:���M�¬c�p�A� �����S��n��<�f�ƥ��9�fS��ꖸ2Aā�̾|�ޡ_�k��,�/�X�8!�6>��a�m<u~��$�=g��C	ˇ��MEEb�ry-�N��p���b��	T��>����М�/I+����)?jH|U�P����2�|=d���L=ܕ�o`'�~��ؒ�nK�H���	 ��hjZ%�~r��&�[�<����A�h�R�:�H�!�����D���]�=�M��r
5Qg
m��-C�)�����@_No�[8c(����N��Т��W�,cz��d�1	^�/{�Ã'(�1c����ХN�c?q(�{��}]�����v�J����t��_0
ޏ��y�;���>"O�?7����GB}ԋt�S�g7!r!|y�ۧ��5���5��k-#�6oZI���9������%|ґn]�~��$O���ľ��t!�ކm���t��j�� ��s[-���^^P���ᤁT�)��{j�A�ŹZ�B��z�n�Xg�6�8��1���M����t�[�tSAG	M�͖>KEQ�.����)3{z�;2�>Jr�}����X��x�(�����W�k�?\f&R�����P4�&��/��R!�NT����7L�3�۟?�(�ek����+�R�ıo�YL"��J��Uj���"�#��T���/p���	����M�9�fi�9���9�H	}�P�T�4��k?>23K$���i# �O�6��T����DKu�&�.��vʍ�x�8�����>�2�e�o����TSD9$�f*^_�L�Tg ��!�����$�	~	� �	D���M�;F����*+�������1��KN��%_�"Y���~��献��Ng�X��~1�tv� �qȬT�ǂ�D����)=,�(ZⅱW����6��2D��`��L�\�X���K�u���Q��0 x~��0�|!OU������w�T���1�=�˛3p�̝�9 9(U�$�n���FP̿���V�zF���@�u�J�p�q�������G��3<��P�B�UF@T�(=�� ��X�y��ѓv�G"�.ݒ57ጭ�?�;9?ᆷ�o�z�`�7����W�'���gX}�f;۰�����\ҟK��z�TX�%[�"C�g�. p^8���{�R�9\����"J��]���T�s�|���wf$vi* {��;���2�����E�E��{ӏ�]����M�7_��d��E��o=��D�I��-ǎ%�#>f1� mk+¯F�SZ��~Y�+k���O�Q{�ۑ��ϵ����HJ��*���	��u��͘BkU|�\0�{�ޅiv���y+5�{���f������B���^�G���I�`���"R�ldX�" �/ַD`���H���u���}�2$�1q�2 yc��f�����ְ�>����̛�\g㭸.�'������Pp#�/���V:�C����t��cMe�	����K����JA�as�H��{�CP�o�p���p��c�bi�Yf�"�!�9	iP���J��T�>�-cp֑���<�'9m�aT�G {M���z8YK��a%�<j�/<~*�X���/ɪ{�]�A=��ʐ״~0���|��T!�EK�g <L�I҄���$�n��� ڱ��Ř���%�~-����+U�Y}U�4%�|Q�p��K*E�צKl�K[a����2h�w�g�*Fm���y\o�JäF�n6<�fXB��U�%�Z��I�ƨ��"N�S���LzB�)zb!���D��g^�Ȳ/��RiƬ����2 ]C��0+�a ��~W�L���5�fTO��R]%���P�谍� �N[�l�z,���D���4�]�-/�ӕ�K �k�����Q��9��a�f�%���d�B�yBc���yv�2˗s݇�I�IG��Zb�-"��^�8\F{��K|�G��&}����!�v9�d� L:�y���D���h��!1ԑ�OWEf\3Py|��"f��<ĥb��͝��t.\f�Rw{i�?sC�yH�T�P|��NjD�NI��C��ɷ��'�T��L��Y}n��e[]�X0�y!!��Ԋ�+k��XZ	o��!���΋����Rr���<���*���V�<����6RrN۷u}�)���G`������-˟(����č#�q�-��&��z�(nD!����Y@eOU&�Tgp���|�8uT�{R9�Ѫ�WBĊ�!>���_�,���d��5�?�u=�0�k�՟�/��Ν�d�� 4��[����"އ���'aw���-ƿ6p+���ҞZ�����a�k*�cY�h���^�1kB�����TQ�>�Ļ���e����G�J�6�1F�
C@'!�Qs�ɼ˦��ɍ�(�:B�W+ M�+����j�<����Q��@��Yfwm��kG�;R6!��q{���C��J�����AF��Q(�$
QL9	�E��=+
:�2"���'��%�EI�������y1���̿������9��x`����1+N���G�6�!�Pܘ�+"K�>@���4����'��K��\�,�6e�3�n�����@�%���#��$�t)ne�K�cO��l*N���]�Rb�Q���X�/<\�.jg�4U�7*�th�NFr�\F�ǌg֘t"0���o<C��7ӣ��"�1g��i�,tnV�.�g������07�W!���X��D�BfTvԮ4�2vI��;�<�f<7��q�i��i(�>,K³&m��;�+!⻁�d�a�c{x�V�{��Ln\� 2���-B�)f��}�-S�_�k���ݖ5rū�>�3oc*`���,�5�P�6������ڣZ�� {�=��M{�i�(�4��րX^��Gr��w���GM⌳N�[�;쉮ꇽO1IP]�_����ְ�T�]�MyI����+b�\_M����&p��k�W����cL��$�0�뫽=:�N��u-�p���ʟz\Ωю�D2�@�۹!d.C�2a�j,�)�ΐܜ��߂� Re7�@@FS���=#�n����p��u�� Y�Χ�<=e`G~�µ�M?qy/b��#�^(�����ԉ禩Rɋ����i�0����i{,C�� 2���j槃�A�������c�Q�oo�(�a gR�[�S/izBs��:N�5h�b���0�go#e9I:u�R��Kl�Q1��,ҹ
 [êpR+m2�ī�;N�i&� )o�5Glؙ�]�����G�Mፍy�&Y�M��N�y�����4�Df�u���
_p�Id��O�JL��s%2��T��iV/�rP �V\�#���B��+5E�,�����&�{����	���J٨1f:�;�^+�|_��G��~�����F�[�]{�?�;0[b���Z�7��sj�+6´�- ]L�5MP�Ar�`F4�&_�c�Y���&��Q#?ͧJ[�;��x��2�-"�7ځ>��JG��z�U�Ky=&���Ϸ,@s�>`g�hۘދ�o4Ja1PU����:�S9��'͖W#�^Q���V�x�1y�Kw\Ũ�vR�E�t��~u�d�n�{�>��(Fz�#bc�E9iD�t�9�nC�� ��ѹn,�8�v�cޱ�G5��B�Ԉ�Ͱ2���=�K������ڰ�_�= Be��_�?+d���YEt&�$J������/��P���o~sQOR�[DK��|�Ł"�WNZ�N��S���B���Z�a"�|�{^V-:��k(�?i�,�/O���]/g����E	�R^�Q4%�/�-ń���/$f�&�"}�O�V6h��}�8.&��l�!w��g�W�C�n�}� ��ͮ�R5�� ( ٥�@����@�7Y{X7_��6��4�h�k�ɦ(aZ����DV�P]n����#]o��ZZ�S�n�![������ϧ�0 \ v�;�����m��x4ߪI\<��;Fk�$/�V[v�w��S�����x��-�-�^X�� �n����
�d��<��Vj�+uL�
:�r�	�a`�������x/ eХjP�;n8�XyLRS���xI0�z���|VV���g�G�%��>�_V=��>����D�`̴b��S�/ih�8#��I_��=� +T�l�	O)��u�X��>�
��YN�G�m��g/d[4F�FR�餮����{�������o��~�]&�G/��M�+)����y5�����RA4p����r�3 ��&�������}-�S��ŝ,j�T{#�[G(JH��Ȗ<GP���61��K�jW��8���#jN�»^|�P�ԍ?*�3=����ܺ���~Z�V|i�|��!B��$�n{�F���ĭ�����0]0Õ ����%�,nr���N�����ٳ��,�����vX��:�}������bz����� ��3&�mSm�|�<��6$ēp�4�f�q|%��$�~���{Cs�N�Q�	�!�ZZKJ�$�+�W�h鹇dV&~����M�������������q��[�$�&k]3��C\�jȶ��^њ �#xe]د�%�l��\x���N��&~ڼ  �t˔]� �$ަVP�.��[�@�b$�On�Ec�컊���lTi̕T3�-���n��R������a6��i�1=)�)}���t�.��4���g$�KG�����1�2�Ӂ�H�H�!9p��6�st���D�/�y韟H0Y�ݡ|��m��2�}�����km�*����4)��ǝ~���bL�a1ih|�վ��.��yS��Ai��k#������!���g�XaW�W�j͈&�)���_�x��;t65eN����D��*��Σ�9�I�w��Mb�k�
'i<;!�4E��V5��O��N��~��IKq�@|aڪ�·���	Ća�./�)�.�x�Rۻ��Y�⡬��.�YAu�zu֋�����__�#ZD��'�)%�J����%	r�Y]�_~��m�!��v0BWE`S���w>�cF���\s}�)	C��-N��;���l�ӫ�Wr�\����+%�6��ci�<J�J=�ͦt��� ��fΝ�4�����������9� �jv|�)~1� j���Z]��I+��̮�і�ŽTI�D�41jA	?�D|����3JG6)HƳ�0�6ȥ$�ѮX�s���vB{��-W������N�7�.Y�?��h/�@F��˘�/�&�K��`̈́|{��|Z�kL�gc���8�̕*���|�9�f��=�>�I-��!2�J:�a�Pt'�X��
��ً�ⷊ19p���.���!���W�s�F�ԧ+��[�جl��sЊMv[n��%�j�r��<^|M�Ju�×��8|��`F�б�<����}�]��s~S��o>A8�tOY�9�</�()K9�t�	�f��e�+o�M��]�����V��i��D������\u��Tf�z箦�T��}>z�-���q	,`�?3��V첸�>K|����*�Ы�Ż�$�� ��R�J�j�`�Ψ�EeQ�)��@0�Ƚ�qd�\�\�C�瀘]M?h���}�`���R��k�i�Jm��_9	����8�	t��IRQP�U[��Cv��(��״q8�gHfL2�ѵ?}�q!�́��`#E���ˈ�r��a��0�d\�9j�hgwaE�"�q����P��10�~y�f-0��?�+NecbMJf�/��*���#w�I��jN�>�wk�R�����~�! 9�Z�����|��CT%xw:����?Y\�}�'\ɿ������'�k1��5��M.�������ZI|a�$.Q��f@	"�����������AE���vIZ�������o��yw%�����۞3�eE9�����0�^y�_x��k�x��SLe�#��4t���z�;0>�~rRNP�i��҂ rVK��T]�W�L�����t���|��!��[(��6={��U��pwG�m&�}��=9_�$�?��o8S����Y�����$�W+(���e�N��^��?�/�N���k^�?�c���nU'0^�.���B"�w��m3\�!^��r����tܪ,����d󐧀��!JX��b���p�bլ�K���^�I�.Maj���Lk=�?K�1��[jߘ�E������R��-\�}��B���Ȥ���\ĥ�װ���Ga�`N?F�Φ�	L�~�x�X$B��p�b��q�Sa���M����T+|E'��Ħݤ�/��pe��K"�zYg������hT�>ĉœ4���a�����/|x�����UJژ�a���I�
d�7�&br��n����y��.�m,�)P�>�Y|?.��"�H�����WǉI*xpA�!ڡ��lc��\�g�/f.�N�m��
T��J"�A�[ߩ!��xf��0�� �V�G��S��x��.��z�)H�UH���}6����#��S���bg�����l�'Hs��N5��
�SQ,��t|>�a�t�/�E����6E֡���薸�\be��n�+�i�i�d-�%Q%��0��1�"��c�֔9{�ገ	��\��վΧZ�o��#�jF���6O%2��(2��G��M~�)��,��s#�����fM@KEʕ�Q���akI�@����?�����WY���w��w��vU#Л�86���>4���dTF�ۇ�?09�m�=F���'T���:v�@8�,͸?gz�Ž�-k@N%��F�*�rTd�Jo�$�~o@�I�+�A �n��Fw��]�"�j��C��u���QA��I�gf���\�����Y� x��y��LgJp�hEEI��o��YS��i����$�� h��EU�\5��љ�eE+:���I��v�H��_��d����z(�����������-�3��{��7do��f�BA����2�]}��>m[D��w��c�h�`hw�*��u��l�2�1�B��@�?�{+��=����Pʚ��*: �E衷�im�J�1Z ���s�G�Ӻ�D�b��dZs���b��5h���چ�$�Ȳ.E0��C�g��C��K��>��x��"��%�Թ�x��g�l��na����}�
hu_�<���@r\fID���>�. <YUD;���P|Jnn!Eͧ|��E!�~ʊߨ�t�7*9���ee�b�,B�C�Ю4ڧK5�oҹ6�W�Z�}
�ݲ�������y�����Y�0T�N��m�/��0HH_q���_һ��.�L2��>z�\��
�<>8rj��S�')���z��B=�m�P�W,�[#�I��j���^����6�:}_qzXg�_gX}�dn>�Jw�v�������Q����!�Ѡ[��3Ns�H��5��-\E���孰1�+y�+ig�Cfb�)���ٹ-���;��QAatd�)>d����W��lUH������/r����E2̖B#NK�<d~�p ,l3HE�#Y�#�q]V�0sCU��2ƅ�7$����=��!���a���kH�N�/��&7�9h��'Z��"��OL:y���HO
T*a��"�¡#>���Q������=�}�HTIm�,���v���{���~����}K�f�(�����/;`c\ى%u�̣I�$C�yH*��`=����+��&H�M�:g�fb�y;LtI�!��7� ݶ�=$Q&�ΫQ�~#@����0�'[�~�[��K_���6��['�v�}������9q%6�A!x�fj^��V�W��o���W��Zȥ����T���Q`ؠ�(�ji�!E�dT��+��Bu�������!'-�z;G�.7�v#6�����H��Mo��CF��*��j���Cx�W[�'M:d:d9k
~�|�������I�Ri����XWmC�F��{5�=A���.?�c����	a/��M[I�����$�����G3�Zq1)�\ѧ������,�
��oFs� y��uԞQS_@-��ܓl���3@�Y��] ��1���4_m�H}I���y��%~�#��XN��y1�~b(Pfh��C�-p>����{'�{�)���J;��W�p���G�ϗ(�k`�t>��0=���O_6�i3hO�P�
��O(j�V�JNR�J{�3bwX�Ȏ��1�2	�P#�|�1H2�M��71�f��x��$�G$nz��Υ�����r<�/�^��4k<I9k�E�;
�FH����)��h��@��PMH劾ڊE-� ��K���Ru�*�`6���2r8ϸ�m�>Z��b�\E����ue���S���_�Q�eYfg���-�|��I��s1�(��p��	�Y�1_�9��7T׸9�Zl�l���%8�Z�U����G��ɐW}�k2�:���ױ��7��� o�z:!��w{�,k��~%��#?K$P'ղ�r���(]��1�7��?,}�^���w�ݵsa�A�~����:�_�7V>���칙�d
W�*�	��������5M��|Tħy@���0���'�x0������Jo����\��1v�	Ȳ&�_)6�A"&��A����e�yd<Vh.�;�8�9\2��t?�ׇ�Õ�Dh��h��iLf]���!G���B���H���wk_p�)O��:>Z!tJ����P�p�� �1A�f��M��bZjQ7t?�H���z�Oȕ��vq���Z8��
���{2�p��Ȗg?oBI��Fg�I���q^��4`{�*�1��/�Z�	,�@πm�k�8�g�DE�_!p�ē-Zd�z�ט��IȽ���a�a~�����Q6���ùH�/Zn/x�Ψ�il�̭\����|��Z�d��XF�O��a�"tFdJ5ư'�)�z9�t�'����Xh��ص�h�<[K*|@-��1���7e&59��%j�aǴ�U4}Zde��,IT(b�3!!պ6�|�e�u`��ԗw7f�U�iN1'�Pz�����˃Y�m�F�;�>Gq��
$��#4&����vPU��'ls���o8ί����9�=��ڱ( {:,�7�����3�#ǍT��[++:�*eC*�}//�׆L[@ַU�]xK���)7Bh�CL��U�� ���}�r���Od���)��-������]�<�~K���� ��A[�?��9Cd�R�����x��y�m"��0���Θ_b�y��6n��X�.:�Y���9�e�QB�ӋH�en#0�C�,��;�"�Ț#)��57�q�;D+P{Ew^�h�@�����kK�ȹ��s��R��E�o���S=v��u3kR��،2�XXϯE��Y�Ҩy�$լ��(L�������.�U�7xy"��h��]�e�;�,�o�;���l8l,9�`�X�vD��7)�R ��V�W9�s�?S^n�����!�`p�e����(ŏs::C�V�+nR�����&�)�}�K/|����Gȃ�aY�2|t65�ƥ!��Y6�����޼���{m��(��R�P�=��Vލo��p��T����8��$���b:�:ẻH�9s�};L����M�=�fVb
�q�ĭ��mn�\�&n\r��y�\���(�fB�K����Ȭ���X���u��?:ˢsmR��ClĊ��@,>Mم P�CɽEs�2}�NJe�9ł�)�M���w[�`�]��	�yz{�"�\uz��Z`�Ch����i�p�cu{�5�~��#�\�X�X��Qi&Q�N�S�Zكk�E�
Z`�עph�a�i�bM���=�6UQ�����(�p�����4��i#Sj&n��äB�4�v41�'S����Al_c��$�A���[E���C������=��VZD���?#�����"�%	(��e�&c�T�j�%��Q**W��6��m>Xw(�x
d\"q1�;��}�����W���q�8NC��������뀫A����H����L��M���C.E^%�p!�5D�(�u!���Ә�C|,o�tf'�jCT���vP��E�t5�(�-�f%n��/��񃾤��U�|Q3��p��M5�JV_͹�s��mG�痝��ܼ`�\Rd���=l1��*J��,Uy����1���-fRiQ��EvGs<#
��/1)tꆌy���|t��S���[�6v��y+�A����n,-�r�P�$�Ƅo��6�V��r���\���o�򉍾D��PPL�z5��D �fpw��g�v�$l�|D�ee)W���
��H���);s�='��A�&gd�����1@fe�v�=mب@T(��ɖ����ϗ��d&6Af�Ԉ��Z��l՟��	j�E�4�2K�!;�����d�c�>�Bf��a����u�cA`w��g�p�Q�]���c/�)�X��5�r�hVE��#mU�V��F�;�����*rp�����{�%\���%�F��XO�D:qu��-�^ȹ�����@iy�0��#���<�Ħ�f��as ����d ��/P�/Y��RD%Rx�Z'$;UG>H��х��]Md�1l=�aޖN�0:D�!�o�E7���΁��n�K�~O@E�W�3y'J'�x@���W��΂�$�O���O���R&����I���n�[h��{]��!�EP�ȓ��.p�|QqT�i��1j�@��u�gyX0��,�Q�E���z]BmE�8��È����~[�H��7�<Dƞt��!]d+{hĆ�-$��շ;ݞH��ҳ�d�)D��D�م��o̹<��h��60�H�t$ �[���z�7*6ȯ���v#�����Y[�]QvD��\UrxÌ8"�Q>�j[;��R��h��m���*������*�g�����Yt f����V��$�Z��Q8�� �n��|�DjSv���Xu�v�<!���]s��5[����h����@Դ��ژ��܋�C��m��e�>�6�3W�]y,P�H���.<bR'�U��XިAq��1��{r�{&L��Eb'���3��H��U� �$B(D/�����G��`VKu�vL�@�d��ڶ�eէ3�v�l���&�ٵr���s��*�D'6[	C���(H|��v��ǝL�q�@=/B��v		��|�ی\�\���y�?��T�Jax�^�b��c����t��Ɓ�Y�&�)���w����J��q�w�|����nX�ٲ�L,1A�[�7�9�۹�ߎ�t���k��!�3BMl�KeY��e3�TY".ȹ�KA������{G,��[�qƦC����4'��#���`��G�e�.��Ƈ�R��؃�XTjI'�a�'Psw/�4*n�uEI|0�3V��>gЩX�S�xh��z�d,(�w��]��I9�`�,�N��p$&�n���*��?�(׶��n$
JZ	n�r[�"�����j�/m��X�n�>�(jD���V���R3��Ic .w<v.\`LG�å� ���ߴ�tk"K��򍯣�N�X�UW�mJ"�����������nn��_�ķa�\u<c�.NҺ&6�}���z�� )���kHH����Hzl�%��� ��X�)�M��A�U�er����g	�UM�rjC��M�B��?�#/�_ً)��	�p�JQ2E�<��'�f����y6$Y�D�=-F��3!Mh/�H��b�%#�i�0�efB!tH_��c��t�k���=2jl���vy���g^yZ"=�s��EdF��09I��v����e��bY=���������Z܀����4q*�bՂ�2�b�]�0�X����u���Ay�,:�j��L�y�<����d"�%��LiĂ�iƊ@�i�KOY菇�m��
N�vk\AH��sg�*�qHS�٭pY9�� �4�[��x��s�=�*�ߪRrgl�c�|��ɿ
7?�����:�u0h��*��~��o�JH�b�f����R�`Nad�˰�Fv��d�＇���B�ju�Zr,��v &4&;��F���V^�F���V���BX"��D������1nBF��F���'��_y7Ҩi���e�k��b&�)��`2�������Yr�sr"���q�m7i�9R����xK�I.�p�$���`z"Y�j�7+"�תcF��:�ș��]�kQ����-L�N�/Ӝ�^-kJ6��ߣӄ��4�{�<�WC�9r�-�Ay�k�o�<ٺ���ҁ0>prF����7��ǉ.��c~��Rh�	�Vt�1
C�ʼ�ӻ��C����]Ɋ7g�A�v
��8��6R��c�k{0�x^���k���s��uׅ�魰|!k�����t�ߙ?R9�&9�\�$���h겍�q�|��NA-:���[-��,<�/ω�ٻ|�K����P������4�\g�g��6���%�=�c��#�#uUl�Y/��`���n�K���H��(c(I�w@sX�B�/��1yl8i~����xUO5t��9�-�M�؛�괗�����?�+A�񢕇�r��>��Ce:x#��ɥ�|�d�=�=x�\��Ƭ�[�!l��P����>p6#"�?��9��M����ͷC��mb�"W�p������JXC.��Ӣ��mƨ��I)�Q|���U��j��^���|�b�<	����{����gfI�'��|�|�9 ��h<>׃),2�V�ȃӹ�ڀ�h��B�p�����ⴊ%�b�ju������=l�
	1 �1�;h�'�k���?�s�>m},;4������6~L\t�Ӊ�'���nKy
m�����}����,,���fal���a��3sK�4�p	��J�X
���m$���3�M�d��0�� ��9��CZ3����ך�5�rf�|��qKe�5����jK$V��I�N�`��\���8��uʾ�g�l�ڶ�ݏfq����l��S{���0�4>����;W}HdC.O��Td�����Zmb\J�=a��	��dk�OGvbMv:Hw֚,�g��V�_� 0�4�B��d�ѢY\e�h!_uWD�R�F�ð�.�n����0�(���8���^Y�B�U�5�r���-V?���IS���6�ߦR32����_�Ɇ���܆���dS5r�E8�Sp����b1�]��R:")	���g��I<����_���u�A�����*E�:*ua���R[���<��=���>��{��~`����^0��F��󤏌jvD�� F�+����ۆίY���GDǣ�dA�l��k8?j����*7���Lp]4�����x����(@�\��<�x����bp*q�w�WC��awZ���hf�������fc�ƈ �G�&H��u��J  X��I���QΓ�x[9O��kZ��_/�2K��X��!��e�}�p�Ӵ|z��w��Ƅ�%�CsNa��@��-����7��~Cf1��xx�)��={�jm�Q�Pa�	��v�D��W���� ���r`+�U��(]���'��Y�ܥ�����P�-g_,�{ݦ+��{RI����B�Qj=�r��5n�#�'��~�*!ΛCi�*���F�|q��S�dqw6@�|�+k�w��jqE�'J�P��z6�T� ^�u󹑄[��u�~-��d�/�%��v����w�PI}�S4/��]��z���;����S]��K'�.P��3BD��^�cT�G��t$�$QYS�Tjd�.;�2yv�u'�hb��	7ť�r����@9��<�b�z�!{pL�����щ	��^�T�>h{�C�H|��(/�5S��H��+���2P��t�jh<Ó̻�(�F�h�^��b?RX�?��V��H?Dw�W�ҬRLRH�hM�N@{������:�&hB��]�3�*}U���p�b}�*�d�D�`t��	7@zc@�����([e�ɕN�ت�yI���U8�t�v��5�#�S����E�,|=qO�tU~��W�1����5��絭��
P�.cm�%@�3G%R�L�' 5�������8Q�U6u���<����AF��p��WK�G"�G{�N��rhn���˖$'���X��b����}v1�9Ia�ݓ�x�U��T� �t���0Ɇ �^}�y���{P��}��{(��~3���P\Xh
ݕl�sg�~���$J�ir�����DD�)�:ܦe(�j�д�+�y=|~���lߺ�"����p8�5q��*[�/�lq_G�o|���M�W�~����
yb���[�}��PbFC^	���DC���>yAڻT�<c�z�5H�.KZI��z���=aXt5H:�����婊^��Z��; �N��^if(bLT}��&]	@	�h"����&ܭo~5�U�j,+���`��Z[̇��{(%A�C��tX,�;��z����y�ɽ@ u~�=V3�e)�$&8%�D2��^�����|�t�\��7� ��Qc ��s5~����n��%)�R���Fo#�SG?��L;�1/8˙��~N3�u��F�MUi~���`],9F���˷�F�<"b����� �u�Uv ��X9,�Vh��Qm������S2>8g�[�Wz	C�FC�M/}V帟������a5b���(��(R��]��f9ˆ;���2ێک��Ls:���H<:�D?$,b�Px[(��i��^õ���ޭ�MX!�#�0��o�"f��n���ȩ^���,Կr�l�wG�YfW���`B�����$������t%Ox8x�z�W�2�а�k�E���^%F�@�P+���E��ɭ���g�����w*��#��rv<5Ȅ��u4ڒ���,��F; j�����Ĩ�M�R�V@�)�&@S�Y����wtwB@����ꖖ�H�S$��+K �W��R^*��~��_XS��\}h�kvnd6�C��ՠɴ/V�gM�D�H1��'#y���0[�j��"�H������t��e������)�"Hѵl�h�^�=�-~]s�Jƚ.��KR�h��ō?�b93�Ā������bo�6g�(Y��N�
�A�� 3qߛsI<��D�C9�v�ů��;c�r�QKs���z������P|e��4Y敃C>Q��*l��p"����2綇�����8؉�����0�w/`҉K9K#���d'%@���\���6�U��&�u7Nb�	�ɈK��v�^k����Ρp������XA4�]��x�J�
�(2�}��&Iް�	�R��TƱ���Lb��׵$q�����#��潉=fȴ��������}��P�K��SF����˙F6R� ��ᑝX-"~�@�H��Z�]��7T�t�%AL0E�d�E8�}��(jhM���bq��:�e�>�Љ2�����[�k(Iu��E�j���8A,��K�L��t�!��Q�V��8��ǰq�N��t�󅀯+B�>  Xdz#<rH�~��tg���.o�	�" ��ű�;��r� �s�E[J� @�������&K��QI��֙Ӹ�5�G��|� ��Y���	v��,�8��9xW���;]���Q�C]�IGa��}K?�;Y��j��c�Z2��qŮ�2�u����+.���cO���[8P���w(.�X"���{��ώы�*�a���\��|ސ�jA�QT�x�j�$�.�k�]�t���<G���-����>?���Xv+�,��=w��76�'^��_��q@�e|8��ۚ����O,�_	L���T+�
�WW������\/�� �^�㙄F������H��䧞p���i,�彅�Z#��n�վ�e[qn� >���4�6�}�<�o�L�G:z	��H������	Er�OG0���@I�^g vM�w�m<Ke6�Tq���,�̱X�K�VK4���m�B��6���nq�����!8&)ǃ���#J�( �(ҧ()>�i��/&M��F���nγ��WI������/� X�}!.�"���;�زɦ-Ie__�z�-b�*IWDw3��!6��U��E��w	�|䓘����Xo���4����C�7U+:?���M�,8�.g����r���S���y�פ����h*g{�D�"�a���(�Zi���p/7�O
�N^&���)!6�ߚ���mT~BR35�e7��g�m0�~Ͽ��5���%L�n�O�a�ʴi�~s��d�l5XH�_���iM�{�{�O��@�}M=�9��a:�XNؼ�n�ހ�=��N�FkƐۧ�~o5.�4�J}�"z�췤��ɹҶ�d�.��8hi��W�&y��L��SZk?�6l����&���I���ù"��j�꿆�
�@̪�V��H[~X2;
���u�e�t��=N��z���(�~@�Οfԓ�o(����4)�<���cv�R� �������������fP�Z��ղ�^�]Bl\A�+�B��(ʬ�9�$l��{Z�M.�8͗��Gt{���#!>H�+i�`��5���W����*�h�Ƒ95��M��7ذ�/�a<o������$�����^"p��4�(uH�ur��=>����p�ϟ�i���_�;mI��"����,cz��+5F�@,�\��������~���.4L8�ұ�Wh`'#}��=��+�Rw���y�U9܏^�h�v�w-������Q�S[z!��<�0F�n�|�ݚ|�����.�Y����]��̲��{s��?_��M'��lp�!l�^���Xo_f���>������H�3�-|0�Y�`J�������mu�-
]�b�f����M���wKu�ƞc���CH�+��V=��QUw~�/�p͓�ͫ�$2��7����(V�|ᅸB?���\!�%�gIϯ6��Y��^�Ruy�N����	`�_0y����U����;���-D���������GM2�p�OFK��I�
��*_8�y	b�-�K]�im��Ue�{^ɕ�y�<���.�A�O(W��	�/&�,o�aCz�vt��BfЁ��]�wT�6j��?E�X��}�!�_�L0g�&8(V����|5�ruAk��Ll::0N���1:z?�c���xNT�k�4��y�Xx�T�"n��8����M,=���aD+?&4���i������ԇ�Y��Aoy^Q��
���z���^���r�Q= ���4� ���?7��^c!���3p�Xt���d@Х�X>�#ҠF��zU�{�ܦ[q���Ճ 9k���/=S�>9�%�&��o�q)͜=W�0xq'���l�c��+7ޔ�=��5��HQ����*c�4�Z���
�l)ػY����*�+tv����Q�p Ֆ�������)"��{�r��Z�Q������U<߈�TY�J'���>w4$�z�?�IO�����`�T�`_���΋)�39�yW-�zy�V�v��f�8�i
b���_���{��[��,iD�w>2Z]Ϊ���P��79�x��A��1S�"}
@N�w���`eTc���3�"�D����W���h�������B@��Wm���^LLSB���21��ɖ�Cq�N�����k�yŒ@t����<�*$���W]
6����^si����kC;�C�.�K��ޠ8$��l�)-Z�r�vV���ʈ���8�����o�K�cF��_߁��:�r�j��Y�>�ǼT��~T�%��mU��P�GFΩb��� C2�ۮM)��L�,�.� S�*��W�1z(E"�[d|�:��Zc��� ܔ�ޚm��Ge��7����ST%h�1�ݚ�ўXV�oc�l�W4q[-���󨯖�9��}��ď���s&�֩�xW��ñ4J�*�'��,�2#��S���d���P�=$zT�R��	����j��M:�������q�U>P��oϑ��U�'�Gd��av��vj��Ʌ6�z3]�i�s�d�k�{g�� an���2��5n��*"L�����ȗ4O�9YW��MG�|�'��>�/{�V{B[����	��w�uF��\]壀si!1����ae��b�z��Eƭ�
9`�.Y��K1й򁕈��4��/|���G�p+�#�gc�����bg�w��R�n�M'�!�"��{���2��`u!��B���kd��T)�՞#���`"��Q$<ĕ�Lߗ��n���q���	�B&��\o ������*b��E�-�pj���"R����5�XZ`�!�tm��*J�λ�tXР8�9�m�2��ܳ�gu�uК�azž/�/�nn�>��+�:̨����47�z/�B�<YJ�`��<Y~7���\V���J�`��<G��O���c��j{ʱr(�:L�ק��6ć��U�i���F��-�[ut3WԮC���)�eouh�i���-�!�zE`�nG$���X�yE<^bY渳+�*�uW�	�~�&
w�.,̢2S�\^��U�[�N�5�1��i�T��-��>a6w~��\�������M'"D�)�M")�	��7��u�6�BQ���1��Zf�� �|�n�D�&�V����KW�tl=%!���u�&��9sN���c��<=�
=�G2��WT$$�HFD��|�*�Ț���Gc���ѷ�b�}��ɾ7����&��ek�ְ�CG9K��R��_���&�I7�Y���V,�dr{ʜ(�TZ����M�k[�7���y�f�2��LD��h���$H;���w�.d�55�ܵ��f*X���{^;�
;�a�A-K	׬Ħ�}��F��_{<�K.[�h�B��~8-��t���gsAr����ָ�­wPS�%:�p*"-����d���/���JϚ5|��U��n��R��?҃8�k���<��r��Y(�[yBi��F���p�Ud__WA��wN�:�8�pb�ٸd��Zbk*)�o�¡��s�`RT��_0�_��!�!}H���q%Mc��[�F�}.���s��s,?�h2��)�.�+Ga}�=��L��F���ۅ\�~�I����(�gT���ꮻ~�e�쥣\'�<`�r���*��s�O�D���<溞k\�kk�F�¿ET���E�:�ç��If`�3AtMg~�q>��P�V/��_�!�Uk1q���:
E'��W��?�ү��A���U���5.�W}�9*�����ܼtZ��k��;����/��������l�[�pٙ���qS��祸�yv�x�O�5�A��z��S�>�(kh]�a��N@v�OL-D��8�ft��)��p����D���A�C�ƈ^Wn`-\�0*Z�`j�S�'�?lG"X�G+&�&�)���S5Z�Cv�B��N�{��ө�4��ZWF��BbE�>�N�8��4���u/؞M����gP�kV�G�������]}=Rx��F����I�g['�D�C�{	yK�\G/a�>������`�T�?�u~Ԏ�Y�Ʋ���>/�<�J�cH��(¤��wFL��ޘ(݃���w[B@؀�y?�Ws���_�s�Yt��C�M:��vhҌ_=QQ��E���wn�$ȧ���=�>V�4��\=���)j�oe���5"s+E��]���؈��l]�Yu����m��H�����j� �1��~[c\M<@q	�y���^-���be��ƪ_��ɓ�����tZ��9��I�����~����t�1��inP-��\�Q2�|z݀��uQ�Q�T��N*� B����߰�Ps-XPX��bL�^0�ew)�I?�ȯ��F #aEk^��J��<��U�A!�+j��=��A{TD6�>����~�(ȅ,�9��s�	Pp��x�9�t�.��%���R9����P&Ǥ+���=
O�g�r"��rU�%��� ��F��t��T-�&�ϨT_�[�q���Čy�sh��j� 2��po�*����)�8�Vb�6x-"�]�U@K�P�j\�$��@k&Ԥ���;S�V�2�i��'C��w �e��	�F���_/��)An��I���*q"aQ�����t2M��(�d��Go�H7��)�l�iI�H���44 �	)L�vl51�~�*L�6��p��I��0���7L�P� �7;��7���6Y�v���Jł�gm4tU6�Ц���_U���1�!��߉�Q9��
�0�X^��(�:1���eGO&����r�8W�&�$"fL#�\y��z�.��A�:�H�Y5�ʖ	-���t�2u�]!��_�5t2��?� [`8Bܥ���cw�H��i��K�
vT�y����G?\���M��Z��*�U|� �g���/6��[�ZO�:l|�]��`*��.C�DN�K^�W��ux5	�gF[�ƙ"�w� �<��t~b?�$]�y�'gy�YR��	p�՛�B���=V���+'`�k(re��[Iٝ�7���o�Q�W	�igz���>�"�V���UIϯ�*��g*X&����!�!���2���ë�*��!K��|R�⢞V�i�!�Q�����@|]p���,#���/��]m4Vs-�m�c����1�S��f�>x�-^�{^��x�Җr�6v�+������Vd���H�����襾T���X��Ӷ�>���e[���9�#�(�]�mCKMFz�Q��ݫcjVqM�\���ּ�}8Q��`�X�G'<�@]����+[��Aw qn�ES�P��=/�?;�|�Z��|�m8�9�Ϸ5��9@7d��C�yb��S�Ot� ���WM�=���W޻��{}9O�dc��CB��\��C��Ș8֣H�c���r����-_� ����&���u����߻��8r�cXF�?�_�V�bϒ.PfK�Z����8r(��e��~�B�^���K*qv\)GCP4���y0?�u�vz��7n>Z����a���|������kg$��F�-���g@�:��'`�+|���9�<R4��h��s5!���5kGI����������Y��'��gUF�_�����;�7�XuJ>�\`=D�h>~�i6�1���`��cA�t'7�ְ����O�e,'~/�F���ҟ(�&�XX�	��,���q�:i�-�;��94�������A������!|1J�(��4:q�⯰,�x����-N����&[J������r��3�|��*m��<k�ln�'�Π�'�U�����5�2�"O�؟U:�q�j�Ĳ�6���YE-�IJ؇�KX}4m��2�}��˄'�(z�$wʮ�4*��nGO�y�=a22��ިA:�p%k���R��xxP���>�!N�aY�A���KS�P4ag1����k��5 (�`X��;�*(�a@P����Mm�rvP�Ʃo"�iaHS�},+���֦�L/2W��a1;��d�ξ
��1u09a�"1��hJj/��0ʤ���y��{u�ȇQqE�iK��-�b�Q�8��jw��,u���b�9K�̨�k�M�e4��fD�z6�ծ�5�����*����ę�9��|6��@ٛ�ǐ�;�;���~�����+�����>]��Ge�� ��L�59ƿ������<ƥ3�k�y���!�;�m�}ӻH�|Ey꾤�)V�2�E#��Ԭ^ݴ��'��7�m�@yP�(H R�O���p�;βܬ��b���gd�����/f��C��	W����}��轟�:_K%�]]7����ԖW�X�˝�����"� ���O��[J]���w+6��J3��t.�&:{�4�9�?|����J(�c��ֆ
�#p߫t�j��{�)���_0�6Q/�T�v�r��WҚ2�x�;MT^7%yF�,7�'E�el�!�N�7U|���I[�O{r�;�5{���zs���0�,���m�X�$���P�f���✃��N=�x���U�����}�V�A��k.�Ǽpv"Eӊ0�x�@^��dǠ0�K��vP_��&�������u�C�:���9��߲�xӿ~]n�E�#$��䙠[}ʝ���2'���+f�T��T�$.|���0Y9��h���F2��)E���޸��bR'M�R�Sp�1ڗ�YfL�9��f�TC*�(�	[[>F�%�@����*��Qy�7v �rE���Z����w�����Q�J����HU/V����X^��mQ�_c��X��nb�S�:�����Ϟ=�����M}�dI���J:j:`��{�g�}�Ug�8)+@��nU��k�Y�F-�6��S'-p� p��(j�S�3�S��O�J���/f�`|�-�?���\�����o�X�=�+i=) j ���t�i���f7mI�j-�Jf�S� l����X˽5@�rVh�Ġ:�ݿA�dv;=�OQ��X�5���?d��{m��l?�問Ի\��Q���t�)��$�Qye ��3��e%�=d������14u�L�}��^�j~���G����s���1��D7���`x�� ��l�9���3QG�x��?4�H�����Ɂ��Q�{����м��"%���,��,��xsZ�ո"�~RK���?�ɂ˃�5��ԋ�e����1^�@W��ӝ��v	Wd����H<l��P#��a�6)[� h:�uu~؋������0"]�x������ ��2
��򶖱>��8X<	ʕDWO�pO7оl����Q�So8�Yfs���h"�n*�H�x�:d�tI��Ge6�a�JYgIF�2X'4��'�<N��Q$y޴E�6.� .�Z-V0��Z� ~*���\�R�>
S�_�!uk}	ޠju��7���;`����W7�����ZH3Z�튑��_�$��<���'b?����6[/�ޥ��j����N��<���h�g����ݔ E��#!b&��6�6����F����S�~=՘i,�D0U��$D�k�EJ�I9��D���n��x+@�6�Á2�?z�T��0BK+�� �S�򬹯	$3� �ZF�x[<ix�0X_��A��M+�{$�!:l_jَ�M��� <�O����^�ݿ��2Jjx��	U��������w�?������d�C[?B��!��d^��s��Xd�u�����2�Xo��T�o�����b���y*�sٻ:��`�ݖk�� ��9:��xd�Gy�-��G���&�$�|\
��tp�;m��J��-�Ě�ůQ���+�p=�bH�[Ԍ���w�)��Y3��8���"��1,�Ɋ�7����/���9������7܅��H�1	!Q���G��qЉ>��3��te��ؐ~P�L�����HaU�Z@'}�ߢ��Q�X�b��x�Q>��.I�.H}El��*adsxq�0�V��@�u%z��R�C��#���H@��i!�M�5y��E�qUM�Z��ᨷbX 0K=�R \�
�E�8���:�:T��6�(Z���$�n4�[��3�%�&p���I���5^M�B5�_w0�*��x�����8�q���=*���"+Ku"�Ȩ���}�>�v���я7�
����%�!����r+eC�#[H�>��P۩������	%ٍ9ftL���`����?;��QD��X��>�9��/����QC�G#K��'����4��������2�"�4���&��Q~y��"~&g�K�C�a�6=��|-��E,O6�$<]��6�����ʖmb����Sc�6�P�5��a