��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�����uK~YSokj�&�9ȼ�P������şd�rU�gb�nEg��e��`�"9H�bLr?\�̩���hVM��U������v�u�<X�yvX	 Y��B����נOb����J һ�0��@N�L��7�W9�3pf=rT`YU�e؉4�*�q�\4��ʪZ�~D�����ӘFy��P�1�ɂa)'��0�;&�@�*��,��<��G_��0ө�����ܞ�$�Zl�cw�G�V�^�����)��%�AC�˖���;��' \e�n��/��f�	v3��7��:���9D�
�2��T��������r��8`�fwl�R�b4 ����Zr��+F�\|ZN��]1���t _������,�+zZe���D���?�}v���?绤��A@��86,7�o�>�~����N�p��ԑ�I���U�|M�+���ɨ�)�eD����H͠.�j���l����;0~d���������QRrw�>-�
J�\9JB��|�D�r�푸2C�#��������L��Ќ��l�fA"���X�;��9e����uAW!ad6uR����,~O�U�
�?���8駢��''���5�L ��J�S�߷��{�$�S�O� NԚQ�k�,τ��W# _��ב����`(��ʞ�W��z�@d$��`*��1���۲�q�l<Y�R�0��AS�fs��X,�m��ٮ��=�����[�g��*����TS/.��F0ه��ƌ_*��O���<w�O�s �e~��������`c�/�r��v4D>�{)��Jع��Bf��3��څ�$�����$a�q�H�-}	@]m6�%]-�>n6	�����
�ɍS��$I���(G �ɄZS�04�ٜ*w��������bG�<[�Q�)Ӷ���ZA���{���siW,���xOY;*���?�Y2:�W<*�ؓ�*3}���X��R	͔��#'�l�i5�M���>���KCѰB���*��𺂄��'	�{��J%�ųy��E�W+�?!q�����@����yZb��>�����P7^)��\��m��ޤ���%`};�a��ɰP����;n��4>ag*D$�ە�՛s9�E}�M��i�s���*K�v8�ѩ.���nC��^f��mቼ�����b����
��Er}��b3�5O�NN%�:���N��������2������������j��+*�(>$�a:d-�Zoq�j�.u4����89x�W�Z�����Ta���T�ᫀ���Ҋ�]�˗�|�s������O�q���8�	��)��y�X� ��?̃�(�h5����_�>E���\[��]�$"���b>EI�s9��j-�R� ���y�iߒ��eR�<i����_
C�1p �2=���m����D�<O���|e���am�^�?�9��+w�M��	��ܓ;�*��a���=*b��図��0m+(��,�v�~ԊW�~Q�$��އ�)#TA���� �6X�%1����$���H�L��ȡ֘v+,��.)����--MQ��i�&��F��g>��W=�U�!����]��He��T��=lGg�WX�Eżۘ���Ӫ�1pM����|h�_�
I�.�&W�����ɉD�{�]�2�i2>J�rGU�^��O,�MӾ���҈���TP2��@
�����ߥ�[����d	�Z�GE�m��T&���*;�9n5���-�ݕ����]�m<��v/���A'�䥤=��O�ݜ(�T	�1Ǒ�Qmyso�� ��T5Hl�y^���\h-�SVޖ�\�_����O��*B|�r WI�*�b�����|��0��j4YH�_.��!v�>��|�RƮrO�IxO�$!>٪�
%�윭��ׄ}�B�I�@��M5-�7��#4�2�r���>�0V�d�"�>*���W;fȳ������W������&ÎT��8|@����)��b�Zb?�q�`x������a�a]o]���Y��&}0����.�4�|BN�pR!yS,�xOQ�Zz�����}'�X��-7�"ǆ��
��*�ɂh)V��7�j8ؗ����Q�ډr�+e˨M>�Gy�,��qTa�f��}��{�s�	�4�����/��.Uۑk�����F#�M(�!�M'8�Vz��(5�F�c��l����
t��Y�s��܍���|ˬ: 1��9�E��[0��qM_��d�"�j.�
#�wA����$4guj�@9d����R+�u��F@`l����l���zY^���W�WvW�@�L`��-(_��:~~׍�ޘJYK��nu=���I���H�*Q��'ŗŔ������Fq.g�P���������
 Q��)�+�)��l&Ws��ݜ��C;��˂�C
/�?��6?9�,���N$�>��#�CF{f�Τ%�s�5����B�bw��.i�c2F�k!����f������8�<�s����Q	^���Y4;�ε��g�#���B�4м��ă��U���]�TB�Ȗ����+�Ó�Ќ����^��\�%�
�.W4�5\��\�� k�����f��Cfbq��tS~�.�]�}5D$
��;�$#�6>�"5�f�x�\éo����-��A��_��Ci8xʑObԤc�Ă��ecT�/��!����^b���Bs��	u��(��[c+<��m��;KH�^^:Mnn�;��^Z+SD��,��49I說4*O���ϻDJ��A�D�e�<O)M���T $�5&�@8�Ī]��^t\���-5�	�¶�vU�R�V;��	��F!��_��f'YM��R��� da�	�oT��!f���"p�w���^�������Xg��U������j����^���v�Ch�3�]�e� r^��Z(32@�59���R�ZSo̊�N���{�������!1�ʑ�7<�c�]�v��٪�o߂��i��.��>�C�ן���̢Hv�R�J4Ȩ>$�F�!~(K�P�"��}���;���h��a��ѝ�!Ө9$�1�����
�"�H�:��7�S����R a�n����;��eH������v�?S��|��m����#�_��?l+���8	tH"V���g?��E����p#0,i|�\�AF�v8s���O�G�]���c8z���Od�U�O�#v�g٪�}Ͱt�a�I�G|�,�d�F���Ǽ�k���8�4��!�D�X��z��:�Ms�!�t/���Jʏ��'��a���Q�����STޒ��ߩ�5'���U<�֚�����d��#[e#]l�����C��0�_�׭@C�x�<�Z�Z~c\̖���ZK.n��r:jl��]���*�
b--j[���8l߽���Sn����}ۛ�8�w�b�w�$��e 7��[ ���Q�B�m<vg��<w?��F�F7-�~>b���#�WX���k��Od��B�n�z3�x�æ�rN�� �A�6��I��o؇g��HJ���#k��vvtx�9|�o��n�!���g��2`����Q
l(W W��{ʹ`:�f~%H(��J����{*�r\c�(�K݂(��eJ\0v���T�� �3clE���4��%����Y�X���^��ʐ�4�&7A��Cē%8�f}vY}�\�挱43�I}��W�����M�K��ܘ
�i4�S"SY�����h��a�r�Z�՞����뾅v�1/:Px����~&�4#W=�V�=��#4�ZL,�+M��B:	��X�q<��}N����o���cI�	�+C(p�$I�ˤ�Zp�ͥ����"^�6��b�̓��_q��wN�4a9F���χ@�+�� ��V0{��G���~��й��1���D	(�7����R����@�Ҽ�N�T����4m�l�ո19_8llmq����F��f����)��sd�GJȉ����.&�/��|�$:��k:�G��mT���ⶳ���s�.v�kY�Fm��I�{[��a���z��p��)���y��tcȸ�\�Y���@rVM��P\�9FU�;����ׯS������/�۰�����������ր-�������J&D0��S�,?2t6���l�e��C�Ui��xu�!��j;�o�9Caf\;���q�6��n��J�Y1�2��V��o��2��\�Ϯ�g;��܅p3NpY��h/���6��M}~��3$�,O�� ���p��!)l+L����B?]W8mGE�W3����"��q�6���x���3���I��K�m���JD��M*M"r�P��eɲC�W�$�����*Q���9հ��'�g��D\V�T�S�������eG5Aug����K�Q�U=MP��֏6�<nEOeF�KP�n������ݻ���[�� >��D2���7VhlodY`G���@�KI����vHxC�۸�Ӗ���.$�P�����Jg7������XҮ�o}!�kx&�g��zԝXt!�(�
�ƛ��՗ߩI�ހ>����T�G�M@űk�	��L�$�%Jm���i�K�$&�%��Q��q��\� �o���S��B�{�\c,a`ԏ�$'[��e��X?��O8��y徺.e���l< M�kN��r���n���]l�E�TBL8T��� 2�P���'��9�u� �?�,qm�	R�d�{x]���L��}�nF����ٸdh�v�\�yFr�z�;^΀�S�;�:�t��Ov��ǬM��.s+:� x=���8����3�F|e��=;��I����Lf�g[���Jw�T����*���g��X?���ɋ!�Y<�7�%c���kN� �£����f��F�ʛ��$K���������D���C^d5�LJ�0�����,49}�`��R�Ti�g�UŶ�p@��$�m��Q$5���>Q��n��c�i�;�bkDB���XP�<�ޙ�uVZ�/O���iU�����#�!���CH%U�7���Ñ���w�<!Ϋ2CL���E�3�vk��8��`�EK�2S�G�6�(��J�H��'ۉ��?(y���m
��b_��I3��[��h3�Z��[�T�������̩�����#	d�?��=���HҷclFi�`����k8[�`.�O�e���z��DBP�_*Ds��� �r$�t�յ̙_|j.Q>R�+R����_�V�6O��e��Q�����ۑD�o&��ܪ+Y	��4w̰����U;�lO�e���I��#������*��@zgW�Y��c�3A8��t�9$/�u����~z���4ɌE>j�o-��U�Z���d��ϋ���v��M�r/�q3>?2M�	�;=��g��D�[��x��A��oR�-µ�sJF�-N|���1�-��܀�����J�tWu��F�$�M��݆�	%"�"a�`����@�'�5(j�A��О�Ɠ��眫�Ict\-u��%!M D�H8���
�.4 ����K�y_���s���D��}ÄEq/DMBy"���6�����a*B�k�T8��1�o��Ƶh�+��TU�� �5�8�i>��\2��X��'טּ)�Hm�#+ ���X̀���BA�U�� �x`��Xm�}}�Zd�
*`����8C��6�(��K:yꠞ�����"SF�Ӓ�H�3�w'�`lXn���R1&R=�R�(΢B�Y��CIή�ܠ���m���Cȟ=pro�hZ�s��z4�j���ƕ��*��`ū'�����3�b�tr֯g�j�g�����&C������]�A��|��6qXh�mM�wQȓ��a��Ѧ�|�:`tAl�k�~�x�Q	=���\�H.j�0��W�{Q%w�
�7�'��vVп�����-��#�D�4�j��7�$���/<h#�β���-OuL��e�q�p1��@���[VF����N*�H#uJE]��k$���fd#�Hl���Y��T�<g.�^�%�hv@�� r�7�f�h�#a{$�����5�G��1��)S �gs��4�\�K��#��T*Y���ʍZ�����Y�]�9�>f��I�����N;�	�1-迃������S<�~F{�k~)����"���($2�k��VpA\Q�I�,�M�@��~���KiP�M�;
9Oi�#��;�OcS;ɪ�Y$F�P1�q+_��r2_��T�?M�"�,�:�<�FD�X"�b@Mh�.��h�Ķ<G@!yGr�f]�_ReC*��r�*�Ԟ-�C����_.�!���Q�����9j�niK'���{��5J�����KO�""ӟ�;���%fg$��� j4^Q� s��E]��TL��?�����)U��BJ��ӿ|LF�������]���R0���7�����ڟ�ICr�t��΋[՞�r������e��!o%"� ͗\۱�):��J����< �
R��u�?2�U$���5'z�2��jl�$��C����)��V�Q��m©��w��!xv[���)�4j��NW!(����_����g�P��oS#����4������lI0�HA=��#'W��4k�{i�o�o�2���")�
��c�����y}�+��ڪ
-rf��%w��'5��}�nJr���Q�qo���I��D4U$�p��2�l�LgQ�E�g}��/pQ����� q��b	��<B"�'���M���k_b�A����8����h���ۖ�*c��;���D���q��$�Lo_�8�)d��'u��!�~ɰ�۵�Q�u����[7�(��GqX�ԒCT�0X5׹�*�S�'���ê��*A{Fʐ��\�����1�1�q"���I��e�!���d]:�E:Hb�����ϊ8��r��C��^���W����g����߰�W*;�*����	������HR�O��G�����U���_Z6�4z��M[�3�?
�����W_�{$�t(���@�޾�,0����br����I�A(u6�ڼ�w��k
�������û����!i>�X����-t�Y[�%���f��<��j�,�{���oJC�)%�`��qY�ӗ��ӤU���qn��� ��)�6 �B�.�����z7�c}�˸����4�RP�晖��Q�"8�]�Q󹽋�8�FB:Jqi�<�tc�h�T�����Z���Eye���H�������M�|�o�5cd�H�?���[�ܶa�	��P��A'F�_	/���n:�X5�ߖn�2�J\	�xK0��
+ȂaA:7�S˫2�����yT4V�0i��#v�QG&�|#�f��??�+z�������H��)���:��t.�� ��<y�j�^w��0�^�
Q�N��j�DIRՄ�0ZxNdW��M2�ȶ�&"GԪ�I�-��o���M��k��AtG��ڽ���"���J�Z�|dU�>m�`�=(�a�P.���G��,n��"�݋J���pT2��5\��.J�'A��͙WE�`'��t�؎���1m�/�OT!�.0��_(�$�Y�`%�&����K�	ɽ/�
��d�
C���im��#�x�(֛D���X�������_�s\��+z���z�)�~T/I	H�;�G��}s�`O���@�r��y�TN;�w�P8�.zT���D�i�ұ�F�;����?Q.f<2�� BvQUn��h���1�j�!��;�`�L��J��.}�Na/�\s�9bl�gC�~�f,1^�����&aW Q���!�·�A��@A6vy@����h23z2�xM�ud�͙��n��^��Ņu{��#��ڴr��
�>��i&��#� cC1}���>�a��v�KQh��wy,��֩9˜J�YQ��P!?(n$�2]�<ƽ��L�Xj����]��#e�Ƌh��u�{S�dF�.��O��e��{|7��eg�]Lwr\���Lc O{�J�J�� ��̙J��*"Ky7�C_�曔6�ar����M1?ї�˻}�`��!����%=��o���?�]bΠ��qI�`�%�����V/�K�/N�r)!���9i����K��um��q���t/ɍ�Je�P�g����;4T%>�ȍ	�c�� Z����G�ͥ����z/%¾��;�ש�O#n��������|��\4�7Q��j���L��#��
�q+-Tb9��2��U��W������xaE�K{o��3��h�zU�'����j�,+M�l���T��I���f|���&�K��_�<�tX�F�@ڧH�@�1v?����1"���3,�tA�2G�1U{��l<�3t�}[l� $&5�ߟ��`wY*�b�����?("5��tE�:�A0�Q��_aH)��Ʈ��d�F �KZ;"\.�������W��Bʳ�>��G���ʯ�Q�0(T��ed'�֮�L5�B�f��7�wEG���ܥ�+L6(q��D����.�G٢�`ԇ��G�ODz@�5�����
aAodX[�T�us��^�*Z�:���^Դ2T?g��;����������E��������>�&�C�\u6b�v���і������>��rby��+x�d�C�3�h�ރ���l��ﰲø;B�LY��7��ҽ��?�'�U-j�3< �:��M~��� �L�a\�q�bR|׭���p���>ڴ�G�j~eL�:���S}��`��<�Z�h�PC�
���k��vtL*�����[��n�o( �9�>�L�䠽)�:��F���I��=�̵���3�_P��?��������,j�sV�Xf;댷t�hk\�k���MNKI�C̰�@�N�ʕ�d,����5E��bH�{�'k�߰�La�G�.}���5's�)%0��c���y.6��3T�Jd���K�u4ЇO���X�;���z��4^�����IQ^���OQm����mO8�V`Ӱ��W:�G�c��&=>��퓅C:�?�W
H�'��~7��ڔ�O������{��\P���D��h�s�
_V��M�K��	��?p������-�����d|����y�!�>��	mp��ޗ��(w��58�[�ANA�$���N��>*y�NGeB�*�
�j[��͑����T�n>4E�����L5@'�!�3�x�
����(�_ğ�r�A4�k��[�Z���2O��I�$1�g,�f�=*�^�*���	^��H��}(��P��J��;s��r��Q`���Nj���jІ��w�	�z��׭�lw
%˿�Ѩ�
�N�Ҝ�}��B%�Uy׆�qʀ>Rz���!A�"",�MCbT�U�J��R���ݦ��S��"�%��ҲD�~�U�
䪇���7Yf��SX~d ?z$�s�lsW��[�x��BW�ɾ��D02-*�:���j;>اt�`��xF����_	Bk��[6���p@<$��'��L<��Hn�?��忟���u(�LD�;P�z�6����삀`8�{���3�)V���V����z�#F��L���:P���$TF���U����#�L>p���%�<��#�Ósſ���f_� �FA�,�|he�����0') B�=gR��<���O��K��#��A9j<��!J �c���#Wo��G�ǯ��^]vJM�2�Ћ�)��˕LKg/��F|,B��Z��2'��]
jf*��6�P�!���*���#aҍ�:�C����.��E����ڇ|�ǔr�t��F��3�_1�̩d��(]�Q���r���o�on��#`�f}�M�Qd'/�*:���
�i�|�1(i��3S �*K�]��0��k�����V��E��ͬu1�g+�5�,o��(̐�Д1N��q5I���x��*A:�T,��5Yw�+=��^e~/�Gk{�̕P8���Q�����%�݇s�\
����?�k[�܂���8�����j;�B��W��ퟔ���̂�RXv������7G���p�b��0�#4�ŖG[�n"�>"��h�F��P��4?�M���ʙ��h�ʽ����7pY�
�����P��\|Z8� x*bK?ŗxm��'�r�d���9IN��+�
�O�oZ��ց5��r< %���r�w�7@/��j�f��k<��'G�
|��Oe���38g�Q8\;�)L\/eɩ�8�a#a:��)�0r?e��⚏����X����Ը$.�8J�{&kZl;���ߟyX�1+���rR��Hx�bb5F�ӀNp�^��h+��P�L:����CD�g,ըVH�ye^Yhq
d ��Yl@��]�8�Nz��z4q�g2��߼oW �얛s�&~�&|"�O�ӂtNPw#p�<q��o��ս�
l�{�{���}uD��/A����u0�]ψ��Br�q�-[yʭ��-��U�6.ω���������L��a�^�W_p����W%�۪ap���72_�F�4�/v?)t�y�G�M�|�!������a��F{�����5���&�2�r��` �j#�Gג�L�O�XSU�A��u�_*L��_�k�ESN�H���|�^ޟ3��M����RnZ�s�K��I�y.6l�;���ң� �ٔ�W����1f��c;�נ1�g6@΄ϒ��Y��{(����c|���\���*��z�0��]0�Nl�CE�܈a��-�gW.�,z�$����nۄ�;��;o�M�L��p~8:�jl�EvÆ�6$��QQ ����,�R�OJ�+ˢǫV��ұw	�h��q}�ޱqF�t�mZ�o�23Ϲ^O� �a˲_v��䝒�u���'�k�|��'y	9�� ���Q'�1�r�x����d�	Q�w�E�	��K��>����7���[��A�	�� r�	JX5rɳh�va�h� �h�S��RA�]�D��Γ��}܅t�� �i	��*���N��|>�[�%R������w7X��/RU�/3eFuS�-H6FX!��(�Q��7�M�@�GU
5u�G�0.v����"��zE���:L�o�7<��?��0
��NG��)�}vUVHLA8�!�b�b%=P���Y�NY���n?p\uM�	���ߨD��:�[�	h��-�.�1S:�K�?:3������Jz]u�$�pf[`��4C��1mh�j샨#��}�Hc<Q�*��[fݼ�7�aq~;ۯ�F���!��x��B{��~�9b=�U��!K�T(�#��-�N?3��P-���,��tz�W�w�%X�BѤ���žJ�g�� Q�V"�P�h�yu8�}<�rǶ	���u���5�-�w�ܘP�#D� eu_ DnF�t���M��gz�v�f3c��>gfGg��, i�*
��]��oC=��*�	��r\g$��E���s��<�2e�@����0a�E'�пe�Ȳ@�
��9���(k[�7�dK�e���O�t,��)�ȏ�
~�1A�{��Z� ���u�X�8FۮO�M0[��B���M�{�q� �r+���5���=���}����_�R��q��Y����6�j�N�^q]V?A��)�v���W���A�(�qDl����ٝ u����EI5xn@\ԗ�e�?3�$x�Z��KV�����ֲ	lh80%Z�b������u�����j����H|x���Yqd������",��Պ�[r���?���Z~�s�s&V�����(��<U�m/�������W�fo~� ���}pW]=��
&�;׶3-߻�f�ԁ!*�({�Y�@�j�&&�1�sM
�_$���3��� H~մ�G�bc���q���S��@ޅ�%�8h<�[*� 
d�C#y��<+�q�<\7$K��L��������G���<�b�:\]6�V��>��"�k�wo�)���6�<�K�?We4��zF`��ū<}Z�Y,��h�sU�A����%;[©��z��U�����}��nJ��j�}�;��Ah.�z ؑ���ߔt' ���:���������T4��v]č�6�?�ll����W��t�D;�A%�����׶���46+�N�eg��+�,H�#*�r��Q��"_�O�_�[H���z��'�h`�>&r$��eȿ�M���N��^9�#�b��Q���O�R�)�!P$�Y*Z���uB�o�����'�*0T�3RkxI���L����pELs�%��+ǽ~�(�g
��Ӏ��t��[�&.�
i$:�&�	�WS��l���ZR~'�1Nj-�zC�_W�8�O�O^&�#c��51\f#ov�IJ@��&79��˾#'|�I��y�nX �D����R������rh�'� È~��U�T��9*N���w�ITH�b����ZY'ф$��~��CQ���S7��8��VrY�g~!��i����7�a� z��xj&�wN��ҤH�5�Un�0cZo�\�xmv=E�l�J�F���������5?��/(H,�8�±P��0��(G瞯�.���kLy2ګ���G;I�.]ז��-��������Р�;]����4\�&�}���{��Z�����_O^T]�e���F�=���A�; o�'�G�Q�OaVB���L
ǑR���i�Y�M6t�����ޚT����M���$��}+�R&QJ��0(���E5�pi6'�˸�	�G������*���t���2�p���74mlD��V����%��h܀N|	@�VÐ��@�!���J���p\�_�t)���̃��u� D��+���)�y�H�C et�ye
+�Nw���ɪ��C�]Ɵ�Yv�M�g�Lk!;�?��p��Y;f��Iu��+���d?��p]�1�2�+��/�.�rU)�@S�6'�����3Xmj���[�Tc~]�X'���JX~Kxa�*�&/�)�����2�ޱ'� 5�4p�4U˥*(�<���_T�����/Bɔޚ9�(��i5�>k�8���_�r��n�XH��U[��yC��>��gw���b�|'�ҏ��ړJ��W)3�����[�ye�E�^X�\
P�� � c$�Ꝃ�Ng	����o���_[?3p���'CUZ⫿�$��!du���Ś�lAKxq��R�"�k�¹�f]%��b�{��LC���Ln�[���!s�j��Ř�m���8xvP�p�
��E�u2Z|uA`�.z�.��>GS|��8$�!nW�ڶ�^� �+շ&�a#�Q�`K�x�n���{yڤ�z>��9�z�]��R�.DĖ� �u��$�7?����@�.� ��b���ZN�]�s���j�O������2���,f��0	��6��5>
��F."���q@�R;�g�w�����z�,�h���F��>TBk煿�0�e;�� �b��<�ˑ��C���|]F0���Tt���1��p��65�`��JN�ʪ��Zd~Z�#`�����m�k5et���r�.Xl\;~�KH���^I������a�0/��(�7ydMF���V)o�_�Q�y�5�Տ�~�ea�Ȧ>m�G^UME�@�#p��d�PXo���\؟�ls`�Qzݐ\c�������k��]LU��O������)J�N�K�-��j����X�瀦�?7L0��e�b�����V�!)��t���&��P�[�7�o�[`!$c�JK��z�����v�s���rH��0��&��Z��'O� V�!�8ly�i>�V[��5r8�5�y������s�rFg?���l��z��:Aq���ڑ�TS�m�3�Z�؇� &U�kL7�L��ݍn���N˸D&x>�v\B���E���#kG�Mq#��o�[,q�	�`��䨇�l�?anu'�T�fER"�+��͑�s�Ĩ�q�	��6�`�#����V	<r����!��1�͂c�3�I�vD=�rׯ�o��l��P��_�－��^�]TLv�F8hs����9�{�c���H `{�C������L0�w&]2OL�L�d�K�In��D6mO���,�}i�����#�;ը�b��2�%��񗚬u2�����N��u75�_)�_~������_���i�MM�� `XV��Ru�@B%���[�2��l/���s�f�q�~��k�7mK(����Ň�JFx�7K��/��(߶>7�%����{�g�I	QB�N���xX�B���B��Q� V���[�_����)U���@��v���x��R$�Ȑ��7�8�맂u$�FK~����+#V�,��DOVg1?�@�t�����W�&"A�w�/�ζ�_Ť(u���Qɨ��%��B�ehg� ��	�`����kS5N�Z�?�t��� q}�,�NYYz��@;�	+�!ү�ɸlI(�ZZ7XL�è��n����f�v��W#s{��6̟���J�7�&�7"��q�׶?RUZ��Z?Ԏrჷ��&>{���)O'FżUe~��N�!�%��@����U�v�ö6'��*�R$��l�?E��k��6R������K�D��J�p��i��<+��4M��:JM�O�P��U]ykT����p;�W�e0T8�"�Ml�ݾ���x����4B�骹�p����\���N�*�Yhp7�^���͑��o� l���1��~4�PPH���K��TB}I�O���	$� 9�34S ��a0x�,�[L�qh=ʑ�C{�~���%o�vt����M���WJp�v,�?�^�2��M/�P.�.�>�X�~l�]�����@A���ɳ�Uw�dvu����ԏ*e�Hq���R��p��Mt�Ol�$�&mg8��'�/��e@������h|�O�����ON�I�'I�4%����~��!E�0��W��L�.�M^k��d���]���P��X�XJ_�o�ą��?��X$����w���_u|[L�;�Ɣ��TE`�����%t��,� �t��M�$�\��/�ҫ�d=�n� �pL>�1��ڂ�Y��߈�&��H�[�G��d��ȁ��V\>F�������A�wHb�B`>��׋xQ���őO�k�.R	[���/�f"@y�@�����N��������f�3�rNdj��}�Éf�����Z^J�1�>bW2x���aa7�����&��N�ш�s�����FD(}��O.������ћ�O�7�h��\ղ� :�_�i�J�
=$sNG�$������6"lp�Z(���E_�k��K�l���������[TzT��v��p��������KQ���m�,���[�̬F�+�l���({��V�G�^�>�_/����[}e��7�1�tM�����<Ì?���9����gj���C�n#�C��+�EjZ��,�C���j���?V��xb�C��=��Q�����:��od=8�M
�����}�����a���ȏ�M��:�i��^���d�t�@�a+��{g��}�$k�|7e���>���P��'�G_x��=�>���w�禊�M�$��Js%Ad��u���;��.CR��o��:pٷ��^'O�V�ė�<Nx(Oh1����  N\F'/@-��N�}pn	����w�T`ډ
�Ț�� �F�(�W�+%^�  �e�3W���v�ܹ�g�,��z����Ƶkf�D)]wj�$�H�a�QJ�6+,���n3�i.�	�c���AhEC��8@r�<�u�Y���!{04ک;��'8�)NvMֳ�:��t6CP�,�P m���������5�$�h<9�qm�Ȩ;�^IJI~|�ďW
�6mm��¸�8I* v�|&E���-A*,	͎p_�%br��ʍUv�h֊WUc����Y��0���	�=���x�o#��8��c!.��31RQ�+��d�_�Yb�U��-p�t����Z�{�P���3�@/���6|"�q<�aI��y�����d��$�7:�P�t݊~�ǟ8�ѣhh"
M��s,��������5RP�j��L���s0��+���1�7�X�g<�G����jg��h�;�S�5m<U	"�ם�×�!تs��i�X���c�P�#��W<�"� ��|���8c�Uv�&����=���`�<#;@����+�	]z����(�MoX���ϩ.rw�?읈�����䳎��,W�8���+���˘ �f����#|#�R~ �)�/|���/������ʖ�l���9����{�le�D�H�´�iH���.Đ�����������1q�x�N�ᴞ1�w�>@O1��R�7�`��͡�0�;d:b�!+���@�0�S�I�~�s%r�Xh'�g��6$��o����	-�Q1l8a�h��\�<|�n�S�Q)��k9���Gu�`|p�Y��iܔ����1Zb4�"�8��R�}���s7H���;��mx�1|)>�n|�L�e���j[1AZo,��z����R�>Pf6�����*���ybr��Ƨ�������+��<����	�XP�7�������o89����D���	� ��e'�.������"3C�"�3-��<���ubGi��,�6�
�B�\BC���Sᡳat���T 1(%oEM� �3�n�	v�D��v�q��;�u��#_w�i�k-ÇL��CM�4��/nx	A���(���hJ�[A	ck�ְbM��lPw�7xI"F�Ox�V��;��2���D|����.&�R��\4���iP��Ѕ?Qa)� ���q��It�e���L�I&k���#uT�f8X�{T�e9Z�D�ŹN�Oqg�O�+��nQi7��8DR�4�Z�j��`=�j<L��Y��rw-����:���T~���07������g�
��oKp�P9���&H�96�@_AO�(�#�S��U�h1�lZ	m�H�]l�#)~�� yG^d"��R���%d�	|�4M�^��_�&&��b���w(��Z�<l{��������>�I<3AB,���8S��l�s2�[p&A�4�TCC0���;,�"�Ե>�:�̊[�JMylۦb�[f4{Y��P />Ȭ-ی�	��;M�bf��R5�b�:��ߡz��	��>��D#y�+���ɤ�6�d�qNS��_s�C&�	�y��K��=V�&��r_),#��ڧkDХr���Qe+�z�yT��F�b����
�S��S	���A8{z�(����]�檒�0sV�=NP�,y�f3%%�%�M�~�"r�3������ŻBi�;e���1z�j�}P��br����QC-{?Fr�*xY���Kx}پ� ��6P����=�!6<! �_�Y!僩����a�����E�;�`������!.�"� ��S~�ˁٵ��D�|���r{Rr��^��D�� (����IA�6��C��ћ�o�w٥���]�@`)�x�7W	\ॶ1�	��Ψ�^C''� ���V|��zì�v����&�YNN�ՙ)���e��W�E����kS�m=|(�n�$��~���4�Hv�8����ΪK�9ޮ���iXZ6�٬��~W��@<�M�+޶��u��-6sh��GNK2.,i��$
L��=�b?�J���Hǐ��US߬�˟����zJ]?ϳFʒ�M���}/āc.�n�8��a>PD���8�fcwF�21i	���T.����r���������Ө�7�-z�.���N�����ܖ;؞�k4s���b=2��f]EU^�8���8��h�֯K�9�i�C��ex����q�L�K��NE�m9���b�C"�1A�U��B�,4�#p�F��.�m��y� �,e�G�|
h%�ASH�"��PT}��1K�Yyn���?��q{8�8�0��,�!t�we
�[�!rze��}�`Ŏ���T��͗�Vv��ZTD銣U�s�����6�.�-��͜0{��0����2V��PW����$���_����Q��&;?8�X�R	X����t9�`�5��&�5��ӒE�Ha�Ě`��Ս{��^�+�F-�v�y����+�E�7<:Z���p6c����FAw�+a����
�FS����2)�򔍝�I��\�}y��ᗨ7���O�S��qp//�+-(tE#B�w}c	�5�:�\˯rm���x��ȕ�{�EZ��F��j��fØxB�>��n� �sS�����	0}�fȆ�]}|���ѵ̲���y�'� ��ԳJ��j9\���b��Puϧ��}��8�H@[H0|�iS�i�Ǜ���>
�d��Ӟ�/Sv2vͳp���-�}jW�f�uȵ=j�9�����#>!Gge�F$4�}5��k�Hukr��9r��9�	���S	�W�;6d$�7~ y.��S����cWx7=T5�fٟ�#�<��N�1
�W�v���G���C[n*ܞ�ޏG^�pS�u��+c��B��.;Ph�.z�د��@�Z��W�޿������3��U��[�)�ۦg���s�$�c�xJ��2K�mto�:���n���ۄ�	W~��(��'g���$!5>D��� d��q�O�?�Ȣ�,;�e4���� cL�����E�8I �(}ޥi�b@?ڮ;Ҋ�+ب �,�o\D5Xl��5� �+扱@�f\�\�=�vi�������=p�@�8o[����j�,!#��8�-���kDcıO�d�c
 r�
���kS��0'us{va�X���f3t`�Dk8�#0�4�8N�J��\me���Ҭ���Q��2����m~�#5�uZ�Q��P��3�E�$�o�3no��L�)m�!O� ���Yb���O���Ķa~�нd����}̔F� �y��3*�@�i0���
/J�6����-���3ðaW��ċ����������EP~R��s4�v��RAJgx�p<R��� w ��P!q4�z�^�Ť��ݡRW?Z��;�$�z/2�O�G�"E8��u�&�.�<~���@��:�@�Z���ܐ��P;D
�=�j1ھU1�!HKJ��Y&׼�F�u�l��^�A�%4=����UO�=D����7�ׄq˔m,��sS��C�/�r��#,���]�^tn�W4i�S���o(�P�K��^�my�%�+�L�|	vՔj����L���v���@1>Զu���#��0.�5�C4,�P�u��d>�i�iz	�v�k50hn��{�"E��y$�?��#*
A-z*��5,(��KaV��d��fA�j�g���n� �����r���ð�����-�ōVH-�t�M��˯9����|q���.��5z'�x�����5����2)����B�K}��s �Ci�2C!�z���$p7�V=��v�)( B�&�K��b�Cl�@8b9������}�!?X��V�LU�4����И�Y)�f�����#A�Zָ/!6&<�SNFC���һ��):�>~6���˄��s����&����J�G��;�*0O<%t�^���T ����d, �7���K�ݍW=���f��0�Ɇ
�('�hS�!쁊�
��@�!��=i=N�XM%�����ϔ~�#���
=����:/%��k3��ޟi�fr�K��_��jS@�'�2�L1=1b�1iu�X����siOφ�&�-��1k&9��Z ������9��Pt6v�\y~����WM҅�rD���i*�4|��o���[g��3ڦ��=�A�OQ�c��&�,������P��9�G8D�km��¢
fǺ�r/ݩ�u3�_�?L?�� � N"۰��fC)���0�t�e'�Ѩ1+y�NE*u�k���( �[U�V�<�_9��BƵ��n.�������U�*Nr��3��ex�p�E�觻���l4܃ݸ0�Rfť�gF�͙5�t�A��p�J��/��RDk(���w�3�_���I�l�hZu��)�'�o}�V/g���ϰ)x8����ݺ{�c���@w״��Ũ��)�>zq� �"�Hz��v�,Y���� a�UX�-��H�����|Z��{�֚��lvH�65M�W����~@JDZh������K�/�{�
G-Xj���h'��c�J��l����3�HBN�7@��|y�o���a?2B���pU|ȣѿ���!�wR�yI���$N��L����P�E��&�9����/��N��Qh��zxS�iۘ��i�� ��ғ���	�L�fqta4����8r�y�:Eކ���-_�lg��ذg#��q��^~iJ�w�o��҆�v�HL�\�K|,�&aZ�!��=��I�M�*怺�7f��*T��XX����j3�s�i	�7�-�Ь�b�?FY�kWA�u ���y�)�)�C6��{V��nv+��ϫLg�؊��)a�b!.��7��z�B#�ʹ���H�
�_��a.�1��
O��l��g�)�L)����[�H� �l�w���J���%�v=�?�����RX&I������;n��,z=�7�!�L�A��&����j���c����!~^�\��~G�f�2�ц>� DL,�At�=�zHy�^�u!��U�rm�or*Te=]�������O��?�݆�k�1b&����+�l����,�����2�G;F�f�'������B=ini4�뷭���^�2pK��3����b�]ϟl��udd�v�Q��7c "��R8�;jDv�����v{�- �֑�.=�A��頇�'�:(~
�f���3k��~��d��'�/�࠯��������e?��0��zpg$��9ۈ8�i4g��$a�|A��\61���h����$�p�T��;)YH`Q"�	mb���0^'x��a�N����p�1�|%�_���/�d$��q�/����(0�!k���{����+<��J�V��94@uBB+�*�y놫�W�FK�~<t^�n[�fW����1<}c�f}H�]tw.�7БU�Ӹ�,�yX_���ޑ��IhP=���
�@���	�����X�"�=0v&&�6©Oo�6�d�a�q���7.����`��˒P����d��9m��`��i���\ȕ2�V�6q�>T�'��$��h�w@��P�O|Jgf��V�Vh�^�������!%�v�����@J������q� �+fPn(����8��I�«��+��v<}@[:O�wH0�c���|7(�ۃJ�_�B��H �]�D�=�S%}E�+����O���b������XL@�8?U3u�Z?%���h�|��vB~�����I�%�bE񖶆�9�mY��\gZ���HQ�N�7���A'�4O�I�o{5$-��taq��!�t���ם���S���|ny�U�ɗ^x��Ϳ�j�'���D�/��*/o�&����R�K��)~7!3\���Nҡ��w �*ڦ!���S0�����Ѭ�'W�-���п]�ˣ"���#��WO_k�$b]��Kݜ^���^�/��Dq �_:��M�U�����E���Ei�)�DR��ޞ1�)W`�<Kt4G;=F�sZƝ�kH���NW�8t��`U���}!�ݵ�.l�N�#�݆��q�Ȗ-΅�j��[ب��4� �����R+�ĕ<��bL��-s���4Ňϰ,�]ƱG�>��K��Κ5ю�����^�^��;T2?�z#�p�;�� u3 2�H+ޕ��?Z�ƕo�;n�����U��.�ψ����|�Q�\�w�qK��'-[=�m�bü/����w
Hd[c�A� jx5���2�����;U��\F��vwk�aLB�4�t��\�b4rWf�8(1D��r�Tz��\��l�=��䍎f1i�|�W�2�Os�~O�wZ�n9�ջ1VmY��l)�EҝT��8�c�R�(H��e���	NI�6�z�tu a����b'�WL]�Ȳ�4���AO�~�K�F1���u�6�|we��RZ���y�Vw��#�������V��١W!lG	��:���1sվ7�h�nrو��)��䈇v����-H���OBU�Hs����$�����^F����OU��&g�6X��#�S>�Ȑ~G,v*Ƌ^����e"��yT�-@��㤊��׻�ܜ���J�B�ӈb�d(�r�M�\!_2p������w-&q�T��h�8;U� �`Oeh�������v鯜�� �G�o�2|r���9��PW+s0h��@N�d��U�d*bQ"�J��Sp�샮���-{��#U��/@N�(lD��0!:P��Xf._�6eԦDo�C1&v,ańs!�C�ٷN����v��Z�M��HKb��I���F)&0d����bT��]�7���E�o��)���n
�zа�_�DȖ7�@�<�x���Z)���\�9�HD[ÒC&�(0�Ph��u%�r2�Lnw�-oE,�c�E�aI%$k�Pց	F�e{�R)�Jq�=ZLP�^Cc۔��i�G� Ô��bf��+!�:|^ɣ�@�濨G�J �ڹ��5R��B̤�&q��~�>��؞}-��l���l/!(2�V�����/;���@�#����q��]�L�i=�,O}�n� l(V@��Q�N�� ��k�e0�"]4�!C���6�/�_��03�tLUx[g� �R���� *
#��Q��|�6˦@ϕ]đ'���k�)�u�g�`��Zl�p�[�DQ0`�>9Ss��eQ�	y�$6T�J�&��֒]7ƨE�a#v���f�p�yw�ƨړ��nu��p��^a��
]O�b�*1H��J��{�l�ۿd��v�
�
i�����G:p���p�-��\6B��,�����)X4�1<�y���AL�#��k�)��p �f,�V��C�`]p�U�7�aM����r���O��P���Gkl[�B^EP(=��Hڔ��f�6��@�"@8��k|�4�z���O�����Z���BG�sK�b�m���8i�@���g���"bz-x���`*e�8-+��b��R�FF��b�U��}�����8Ia�ɨ��Ki�. z�RZY�ARw���ȜL�^�R;�D�^�W3�m�-��P�['�����մp[)O�E�ڊ�����X�^X����`�
��3{��FR�0 ��qẽ�_�q��В�?�K]�ҙ$h: ��༮�dv���ߣ�vq#��2c}���.�^��^\�6�J�O�̕)5��Й�	����l�Sq���-K:Ě,è���RrH8{��Tu9;��,`Sg��h��Pe��"rf�
�"g _��y�'����/���T5�e�楔�wc$}mlV[��hKAp�����^UZb��0����[)��몍���G� �`���A�Y�����ā�$*�ĹCo��8�(������ȥ=꼿Z8s��煒$˖�f;M�'wt<�0p�.�%�-�S�������B�=����ɢ��!p�:K)>G��!(�D-^�.�/��h6d��B�[�k�X!���p9�5*.r���7��,��N����?:l��g�a�\��m�&1~�� �c���Y�6/��|�`���.^h�(J|%�о�3�y����Ⱥ�%J��xϦ�I�k�41'�����j�Lr
�!��0�DH�Ղ�p1�Ĵ�a�H_
�]���O�yL���4����<�J�oC���q��p�D
���i�����B�'�%����^smx��U�\�(C-�P�%B7E]���=��Y�d5��Z��%�?.�(n�+�.��<��
v��$jI���EwTcA�^\*���[X6a2}	`IG�e���0�sG� U������k��LV�2R�\p���wiϱ풪]m�(�j�f�J�����Y�`��(&�hZ���B+f*4jE�J^��E�v[HfUo�e&�w��O��dc�����T��/�Zh\W�ܽ�d_��ZHB���";_:]��_Ze����|���y�����^.G�u��@�����W�q����߰����z/
㜞̦S�U���\s��9�����@�wu�u�R)P�����4����|�}r.1�����wF5xc��x,�i����~��A�t�����Amٴ����Iʅn�J:���&��8���g}鷭_����-��s괌=1���aE�`�_gz_M�I����L&�E�*u���0w��N����
�
]M� �w,�%�7�zoT�
�i*��D�C��c�D�=忺��-Ksu�����Te4�,2(c��y'�^Q�pX��z��j g!�^$#z��2k"֩Ӂ!�Ku��!��G��z]�6�a"�d[*�thiɡX�6���7[{���N��KX��]��5�8ʎd�����[�޵��X�gn�B� 2$qp�G�ߖ���0ޢ:��
7"R����"�[��i�`3��N /�������P� �s�m�Щ��;Yq�qX
��{BP��6E`��'Z?���Z��Px��!��ւj�,!�#x��=Ҝ:����1	���yA�a:���`8k�+��;s��LڷҴ���E�?���m��2�>��S�(�i��#��q'���tMk�l�K?,դfY�8�zpAτ�Hmmm����ª�@�R{q������3�Ӭ�:o"�2}��G~��(PO2$P����v�?�N�f�E��U��,-:��utܗ1Of�z&!�#~/U[�:s�h�B�}2xf(��cvJ�y�u�L�g�C�[����h��M���J���Rpy�c�ۑ����J*������|#���\�%���>�5���jSm�[��+�@)�عr0�k}�VpZ�)���{=���]|�@�^/C.���^�y��W��>����c5
O��^=��]Qw����ܯ���< �.�%��o�6���w�)Q���KE�:0�i3u�޾���˸�&���Ӈ�J���v��74g�s��D�Q�f��Z+1,��&�j��,�ݻH�o��h�K�l?�. 1ީ�NN6�!x)��0�YZ��@r�R��hϩ�h��GX�r�-��17�����8i���oQ�۬���X;����VN�g�K:y�nD�_�K{����ۀ�8�{�P�\�!fv���3��G@yU��(�A<�P��S��
����O�: )�(�B�48�DN��ėq��9Z5�^��;�Y��H�AR�f��7I��1��D9�I"�$�p��c��Oh(Њ�!��6b6#�ؼ-���&��)1� ���j��]��PI-|����%aDp��*v��,?pP���{���ޅ�L4՞���K/�Y4�'D�|,*B5��̸B���Q�gI��0DF��5_0����9�e�WD�PVv:\��,+�|�� ������)ġb���lB3��ycHi���������-n9q���2�X/a�DR�(��b��a�2`X�[)*ִ'@��Hz:�_�*���4�����=�`D�����F��QUo�L���zTta#9=|�1(&�߬K��޵���?s`��d,4F�=W��!͒�],RO�A��h��)Bst-��Ϲ�v��y���X���/�D>��p�_T��No=�*;|�p�zL�����1f�^I�z̿Kq[�DG�R<$u0ި.h\Υs3����I���Ū�yH�F��Ծ��FS�K>嚀(e��H�.�/b-p��7Tzc��b���,�R\n�8�N_��1�+Z��L�k�ݚ�H,�>����B&d��l}��p��XBZX��{�[�)\�4-�I�/bт�����8�N��wS���_���c�A���j!��Lҧ]n�fоѱ��H�/��&��_CYơ����A��Ȝ��ʈ�ԶH]��o��ԍ|X�� KxG$�\�m�����A���|*!�Ṉ�ᙋ(�mwl�X:��5��ESr[#ɶ�Me���~WQQ|�Й�����)$�ʷB�ګ裈l~�O[uk�=�� g��lSd�so��O*Ry%��ͬ�t���RFY�թ��7P�,�f8��pb��J�a��'����n���c�OCXw�Z��-P A��ȑ����J���u[��Z���HB]�Ϋ��*�+^W�^Wi��n�����/��K��-���]��[O�:'�н�\��|G�t���y��2Xckc�Ӈ{齶����g0��=O�b��G��@�����o
��`�?�sCb�h�5E^ؔ���T�*�Y�OJ� ���ˑn�ҥwJ԰�Vi`f�B�)Ή���*ai��6v���V��E!=���ܲ���
3A��>������a��d:�D|�?	¢�B�nF&��ƅ8M#N�+�{IqA�5����a �{9Wɀ�y�x��|�r�����W��-�f�1Zm�Qǋ%tO�e���㧴41�a�B"�Is`�P���9�MzYw��CQ�&_�n j�#����1LՒ(V��Tb�\�(3g
�'�陾F
 .�6�md�}��� ���z�u���3��1Ԣ�q�_����kV�j�9���K>�'���@�!�4�P܉�Q0T�#��Ò�Y�7_��LhrM{��h�i��do����r�M�F�M���@h��|�M'�K!�b�E�ݼ�k1h�x��&�^� UB�h_�����W�PIZN3��>��]��B���=,��[����$���3I����"~/cD���&��WG�:��X���ӛۛ��e��<�K���T��5��d����k(Q5�d�NS�_5�DF�d�-d^����d8G�l�jP��,�W��bI��Ts�M����/V!�W��9W���Z��ƍ���z�x�����XG%��!�6\�U͋\��QW(������'Ʒ��d(�}�}Xl�����#��a���y����}J@Ù���4����.�q�<�~n�����+S�RK�'��;��NzD�nUW�S7�:H`"*�1~n�P����o�L/Q��6�\����s�͵+ϳvy��o&�x�v�������ǥ��q�@��S2OI�ֶ h>Cf���*A�P���f��X��g�1�="�Ӳ�T�c�Wh�!δ��Ӥ�62��F�[�V���o+�Ҙ�Pt���P�Qd&�|�ZB�����
��� ���熊)!w�p��ꕉ�������/�%�3p2��]�F\)��S�^�k�G�Cl�%��|K�!�f�4�E2v4�'k��7,����<�Eۜk������.��Lס�"{Pz�N6S��\�Qw��	n�{l(�Qu�_W�����LZr�"`�w/x�f�.�}.�0W_���y���ۺAM�{e�H�� �]B�	�~������$w�`��?���P�'�t9$��+_��h���*H=�m���f,���>����0�N��*�o��n[8���V�E7n�;��Kb����4�FZ]v���Z�(��D�xf�Y�;,E�-G�<�O�\,^
nb+�'9�gm�0�.aa9�/�w�����Y%�����$�ҾN&j�K�.�#2�^;=��{b�|�2�Q�ZT�	�a���E�zy��^
���9��٤�P;��s����HQ�# 9K�y��(S]n�`l�T1\�ɾV�6���F5�k9�<&�0�E)r�)S��?�b�w�$Ǜ����G��Gك@�j�k�=Ҕ#��Y�{.��5�Z�y_e�¼Bm"M>�'���8L-(�v�z��}ѯ�ȕ�Mi�#6Ե�kbVv�k��Z�%��.L��0{�XZ�k�%�(���������s.�h4UWt͖��[������|�|��$Ұ��(��o��a��Ne�3C*~��v$(HviZ�gR'�C�7y�*/�N���Q�ZIl)�D?]�|�Y)��)�G�D�B�����e�۷Rmrs]�v���� ��L>�1�
SD��c3��Hp.մWDw���!ָnm�~N�\�d�kC�w��흂DMg+��9R ��{��L�IŚOРd���������u�	d
U��n��?#o���:�!D�Խ��¯����w�a	���E�*ţ�`�V�B:,U�T�Q�An�#D�$�6�. jlQ�t�D0L��d�(5~��/I֊E�@�i�/�u��u����j�������$*����JXDKd#�	sc!4�}A-�$r��ۼY`u��T�'2>����K&�[�H�+�U��0{�Ip�7^�:�Lcr�}X��~!�Qǀ�&�)?�S|%�x_s��+�:?�$;�р�͕ ��cx�yHqN��$+q1�^�#O�U��)�j�s��-s�d�z><�?�P�-���=�6����}#&Aa:c�n�C�J��#�L��ͭ�����2��qV_��{�h�����u]Hv��*�W�_��E����Tl0b���T�ٌ~tV� �`�(P�;�J����936J�C�֦��L�_�T_�#�/��N�Z������S��f�zY*�H�ߜ6؁��_��˘w�^��jk@mzO�P�@"�R�~��w��TP���\hM�&�A�p���8m9(��	OՊ���CMC����7(4bi�
�{�َ��1�^T�Kʞ/���&K"t���g#G���z�KF������%7�f���e���N���^+]Ey�8��+���$��DP�#�@����ǵ�&4:`pʮ������xiQ�{e�*¯[����Gi�_d�[}����q��X�+^����?^M}as���$���{����X� (�,������v�o2蝌T©|k��p���<��O�/��*����̢��������5���;�]�99kⰩFc2D����g�^�Z�Jt}P�}��ݼ�d-i����+� �3I��^����l��;
�2�R�\�pIh����H?��SmH>E}Oʽ���%%fe�2��0꺩�0\�ԉ�4iQ@ʺ|Jx��C����Թ��j�e1��ȣn�=��m���6�s4�a�,<M\�\n+7B�o�q˳��>pz�-bE!;���kd>��))kN���gz�̔<!�ˈY�5�����oJJ�,^���$lh�Gn`M�e�,���l�h��[
�:{P/ʋU�q�ٕ ����'[��6X�mr�'BW<kn�t�@��'���q����7C��3I^�����u-���J�ImjE�[�X�ڣ���7XR��#��il�	vZ������U�����U��_g��כ�\)B�[ѲI|"��9o�+�D����b��V�k���z�{�6 u�@��}0OM�s{\�:�.�{�-��P	��Po� �t��'��|�|t����˭��N��U�o�9��P^<�x)��i���H�P��?IU��	�f�Y]��:��/h�^�!2T%�@m�m���2�\�(��Ѻ�O���Fk���LA��m ($a����Z�,�J�t
��d���k�߰����]jGǟ�8�wJ��Dtʓ���Q#{zno�m���_���T��A�z�����!CЉ���8
kO�\'ܫ1D�~�L]�C�`Y:޽r�ۉ�ck�k�Y���I�g��a�~/<�� ���m��Q��x��
��#�Ł�E.mf���#����o�0���kKp�"3�) &���(��e��CD�ǽBY�#Ի&�C*����f-�_a^v�N��t�(�1&M���&�BI��KmRXX�o���k��N���'P��rK!p�\�lT��;E4�9�N�P|�jZ�0�o?˪��c�W��{��&��N�����*���"I��O!���:��2�{t��r�ԗ��1=}W��Fֺ��R��l�I�8��I�v�o򎐘�b�����Uq˽�A�6���Ì�&n�?����?����]�����JJg�0�?�ߪ<ש�9�#:a1PL�vd
�҅����62�?a<A��M)��G!OuEqoP8�`�-��y��wOZ���ڢ������{'�p��G�d_\��@�06 0�Ϣ�Sd���s��D�h�,K�� B�l�^�F�yJ��ϖ�����2���B���Fr���i�6v��,��
�M����*Q'Wפ��w�gX�B��,���?@k$��$Sʕi��r���aNF���	�B������.yq��M}���QthܺT!؃H0=x�R*���r���5�`l�2��Uj<�a4�]/�O/儚j��[*\���̵���MF���`WK�z1L�lE�� ,��e�QD��<X�f"oZ���x��F�4��E�+0+�IB+CMYU�Ga�\�>L��v'��O����I����E�F$zA\�İ�6X�Fs�늈ͩ���AN
����n�\�2k��#�U�wd j�F+7���|����t�\��(r���d�Kz�U�^u�=�|S�S����q��Ytbk��L��\��-3𙶫�҆!x؀ s�}�T�?���pF��T���0w��B�N�?0�k3{�)ɫ�XF<�ز�R$9�E}	N��=E��{���!{��fP?��g�$�E�s�#�9����O��
�3~�Օu ]-����v� ��֧�X�ZPㅊ�3��jr��H��|VO������tƷ\0��*��O�.o5PAM�u�@��K���|#�!�� ��,H����?� �/��^Bݿ��~���NH8�8NgI��ʀy� ��3�7s).>r���IZ�y'z�10*5٩��Dv�q�&+?������ɸ r}o6ˆ����MA��8�~hn�VI�r !P��`hQ���ui.EB>�
K[��R}3:��e��S����a��7"���!���KCT���&*�N��A����@�M���jj�q8�L$4��I�Tq���ڧ6�_B1/U�9�����ǆ� �5G�뎟�d����eU�Y����)j���7�k�c�-Ro��
k@�Y���)>t��/�9'�L��^0N��]��.F�Χ��^r�,L6�ˮ~#�׆qr)��VQ�<yL��.���n/�Hg�c�H��-|1��b�R�� 3�2���K{K+B2�*�<�F��&��0�C�Eh9�\����TO������Al�nO�T	7o�n?i-����:#�0k"&K��E��g���g6��~`����Z�LӶ��|���E��r��/֖�Ka`��Ǫ���6>O�i�~�ר�$鉺8*v�>[�HC|��YB叜ށ�����������У�b(`7�hϤ/���^h��C��X�c�� D(���0��M\���e֡%v<$���XV^l���"cǹ��D�������b��1�ݮ��Er���$�����NT$�_r�]�,��m~�M?��bͥ��炖��Ըb4������'���xp�>���K���[���Q*�
�S����u��͊۽����(aI��9�Yp��լ����$����,�S���['I��(	���J�<rJQc=�)91�+}�|�@�H�U��T�e�ܐ�������X+�����n^���=>1��x�p>b�w�8��+������|U�ځ�LVκ�N˚�"q�{7��묷�ٳXrek/@&N�n�%G��:�]Ի�g�e��(3�+��(L�E�]�˗��Լ���x��Ơ�şj���7��hC(�)L��۩Y{;	�cՠQ�'YK�^{K:���/����p�!��	������(�ޣ����x�"^�ø���N�=m��o�i��tDx1���4�v��c6������Y���Y�4����E_C��;W�VvID� �����OT:��+�7"1������v��ͱMhކ'��w�]��X��U!�VR�z2�����|�����ò�v�[$f,qo�+�0w|N$bӟ��A>?r�=��A���F��a�%���R#r�W��%�n�v4c��!ց���������@P�)���c���_�px��U8��BF�]	�\K��tC��e��Yfcf�N�gi~z��0\m%�]��wGJ
���[Yؑ�k�丙̈����]�E��޳3��MF�NS����)ѿ���fO��U��I!���%��2�g0R�Xc�}�#o��b伏(�g�v��q��Y��D
(Jd����pt�9 �T4oc
��G���L�x=V�^���#M&k+�^Ƃ�����A����ۮ�Ӱ��H0^�H���o}�Y�0	/����E��)�Rw�.��=Η��MY�e�ᛅVw`�`=x��В��!����k=�����9&bLW�HO5e�ЍFy9��b[*S��}�����C�2<wKf*�ңN��̬����60�T��Y�`�E_��ߥ\��}MB8h��4Wo��|(�H�ΰ��>~Z�υAX��f;�B�a&l<#2XE��z�ĘpJ郞 �TS��rҺ��ks�^����0�G���a;�_J�Q�J@�wֹ�]�.��C9e�&wgjF�a�?��r�����`Xj��M*m<���-���[��8�=8P�����\���Fn�Ҍ�F>��Wu�W�����O�w�)��p	@��G���4�<���5£����r�W){k|�onN�� ��uI�$`�=YS3�Ǐ6�]��p2�3F����h��1h�[ ׈�I��34Ρ�GO$����[{������y�.@���z5ōEƍ�w]@Z�r��E��k7��(��m,�>�}� ���G��Xw�,id�P��@��]��Jlx�W*�<�V�Y�������>I�h����W,��x�p%���l���Hu��c�~�Ef�eh2uV?w0�4_>5�6�|Yf�:M����lc]m�u�g�kM_�2�TTU�P&7����_��M(�K�Y��SȦ9���R�/2'���Xdix��b�?J{�*=�o��cۈ���FyF6I����@z��6p~�kZ�|w�E�<:/�:�g�c�X�����J�Ua�Z$F ^qUd�^��#�k���p�!?�_�wy5�v�X���bh�ƅW�n���Uw��Z�=���vgTk�lt�-�_oM��a���l���{��>�A.k�a�;W���2�E���$0F����@��~F�^�.���:ST���a�(n�	��Ol6��*W^�z�jg+.�PT�ڃ���CXS����9{�/��h�7�	�~�y~,����\t��#��uR�#r�9(���jMy�٘y%_������]	��bU��Y��0�I$��q<~��N�� �7���ɮ=>�s�U�4Z@�Rp�G_QR���D���K�����b�B��tW@)]º�A��p�����Vƾ
�Z�w�lbު��@qVCe��h��9�s8�b��̜Hy��� �>��뚻�;áN���:��$��{��mXra���v���o��|�ZZ?���R	_F/��\*~Ǔho�cOu�)�o��۫:!T�h���'��<־�n��-H����5B
�}�qq�&X����My�����T����v�Q�K��>�tJ�#��K��e� ��4^H��|۶ښP��6��ߍ��Ӥ���T/s�R*��Ol<^��1��G�bc���f�6.&㗮dO��������w�n����t��T��m��޳w}��]�b����Z�>��@�k/�gw�u	�?��8w+�z_B���9���Rj8ΌW�#�p���@���ܨ�r��$~\��#�8����Ha�|9Rɽވ����=oO��R*�\�Yy��<�q&�Ep``��
�oY�p�z��$H�E���H�h*�:dvJw���_�I��L�;MB��|�r^��� ��QLD�a�Zg�X �%��-'�1���4�!����#���:-�ĭ�scQb��	��Inǳ�����A���Hb�I�A��7�5��:�"�D&&�K�m �]��33Kh�MÇ�T+S��ũ��Q�3݉4ؽ�)�Y�J.�#T�r��V����M	_d��+��F�ؠƊ�iK�`�[3c�Q�ۇ�|���h�޻��p(N7����B���)}��P��p�wԨ2�8��]a��b3�k*,��4=�j��qn���
����)�t�3�������(���(�i��y� x��2��P?j����r(��&nqQ�f�T#O�V�3g���F�GS��9b+�^�_]�{PΣ����BM��nU���#����a���Fo� �!��T�ɿ!��.?���\ۊ�:\�vd)T�+\��Gm�(�܌�A:(�=�1��h��(6��>�n�N��&��p+NP���{�k��{�|x`�L� �[m��R!�R �����:�
^%�Y�$4&�fRͶ���Ov
��S`SU{�W�ad������"�Pi��`�:�.�Lc�h��f��+k#�q�p�������t��%��ᡤ����	�J��G�aJWŰv�CY���s��x�QI;�]nѡxn��i�T4�ٖj����V�j�p���O:DE��K���>̘���.�"ǂ%jC�E�e��t��ŗw��l�%�ъBKw���^j�D����d�3D��_t+<i]V���IYQO�ÍB0��^Q�3Y��?�7�a�����ܺ��Z��� n�:��n�-3=�w�TNm��[HRj]�/Xe�yXEŌ��+ӱ�i��6��8�j�ƚN��\
n���uz����?fթ�-ݢ>���!�_�aIDO���0a����_jX%�[�L�[{ዲ|{'Pq�0}�$��|��~� #�|����P���8�����mq���[^v�J�~�?qq��˽��lf?�Wy�h２GF<�)_�=O�k6����ˋs�\���0,8��eu3=��φ��_�C"�p�_��j-]{r��ݗ���|u�x�]xj��d03s4����{N}vX�Y��jҼ����)�q��M���yw��S�O�����e�=g�K0�g��j3�h���WJ�5����e;߾"�3{�dM�l���Q�5C!:�sJh��cP��WY-��T9����{M(,5�����*p�i�s�E*�H�V�7S4�RQ�u5R6�=���L�86�F2�J�o���kC��ސ3mI�7�(x�w�p3,��a�2���t����s^���Q�8#ؿ��܈q��	�S�\69���y�٧N��^�p�^�^����e�B�"O�ޞ=B0��D���?��Ϭ��l��G���7ըu�tϲ�R��g ��/��;a�S�������$�&��}�PB��`�>�4r�׿K�)7���K�|mF�JU�b�p�������1� ���[Oh}���c��â�?���i�h���6S��F�c�gg]�)8a �(I^Y��E���+g�%Ʒ!M�����<��?��I�~ll��t�@��7��3�-"�]���0<�Kx���$�a�j��У�_I≱�w$d�����~��T��#�J�� ϘCm���>�*��0�y�t��&��#��*&���s�n�^���I��X�rl�zC��O�u�-ݵU��(ik뾣���6�n��nQʳ��l�������Ǚ|q'��QK#�
�X���5�76|3Ma:-�͙d�Cnuaa��dj`wG��qm�|��4ػc��mΠY�N�y�4�VaɅ9�w  ���/�~ł�x�@����F/���3	����M��_i��ȗ�c�yR���,��.5��;��+�w�E����FM�/ck�5��R�RxA��w9�0?����:U�5��$-'F֘���t�̛���FmHw�}��H�ʬ����`T�G��N�K�/��׉R4��B������f�7�X2����CMb������;!:y�{��	)�lB�@�S�Y�^��7��
Fuկ
qx#:��,�m��9������՜�mB�6؛�R8&�G����A�F����Ǣ�/V'�p=�S����� {�<f@�&�[����V:7x�T�'2p���zφ1��#߲��5H���p����+Ό�������Ċ)��� d93Y��F)Q��$6��x����)�t�B@�WQ]Q\pI�5�#���>֟{\��Ba>��%Ύuuy�y�5��6�21���[���>�d��R'œ��1gu���<���<�&�v�a�d������L^J�;��_"%:�m3 ,���/���td�el��#���x�7�
H^jR�j�����PK�./��%�g��ҪwRm�A�ż�\Z� m����5K}Fݶ�	t�t3��Y�Vb�,�M��JU���J7S�0�%����^�3I�'���J�v׀O���9N��6��2������D��h�bX�⵸�ƽP�z��q1�_Y/���B�k}�2\�N�	�Oܰ;�Op���o�ULn�>*�ROn�E"��O�?�ܺ�������RD���ݸI+���̴��Vۃ�aG�*ȳmU�vZ��e��	�7=h���͙rc�G\Y(���a�����י� u��K��%���h�q=ȟ���Et���?�P+����Ks�V� ���3��Ն,[�<󣼕�n�L��	!�7�UXf�_�D}�d�D
�,l.U�L�鲲��DM�2�����%��I��$���[�s:����UHi��}���c qp|� ���r�O	=cG����L��$@��L%U���Y�GH����]al���w`���t�����)Ž��[�N�tSI�����w��ɛ�8�!�x��P��_zt�.��whu�իI�f��c�n��C�_��qa����4���M�"̥��ͯ ��Sۮ���M@x�i������W'�7�{<��T?�|G8n�������#����T�A\6�-��mֿJ�B�w�M��?,{ݜ�I�*����o~�M�ᴽ�����ތ_$�<��%VzI���s<���_d�q(�^x����؝�!��X�yHUɮ$�{���ӎ��,x����!	6���Y�4���~�a�ir���S��I�].���S0^�"�A�����Ozi)z�l�\���R�&�l�J�V[���.��+�"��V���\9���̫�ɮ��_�|*`�Y��j��=���Q�-6��F=��-�0OS��Ͻ�y��OP�0ꛃ�ޫ����#��:[(�.q$MX�̚K!�tY�$"���|	k˩pXq�����56�Ѝ�y�m�1B[5O6�._�@%0k�v���~�0܂#���H��j+�QB*J@��]�P[m��+�����\�e1�o�Vd��-hm�xw U����E+����VB�>�I��Ҳ<[�49!�B��)V���������Gyjx:d�,
0ʷ�"��ٳ��߬è3�3K���wsȏ��m��,%��ҧ!��}sk4��r�����ڭyn. e�x�8P�UlȄf�l�Fg9V1���v#]u��B��e�n�I�o9�~�1��b^F��a4��R&p��h���z#c��ꋱ�_@C���^�V�;o����*�������I�.����U�q	\�r�\wy��K��,6�$�!o�5��h[�]��potZ��ze}<�}��w���52�Q˯��8Z��m��ȯ���8����n�t����ru�b%�����?p��aK�&N��8g�ޢa &ٗ��F:��ZM��])x�D�E�/���ۢ����a:@�4=���5�����j�:�+��A���t�8��a
`��)��7vy�	F�
��6}|џ�P�������S`���O2����/�q΃�i쎨�<_+58��H+q�e�T<�����l���mі��!M%�[N�?Ym���@%~�k)��g���bQO٠�&̾��3��SzX}W�"Ř&�$���kl�^-[b[�j��\�H�*�0?���#��(ɭ��j�T��J5\5E�7vr��?�sŰ>ƃ!ǉ?�I�<l"Jo�����Č�P�&����i���7@�:��ɓ����[b�ׂਖ਼pX,&A�ȷ���E��#h���?$*2��r��"�H����
j��bS��:+ �B�>�!ݖ��dx\Y������
Y�Ըݢ1���̜c�PV�5��/�;)��|��!F��J*� ��F���rǇo^�Au�j7٪�!ↆb���i�:���""�u#�T��f&��&��u}�Ȝ��@�~���ӆ�cy�U���L>~I���%T��&3����=�I.�O�pz��+<
�>�
�{;��803/�#��9Xx?s���Uo���c-*�Fc[��b*It9yK����Lc���[㥥Dy���V=A��� �f�3
��U<�ISD���O��9�Qj�<�G��\/!�٣�ݑA�1���%zF2���zD|�v�3l�wZ�����6��5�׉�`xr�O>x��+=�F��2������|AS=q�e�� �v ���Mۑ,4��N�2�%�4ư�Ni<��B����`g�Z�����A�~_��D�7��GN�.��(՛�����h"g����	穌�ި7��y~Mvh��7�s�ru�6�E�3��Dmљ��m.]c�sl|ms-�6�z1��l{ە*O8��8ū�x���KEG|rQ�_���FS��&��H��u�(Kх�@�ZK��6��4
��N�]8@0�J�Y�(���K�A�,1T�_��}�[�R����O�#��I�K9^���N�!�􅒨�(�[?�������b�E,h(��ثsN�9N�#���ٹ��$R����4f�55�uwjc��02��s!S�S�tSdf�b�Ik.�
H-_ru7�C���fLו��2�#���֞m�����F�UB��a$PA��$�{�v�����'�l;��[�yOE�~!�׭��m�QE�Ԯ��i2A���nk�t�Q4h�Ϸ�~F�g� [7@������n�����)���_8�*��M{�g¦]�/�5�(סg<W��y ��E�A�"�=�q��[L�Z�AQ�@�JL�r��O�+vDZeS��8絮�p4�裹��6ba�J�d�I4�A������%�md��� ������l(�Nc�NX�`ܒ��)
K�`ӏ��V14}�	֩��s�pjS���T���|���2���$.\����f!u�I<r^��A!�8=q�c�8Ǝ����EE-u�_2[UPf�Op������ ��y��� o��K��#����g���Om�w�!0�,L%�=#��%H��G[���>5�t��~o����{�+��5	��/9<}�s�-����qN_ۚl<�2|�ľt&r����{��d���t2���v�ȷE��舏�t�,���V#���<�q�^��F6{ːw]�:k�i4B㗉��)M�3��)�8X���m�i��	�mm��m����G֗s>twV&�?����+%�bo1�t�i�q�&��<z�d�閧5�;4���^z
�����ho���Y�O<gӞ�o!�DO�p���;
��ޏ��5�n8\��gH���Y@�u<-���g�$}A d	8Ȫ��R�����`L�	@�~z����xì�;. �~0qj��=/��Yw�j�?f�Ie��`B���q��t �*\^ԁ��o�� � X+gRk � +t���������vCj=���WN�M����CH�}+�s`1](�g��>���`�C{�W��7 t9v�^�	�ї�PifH���T�:8\��_�4���/�N'����� �sQ�b�3�f��^�z�&�Nd��0���]�=:��� ��?�l��Q�Q%��h�͘ĩ�<oPm�rz�D�d�_U1�l�՟� ţ|?�<uv����h������t���z�c[[^�>G�]?�7a2}��ֽ�K��%��b�<��H��U��T^�Jq�n-&�|?��C�r��j:9�æh p�R?�a臥�
HH��MM}�6�6��__à�e-�����c�����ufӧ���=�~"! 4��D����'�Y�b�|"1`)u5�k/�$HpPy�)Y��Bu[.}�f�s���W@�/t��o��P�rKj����F]*E@E��ʄ��=�W6!^�N�!W&c>c ���$p�E���AW1��z�p�+�ar��
��R��g��5�ϓ�;��Ë���{rJ�k~��t�p�O �#��Ѐ��˳��-��:�O
�	o�4,�������)�Y���K��s�.b������z 9c��
eO k@9&���
��㠲4mh����y���A}E�[���>�Pz�߇\vo�X�
��'�<8D��6򩭹��v�����h%}|�.D�XMC��u#���W/�&4)��h��,_;� �6ۇ%w'�A�=�A�2'W�j�#����w�傖s�Q��ɖ�O�dY��T[c|� �꼎vV��v.z[�~Ie=qxXEz$������r/O���{J��HDLa~zX��f5�V!��6�Ք�B.Y�J&�A�۾]+,�
����,<�T�����]�ihK�b"Q�#T���n6L�]d��n�=����^iUػܧ^��Yr��\sM��ͷ7K�TƘ�=q�ւ~:ʧ/��W���>J&Fx�0�������-�m1��~�e��a4@ߋpvRI�0P�,d�o�Q�vN#L���-4ǯ�p�k�+�OIzGVƂOz�ǔ0��n�@�Vy��o'iZ=��X��`���R8`/c��f�*�Ā�Gj�-��8����D�4���хӿUط6����{2b�8t��ܬ��x���*t?|��-L���Ʋ^��GɥؗIޔ����5�!��Y>j�a��j�b8��M,ɟwp�����}���.�>8D��vl
��z�kv��S4�it�>��DSa���g��i;���4,�.9��*d����`8���=Na�C�vl�ša9ޣ2�oEp��F�g:� �����h�1��`,�'*51B�P�����W���
R�2�=�Ak��>� �d,D��� �\.��5ԣǛ��Ds����ͬ'j�~��`#��C�Hy�A��#�����c������(�l����d0e��#R�Bυ�K���p0X����n��kk��Q�;�#Q��	IQ�����)�ܰ� {�o��Mb�ƫ�ͽ3%��&�<�bO(�h!w�-�l��o��A���/���x���oO�y۱Z�"3k�B䉦��,ٟ��F8#8e��jrM&�;ȝ�
.�N[���t2�<�S����D����D�;�$�����g�_��qh4������%ALҵgZ�]y�d��9  l?���Q�@vYx�
k��pK|��.j>v�"�j���1��si�"-��k��ܝg'�a9^bW���`q���\�S�+�"^��?���aŝe��[�����]���̷y����轤�N��ߪ���=_���W4`��ap��R}���rx�? ��r��3�*5�$���|d�ʽ�7�el곲�{o��zA����
��Z��Wr\���}�Y��FͰ1��E�ǚ�F܆@��n
�Nn5��y�k]p�����R��Q��n�U�<����l�.��iT�,Z���g��0����}!Y}�ӑ�|3m�u�ܘp���-*����W<���1t��/N"�>����ۢ���?z��} ^κF�(�����b'f`�Y�Y����v����q�)D���.�\#ej�z�X�q�n�����J^�Ȥ���e8�AP��l�;���M�*��_�
qɞ4��ft���+���������w ��E�U͍�qu�����A{݂T�b�1ģ) )�d�Rtf�j�����`��N�~��}'�Lk�L��5�)W��x,����H��v����?��0o;�9�`�%�Q���_)�!���ꨢ��lX��z�H��(w`!Q.�IAc#�.X���=��@�k�|]I�oo�f���l1n�2J!ڥ�z�a�H����й�t�q�I ��z���d��o�w�]-X��@�o'�t�E�؊냺K��/_k#��U*Xm�i��Z���X,Da}��� ���O-C�ĎG��rݤ�l����N!fl�2�~3X����з��	�v'>��?������0!��`E�Oh��傺��@ND�$�<�@��ѩe�z�d���I&eHH���U�u���^~8��QUC�Ҟ�K���2c	�^X�'n��dnH�����p�5~�H>���y�1i�U0�HO�y8!�N1?3�;,_�$�k�AQ����K�㘪*l"&n:m�y��l���-����z`�|H��(�z;)>��C2ـ��$5�L�l�s�����-��\aU��ŝ���Y�b\¬+}�R(�o� �)}�*�o�_�񞝐ҫ�QV�z�e�\/�E7��J����l�8��.�i�z�Jh�6a����C��[N�W��%������ ����D���L��6P�����σ�T)6KuJ�i��E1����3�^�� u،�P�kM5�&�o�1�jz�ψ�ܵ��I*j�p�Kɿu
�����J	xn�To1����eIHZC=֕�Bu�eqN��G�!�5�_"�t�D/�'d����S�O��MeiO�Al�q�8��w���AU�h_�bl�l,W'��͂��qa��5^�[��ц���=����:Y�2m�k;���Vd��H��J��?��=q��L̃.�pv3�I(�u{�w��YU��Cd�0�D^�$X6��:���Qic�m�p<"f@D��%�L�g�������	��}DZ�g2�i�J��AS/ה[TkL(�3�<u�++m1���U��K�l@ r��	���t�l龐 :�����6�}��,z�5����1Zr!���`CP,�c�!�������G$2��_8Y�-��	���RIH$�@�1�C�<���k͵��=�좭��HO??>�?�^u� �� �%���t��W���M���E6{�[�9g�
(A��k�`Ƶ-a��%��#��7e���m���``�QD�Z'~w�������T�T���=���'}tgIڒqڠ>y���0��%�B4_�FR�G�e0;N�1s�Ŷ�{~�۵ꆯkb���:�7*@f�Ά���kX3�\'mO�[b �U�#A�hU�J�b).27�\��%��.�Ҥ[#�����X9�&�(���f;��L��G�
��㰑
�{��"
I�P7��'<�!�{�p͚(JL��aڪv���ƿA�J�с+�+��Ô��'%s�ߚ��p�q~j�i+TJW�0�C�ĥO��ͷe��W�s+IL��he���Rd|U�%�Ƒ(��Ĩ�%2��Λ�ƛ�b��},�3BHY쾄l�%�b��	���W(�5mb1j�kA�Ҙ�Q�M�Q{r�e��c�J�R,�z�jh��!�]boq?���N_�iYF�B�6M��/#tM����p��Ӈ/�E�j���6�%RA{��o���AW�n��2֥�#���~��&���ۦc�mY����nCF.��M����+��%�YA���F��H���Ft-��Y��lݟ�݄ƶ�"v[��2���l��X\-Q�c3H7�Q�]����4��-���o[�J���Q;3;`�g8��/2�h(&�O]+נ�U�+;���MH��\څnx�)�r�B���]}����y;�M�e�����*��V��0����;6��$���K�L�Ɍ��Rr|���W��y��IBcA�H�J�SS{��~0��H"_�w���e�v�?6e�At�A^�Q���?���4zI <t��?I�&�&W�D��V겟
����������j;R(̯�C͙ݕ�Р�A����V�Vݎs]�yl����k��������)���v8Y��R�L�%�����^X�U��N���5�����~�G�]��X���IW�	� ��ą���$8=�p~OQ�pJ뎮n���F�#%2z��`�pa�Xja�φ�jQ�O��\�ƸsA�x	W�B���7\#�i�[������! &PU�2w|���
�*�_��j=�Ӈ���iO;*n���~�)A�^��z�����G.a8���h=V1<��@PtKb�>���+s���4M��Q��o=�n��n��ғ߼3�Z�đ����|$Iy��[��] ?Q�Җ��M ֔�c�����cJܠ�M���mUo�=�T#(醼f�\yS�n�t���uڒ/DB�r&/�_�Y�L�e���(k8}��u]A��(�.̒��]pU�U���1�vۆ%�g��@k�\ ��ga���F��@�e��u�S�O�������8��dz�XZ�IPr��z�5[����	 M��7D��sQ࿫H:?˴������q�r�3���Y�c�;�x��t�7��xڰ���U��^���s4 ���a�z�Jx�־�c�x}�=<�$�͡�j�2�l�0�NH�W�<���x�.�XH����E98�_>1g������Z��	Al�6�F�	F��l�&�DR����N��}Qt򴔂7��@���(��s��?�#����i0V�2:ބ����I��\���ba�S�����,sME,*�!\Sϼ+��,������� K�=���N������MW�$�����Ud0����z��2lͯwf��:��1a�%���f�0���)$�l#�q�H�G�7xTb�g����\$��`�1�p��#N>ʮ�A?����o7��m��h�J�zR�sEI�y�l������q����ț�VMɿ4��2�c�2�T���'J��[�]�) -�v-g v�s�3�0��-`�ShQ4�Z�_���D��ky3pI�L�ɱx���#fz�Fͱ�������
@���M"�k��v-TV��׌�n7�����t���w�����6��">z4�J�����IY�`X�*��O���P,��א$�$4Cw�	�1"�woC߷�}�#8�lų�]LAN.�W���#3x'hE��!Δ4�����Ew��a����]T{*g&�`�_`�e#�PP����5��Ao_{xO7�2�-����X-���1@�ւ��>l}W�ՠ&ư!�����	!��[��A3d Ob��._��xOvr1,�Zr�U�ؾT)eȑ���������>BRL] �ګ3�DnӪ_6lC<���qP�ٶ/��j/�o-q��ۤ���G1{�;x5�P�U9kIj���s�7w&�nD����C!�؀4���xpW�1����Wn��-�� �A�������G��I ȼ�6��C��Z�%�zA��L�Na�8�>���|��W�:�q�J�;�t���:vZ��r
����Y� L@M�䗇��'q�g�
�Y�MΉ�&�����]0b	�^V%'u�t|� lC9�F5ͱ�]��3�K��膫(�+�Z��rw��8�Zl��J�E��D����w�N(s#�7Lڶ��Y�d4����}���D%%q�i�yD�D�;��P͆&���������2P,Z-e�H���?��)�q7|0E�%�ڵ.ӳ������,����H[�Á�����)!�d�+c��
�'�G���|����߂���b!N��������t�/oċ���#�VVv��z�����a�
��џ[���kK��H�k���2sʲY	�����,��� x�B
��� ܕ�ԑ���3?>s
�c���#�AFو����a��l�Ώ�b)�ڗG���V����M����Zn�ƌ�?\Ap�){}v�T�M�]�g���t�pU����V,�${�8���Er���q7�
�W �T[����y�07P,p9�l
W��B虇�
�#���~�o�N���8�BH6e0qC�b��Nx���_N�?��1��+�=j�@�C�a��	y�Z�=�z�~``�o�#�K���Hxyn�Z20ݠ@-2PX.:�$�.R�~�,����e�Y�&H��ݗ�b�/3�������y�,��A1�5��4�Mv���J��@����J�ڸj����VSp�	��E"~�
�2M�1�n�	�!}�sD���J��!ם�k��^�|����8�˛�����X>}2r�n�����G�q��ʃR�z�V��N�n���b'�[Az�N�;���r2����#��|B����xfmW"\t����	��z��J~��8>���>��/S�`��.	��`��샄Wz���U���"��K|�`^,�K�F��p�I�:q��?���8H�hĶS|T�{E7��l�ŉY�
J_���6!�R}理������l��~�0�Gn;�Ǩ]���]����cvA5i���rr"���mr\����@��%5��9���~Ր�D+n����g����!��`QvS�%��M���1�۴Q���|�@bP����j���_PY_B{{ߝ�?��	0`�$dw�t�Y�c�����g��8��i�i�j#m#�0.�$c��E��e�5��plw���جb&�#'�H�Ů�3x�2,�q�t��B�Zmu�Ҁ��V4����ۍ����Rli�`�؎*E�*��SuY���A]��;~�ߖQm7�&��*�͸���58S&�"@_��3@�,F97:���Ξ��+����WsI��=���M�q3�h�E����2U8�1�>w���kX}�>��캞^O�h�m� �fY m��K��؇��U���p	�cl�/����8�������c�\|s|�������gM���--]Rd���s��ȴb�A���I�߃�q�{ƨ�/ˊ@�Ai؁g��"0�@Ǣ�m�D+� 1����*�Ru�(�dزl@h2���Uj)V
u4[o�I�f�%Z��p�07{X��߶�ߖ��;dz&�\r�7�^�Đ���<�Y����r�B� z(��{��P�U7��NL"��=}e�
�@F�[�BpK���كSKG��:S��Ƿ��|�8N�6�r���o��gP�X���	��e�pl�El۞�\D�����t�,�,3%�V&�e�X�%`��h;��hĆ�}�:I;4�� �Kn�S������4+�>/��s�k����uɼ?���`�S�{�Q�O�ޢ�9��_ �̓(�,�������-�e�y��X۵e:=g�����Bi2SH��BCѦ���KL��1��q8V��A�T=�t��y�w�
�����9d����L�z푖6�Qi�B�0|�d���1�dXx����3W��j��U���Fؖ �y��k̴��JA�'x�rn�y�멝VC9�Uô�YfEe��e?����!+�,*�Ȝz��}�o�:��f�7����G�w�y�����ɯ�Ѭ3 '=[���5Z�<Z��QtFA��SքXP���<�K��h����rQ11Mi)V�oGb�6��<���)蚥E�T�l��%F~��я/�9�	:�G��L���_0:E�dXU=�N�:�/���,�|�0倠"D�Bv�Z��B���k4�Ɋp����� .(����+�]�����rrW���S�Pg@M!Z��=��+8��0��i�����YO2m��H���8�v,pn�_�X�e����i� �5
��@�6
���۾�}�>$5���q�U:W�7;8��5'������&W/b��$ȸ� l�����%|����&�����6rQ��O1�q���M����<,t���u�r2H�h���c���!�Q���z�"p�+�Rwl��S�V��U^98 �+�����(�8��\	V����q(!��J��@$ T{�*Kt������������:�iu�+�m]�Y뇮U� �I8�D�&����u�{b��i~�K�S��xqD�Ӷ�}A�r�_~������&e��{P_n�ÄQ��Gh�!4�6�
� �l�l7r�jǦh�s���ڬ ��0�в~��VB����K�}}�;�2L
m�J���! Ξ�qb�"J�4�0��M@aa�iU�@CkI���O�$$�zYlG����5����IW�!v�ά����baC~bh�Lk���)L	���i�_��(�(�x��,R�j	�#��0���d��z���I����[�#�k���J�s�=Vo�D}�_\WoB�8f��Gr}z�"�A�h���Ϭ���O����0�>��6R�����}��)��$Y�m^C�q;��5L�?)����j���qN�'���[�R�o�7�W赳ix��i��ɶ��=��A�>f�Oi;�$��ƙ��r^`�O���t��s�Dn|�b�(��A�����y��X,-'A��ኴd�a���	y��8vѢ�4J1r2D���������~8m�A����ϞD�g��_�3�t����Nt�l��q��Ԥ�'Tq� L1���%����vhd.,P��X�������ŉ"��SF],u���d�!'��FV���O(6��hM�4�e'73��s��<�qQ�ו�]ɻ`���YҦ�Iݥ6�u�������Ɉ��׈S�|� �����6&o�%+<�^Ih��2������<P}N��J�`*����y�C_�R �#�A(�(}6<�����/�ǉi������Wlf�~[��������yO�x�����) ��Yg���r��#��IES'�2F�	n>��X�/��Ft|q�w�Q�jL
�6^�c�l��I�9�
I+(��Ӝ�+q���m�֟���R�-��w:/�A��V=�w�I◺�~%�7�u\P0�?�cQ�3	ae	H<�oW�Oʕ2j�ԯV���~�{�֖����N ����;��t@�{�g!���������렧C��=L8�2�ڽ")�\\��k~�.\�v�e�����HW���m]۹���_��+J�=�2&U��$"��6-�{�G6W�I�P��Ndmg�#�?�\�� �2��FO?��&%�Mw���� ����]C��FQ'`VY�`8��2%4�)���Ǫ�̪�eל����-��h~ɧ�H�2�� |�c�݆�U�ɽ��J��K��[Xjz�o��J�R����6�*ƚ�q���������bb#��r�A�G�!&f\����}X1�0y΃=�vh>�sv� j�~��=l�d;G�,�"�r;�<N'�S-B�Ԗ��j����'_Jq,D���}�R��3d���6�?�rR_Q7"��&��\C��yR.B4�ʋf��>q��kC`��q[��R뀋K��@^���k�o��W�6����$ɕ_�N70uE+O�%j>lIɂ�GZ�����vt[�T��л�B���k�����k��i4��_C2�4[���Hy��c��+w���|��.��BT�ѧלb4�/�kl�I�~?r���(5f̘�#Ą��$�P����6���4P��*N�Rr���x�#�!Cs	������	u� ���"��c���D=]e�^����[#�E^����T�}���l�E=B��i���k����g`�zr�<��@�:��5׈E�h��`�����'r�D�q�D�l`j��O]�w����<�g�j��y�vG���kYH����zѧ��{����0�U�}�0�ڗY�x�zʚ"sJ�@|x�2�l����",�d�V����ϤG�j���VŇ��՝�?��O�:�UKl����	U��C�z&��W��<Յ�m^���s�|p��>8��ŀ�iӠ�Y�)$�������|0�⿍2�KQ��4r���w���f�H��2��M�&�)�VH(<q#�*N����6AC[@@m0ˎ@��܌?�۫���9��nf`�{p5.�?R!mTD��Jpѕ3Aa"��ꌯ*�Kn���Y�� ��ݰ��}�����B�#[��b������/��pg0����H�L"�@4j�Y�Z>�������l@�4W�~��4��&�q�XL�o7�kj~%0e���&��al���sA���m�溣��d#�<5w�bk�u��t�����c�z�O"��il3���c��{���m���	�"��Z%ڗ���򅬧^���R<Z!�s_��*�Ë*�a�$�P9�+�f���x{��]"�cu��KwҢ/�)�Dy�qxH}y�r�}��c�4�]����ň�Q2�K��%��cetbq�;��-٢p(�Ro���g��%&�W�A��4��[z>��n�/�m���m�C|?��3�S�u�p0i���s�7i�4�Ñ���F�hg�����GfrV�t��dv��_� �ERX��B�ᄧH-//���y��)aa ��km� ���&�nFR�z.m0��T��D��~�,�a���,
��+ȱa��er��q��47�}ߟv�e��V�]�x �F!nz��D�|T! WR�Ǜf���i:[`5�4�ј1��s܉�ܩ��B���]O�����r���+��[P����O��ʧ���wh/�(��؝y�rF��{��"}X���c��va�ŕp�V��e.,��( w�V���(�RZ����[�ki�b4����n�}�7�ʗ�SE�Q�Z�~D�;k��zH��$D���6�3��*�bYlƭ� �c��c+͢!3./=P�r�깙���̛WA�����µ���LR��� �:
�n'�"� ���=2h�.,Uaл���o�w�d�U�P��:D�_#�g��I쫿����?��'/��g-#4����樥��'��,$���ɡ6����Ҥ^���������{@S<�gH��DW�����'��9"Z6�lY,D:+>��E4�T���%H�y�F�!Q/u�L�D�[���ۄ1���/^�9�T�D�x�[Q��R��D�mQ{7o�F����m���o�� �q�e��2◊����H�r�!RT
�̢� 1�y�'/i�_��@W>U�q^�oރ[��t9c��_��@���<'��Qul9< '��@h���yU�h6ՙD�QU;�n9棲�	������n�x�>�BO�2ۭ?���?�֮v�n�c�𒾽^ܣ�CdO]Q���85b�Y�6
'����l���Q���&r[L�2�$Ȩn�Ń��b|� MO/�Ec]X��3U5g�~5�
�w����Fh6��t�0�0ݵB��]�o�_.�̚D6u.2�;�ן�@����}�w`��vJa4r�؋�>�h���D�d(*���K�p8G�n?�b��z�O�2������'*h��P�;��n�7K���LJ��x�_>�ߤ��8�f�Zw���@Jn��rԀ�̞�
t]��,P������d�c�����s�������O?�B�<�5R�N?�,tV��qc����y?���p����]ʴ�ʫ䭡T>��W���+g˃X ���]-�4UAz�u���N%Oe����l��=��2��	��L2���w�BT�`/^�"��G�:3�<Gq�N�2��' ���_�(�`!M��h�\^K��zd�O`�v�^'3��DL�ux-n��\��'��p_2k�f�qC�N%%���.���腫�Ɏ������39~�	��\����� }��eZh���D�3�t�����s �I����#��#�Q�?�҈�S�*����2�9��<�0_}��k�_�'0�����|����'[{�ۋ�c��-\[!2��3���7��}E�v�jQ�[��B�,Jo�{"<�P���o�0<���:��O�}M�`3X7 ;5Ҍ��P>>�6�f����T�A82_��8cHl�@N�6�V�j�_ے1:�לk�2b*����4�+
�j̓I���s�;�j6��Vr8����0����V+����zq4�:�w�:��rn�:����^`�.Ғf�T�����^���ǐ�^nߺ����J�����*%���l��թ�m�fuV/�ت�9�gmtnѿ�T-���t�2g�6�|�z�N�g�����2k�zI0�0R<5���aj��f�W�g$e�ȇ�#��kڄ����)�G���0�ț��1N����3�dZ�)E���kɊ.�Xwkd��F���(�n�����!�Zč�:�'����uB/:*�m�7�G�����Ϋ�	6D��*��5\O��M_�>R�|�4���˜�K�a�n1-s���ŭ܆�XI�@��oGD��@�u�0:Se@*��E�пQ�/���h*]%pA�m��i�1/]ZW�ʎ�g��/�}1a"�RM�ן��!ѧ%�r�S�nR%���J��5�%
 �,�eH5��h:pD���LDߚ�h�a�e{�F��Y����Q��2�����uY�Ή$��8��gۋ�:ܮ�!	�q��ɋ��k��],��:�l��H	��E�O��ĭ�~_�	��N��mwj�31���H�S�"r61�((����fΰ�7�u<��<�r
:"}kiZa��H�S�G[
�q�}��)<-6�+D�HDL�Ȼ�%ٳ�NM�V�=�5�H�
����up���C4b3l�O~!���~���x�d0�Q�
J�����e�TM�ł�ڜ�Ddz��R?e�w���e�'s�Y	��S�ٜ	R&�6�V��^�i(�{�#�D�%+��eLU�DV�ga�x���d��xT6��Y$�0"`��]�4��-\�X�� �]C�z .-_&r)[e(pN�ɤ[���#E��D��2њl�zM�gvml'�$.#PhH�L���Ǔ6
Λ������z�����2����r��D����u'�y?Xg�����s��JJ/g�:�V�p���[b9�"h	��U^��ffb�
5P8��37���2��[��)�F�:*�+
^�0%��i�/�9>2r�Erw���Ƽ"YD9�}5����H�{]B@@tB�i���� S�p>
.�6�G�p'?�3�!-�@}��a�vs�8��o��U)A���~��ҟr�̐;v�n
�� ��:��q�9��� ����.�h�|��Ap+ɻ��k�qe�^�(�M�a(��?8����ߟ���� ~��f�>C-'��9��;�������A�Q�|0,^̨'�	�z|->-��=q�˰0�Q�Q�j�O�Ӥ*��ٙ�=`��m��*��� �O���m���!�/Ы�؛d%�����7W��`X{9Q��BrIR�O|;�="����J��$5?��\&)^��ЕB���CI�����Vf�!M� M(���­&!�A��j.�2l�.äξ>|�;�ԁ���巾��D�#_��(�'B��gE���\å!DD �:ua�i_�)��)��(���0����]�7��N�ۅ2�	=l:W=ܞ������;�j[��W�Q�'�
;׮���>̪�7�#�E���\%e U?������Qԣh���r��� � H(�8}�"55ZB@iq�u�e��h�1�2�gf��5�+��V�����}Ϫ��ͫ�)R;�����wא�5$�̫ka�"V��>���j�n��m���v�xL�K�b4�Sa�4�w���,��9�%�&=�Cm�ɦ��)���K�e��B�ޓJ��^�G�!���um�Ad�{�j���ǽڻ�N���T
��pKMY����J�i\�C8�&�
�� ��fPJSN�1׶3n�Jb�.jx�G���ڱ���9x�4��_H4k`X��yʛ J]��2l��+Ԗj�2���T`B$����-cA3g�j.�0�RG;�u{a�i��WNw(EtV���BŮ0�m��z?w��"o�YIv<�63�����j�s�R��y�]Ū\�qX*u��u��Ţ��)�{!��u�(��\M��L�%��ȯ��+.��H�{7F	��@�qvZ�˅��^�ԖH�Z�����^ގؘ�獅���ި�_�v<�~^���g���0E�N}�����U��2�n&�98z��jpA�~��`���o;Ȳ�і��߱^�QidXhD�Լn�f�fK�̾�<gA�5}����ǥ45���YE�q���&5�%�}J�ޥ�$���S��EZ�R@6`I��3��u��yw�B-�����5,:��ڦ$�Sx4m���P\b9&��p����'@��Bրq_"��(vnUZՙMF��x��6����dw��)�w��|���8j��$*�}cI.?|'�ͬx�!{����ԃ���0ER�V�WQF�H��@|�����Љ04��킃?J�E=��N�Rs�JW�f�t�G��DD��ܹ��4H8j��x	+��̥.T�W��jI��iE�6\O���������чX�̡B���� �j�,H7�Kd3��Y���?��H�D��f+���[�-)
�����β�0��[`�X@��I0�o��Ʉ��K��on�i�{�>k�	�	�5@�u�4�^k($� /yc3WT��L������0�JĶi��Crg�J���u~D)Bj��7Ե�m#zs5���	��V���d�ż�J������3ӣdw٠&
��l���,���";n�&q�aݲ�n�@ZxK������X�Q����rH�H�uV(�,a	B�����v}W�G�T�%��+�j���8R����o��f
Hd���|k�C�0�7�+R�l< B0��dc{V�,�v7��"
��+�\1�y�(�q7���*�$��� C�c�h���tc^z�Vv/4����(^��8W����>�]f�ȸn��3[��Q&���Q����f��v�@�����1�ת3��I7�ǝ����S�	�>�C_��*E��������q]�*�-�G���Q�ؼ��������3(�W{��,���ɪ>�'����l7���| �y�bΞD�99�_9ze�P��,�V�N��$�R�4@�g��S�<X*�!���c��4�,.a�|�o��
y:A-�^�d]�׷[��Q#`;�`�n�(�Y���_�m`TH�V-Tܭ	ۭ*��V�w�]�cվn	M����@K�\TK���+����⫌�ׄ�n��y�{q�2T�{Z	��n (O�;C�-O��2���Ǐ�N���?+��+�֮������԰�0����/P;�.��CR4�%?�����pG����F0]���ҵ��7���:�̈T���0��	�Q��� �冽�� ���ۋ����fȡ~����y���7���t�����>?y��R�9�'��4����UN6��<��qn���8����9���[&4�4v��z+g��i��5�5lPt:���>S$�ջ'�V\��8�^`v��_��M�Ȓ�
�/��M�fu�s��;`f�d����0�P���@�Q��s�>�ɓ�l�$g^�ȫyiP��	���[�г�����1��7ZZ�X�~���#=��xĠ��~��;U�4��k�;���g�4\�_)��y/�^����`Z�G�ɽ�\#���__�^�m$ƺ�Sy��0�"br��:x(v������t���6Xw�r����5�,.b�����w�f��V��C�Tα�g@'�F�'{��vX{ج*ut��Y~.N ~�*W��~@��A�趴�b�[���X`y74����ޗ��g�����m<B(�{�s?�gX���]�^��IB<���X���p�BSZG�ox��M����)���|C��c>���v���1�Q)�r -\�V���T�^]�nd���f<��QbD��8Il�ӡ��l��Nɽ3\nnP7V��^_YQ ԇ�ӎ�<n�c@�/�yy yf$(�Ä�82J��ϰ��D�����ԋYY ��&������El�����(��&�h2�	�::���'h���G��8���T�k�<��H�������R�m��NE�`��w���SzA���h�Ҍ�}�'#%A��0�W��2�=+ַkG.�P�lǟa2j�oώ"=>���g�7=%�A�kj��-bn��ֿ�����g��,A�&أ�:C�OKi~&.K��o�j:Jd��טbӛ�@�#��]����h��Hh�<��BF;�>��DX=�a#�{L@�M����%��{#՚�
,�m�E,M�df�x2FW�6H�(�H�Iئc2���qC�#�F���vE~��s��8�x��̵�vq�M�J��'���z�����|mUe(1�1�U!�hl\i��W<��$̇=�H#���z����~��|�5_{3�������i,!��>��v��<��S��6��@IX�U���C��i��	RH)h���!A\�����rS��Ь0����mߔ17�U
�;'�@]��B%�P-%�moEp�7g9�	���,S��Bb�6H��.'���ٱS���(�/-!e�r^�Ł�-��OU1�Q��Ł�w����d�����F����@Ju�Ovsz��[���Hȣc.�Әe��:md��PHn겸k��裹@{8��4��1`�b�,�v��W=����n�㈦�z ����p1un�M�z�~G?�����qE�Y��N��C
��h_����7��j}���Rߐ�f���I���'��Ꮼˉ�[�b����m�B��-���.`�����_���q^�݌Ϛ1��X�V�g�,�O��� ��~cj9\�Ec9�f�(H��}�Ր����x��9�m����}�d����Y�����k�mmW@��8��&v+e��u���{��y��3F�'�ޅ�oZ��3�؛!#��
(�������~8w�݁��1�(ٞ_��<uv&����y�fIb*G]m����l���>2�E��*`�%D����c%i� q�>�����[��!���1����A����D�T<��_�� >W�W(iё	�q���g��ry���J@���?�S�׋�N�9g� ���<nz���}�qG�%V����#ܘ�e*�3T��vv��O>Vr�Q����#@��D\��fV67�5�X0 �L9���#6U3ePe��Y�c�W\,#�K�ܼ�ɍL����@����Y,KtB�������x�מ�+nUb휇��~��	W�Ⱥ������uKo���0	E�9�S㵷c�K3ܩ�p`%#�22����7���-~BP��V�&���lV�a�c"b$䰘�ăքt.�m���x�X�W�E`��xVh�SԠ��͉H�:��`���u�3g��k��P���'� �`�({����[��M���^���ʎe��8�4ɧ����;
I��#��ژ�%�DX(G���	�V�6�v!C�� ��U^I��k���ͮ��vv�x�����ܛ*����F�Vj�y�'c��W���ՠ�'�Vm���/3�c�Oy��݄ho��H�2 =d��F�D��"_mG�	o�u��G�x-��V�;��dZQ��=R0���k�N0���(z&��G*�6�`�[3�[hK�����%�\А�z��R���b�����7]�M�g�}���Ex�;��+�[A�$�6�w�t3��͒�𔵁#|�*�"��!�#�{�u�lzPֿ��L*X���A�n��w[1xz���B����>�񌋉�D)'Xз,�}����|l�C�o�`�>��1��b�Z+�MѦ���E��Us������ M����bi�i�� bQi�����V��%����<����^��呱ݮ�A�g��8V.V���:��	J�I̔�C��頭Ը7ci�������,W��M��r2�.���\���ʪ^>�?l�ڰ�;Y�*�Z6�qXs��c���Z�-F��8�>�ԯn�,��?x6?��V�p�[_~��-�� �J;�z��,�{��p+�'�b �0�fcӺ��]��+A����`�*J�V�Z>	���KG�&�B�K(��ԯJ'r�]pߑ���]��`��vB_�����<ce��,��:�z��1��R�5�M��%��=(/Zc�Xn��`9�nGN�O�l\�S;S��S����j2���4�l��d�:�x�Hl��{��Hv�s�O
��y�U��b�����έ��]����wg�EQ�7�:��C�9j#�����lAm���7��pgѷ��d*Q@k��j��]��LF�~�$(�G|R���L� ����e��X�( )�L1�8�=�f�a;<��Q��0k��9��x>ߑ̗��R��.���\�h��>�cA�}�5I:M�����B�w������ �'[��]�	4�R�@e�	��`C~Es�uXP����,��d�L�¡�
�Zۻ
�x�T�0D3���MQ:;%��{��KZnnٜ]���.U��0�WP�+���2`h?�(�8�@���.֢"�� �_��D�fO�8 �^l!މ\ZY��A��A}�>{2�.:�tP1F�yLAA��.�2r\ I�T=w�t��x�b��X9�|��
)�b>�&�҉0�������Dy����!:�����ʊ����4�c<}��6�]���M_Y�h��$���>6��v����D��T��8:USy��e� 
���F��)<��{7�J��3z���&j�8S2�2�܈�@[צ�_�c|�3���&�X�lO��ۛ{�rb����ʅa�~��v(�wtϞ�;{xݑ���Eu��˽�aaS��Ѭ���#��m�6�=7��Kգ$>O�ĉ�����AcQ���{2�Zɮ\)�}���N!U�y�u�C�93�;8�+ܙǈ4Se6��G�?���R���ǔ $�����n
`�ˀ����&�v6�6�  ��I*��3S����B�x�,��Q�4.WC�*��}Pc���<�VE8wHq�.�r�2��/}4XH�ؑ��>���F7E~\�@�s^͋���|ی�y�í�0�9�j3#�Ԗ� �#]i���}�\��\p���	 �{���_!fc�O�7��)ψ��N� I�A��7p�����f�s�`P�b��	<L�)�k��!k����׭A��uIz����6o���r����>R�OI���"����?�g	��ޤ�]����1�w�UoaZ��x�7o����o�e ����g =�]���a��*:�%w�+ь�-��B᫓��֬jǦ5iЛ! b�ߤFo�"�1����pe�>�$#8���Q���2�ls|�Z��0O��N,���O ��G������<����4ś,l�]�|_Q�R�M�;����Z���\PeD�[
�1N����rDb�oD����#�[��D�D����,a�js�U���6��,��qL]m�á|`��|��k�ʍ����/�I~D7��5��V�!��(�χy����z�h�G��S%3������I�������5 �rmx�2�	���9��xZ�� ��cn��eQ;��_��;��mF���m7×�h��܃j􆫠;�~�:Y�ASw��4�i-�u���z�!Q����q_��X.�>�
ȩæp�n��n�Y���U=/�Je�D��H���D+;���xirz����ptvk: :#"���Y���Å��_j�\+��ˀ���Ȱ������P��VR%��&6��Qz�ҝw%���!��Ԡ�کhN��}%]�-uX�,��S�g�Cʇ��J|�w%#��+�˹W���.��N��A���b?U�X�C�7���d�/�"�3E�O��ac��k���QӍ����m����<q�Bi�l�|�.�����u�4�v��S�-��R���%����q�� �t���8�_R�`�O�'��mNr����"X�x��@�����'lC�H��ν4���Xf��3�:�9��(����	j�ӈE�%��6����3�Ɉ/nX�e��LFZ+�X�������`�f��=��N�!�mT	+X�>5K�v����k.Ȕa�9�몤�w���b��U$�>'`1Hv��J���|��>6�C#�{�x�K��}%�����Yk�O�xxbi���lj��,f[>	�2��8I�O�
�}��F*��Ɩ����	�ƍ�j���$��@h��q���Ͷ޳��%c\���
̙ضN�J��d<bT(:h��dAY��"�o�71�MO?��&�\X&g��R�'���m}�2�Ry���{<^ړ�A S�L#�EqHZB,߇'v�,JX�=�/j��c���̮�wa���P0v�G�Z"������l6�����[L���J�ɘ\�&z�Ā�H$I��H��݊�|w�.�=D�h^	���'Y�i�5�R>�,�7q�j������V[a��s%�p���-u?�n��+=8ge��Z%�e��]��J����-�]32_���:��2�a1փ�@����{c:�-��jA�DD��<����8����Z!L�ށ6��V2�$������V�t�$p.���PLasy�v� o-v���G9a_��H����_4@�� ;�������?��3=���\�9�
�>�:���z��b5S�b�5|�h�CP�)?tT*�c]4�O�5���H��c���7��$ +K�y����x��km$�)�bs⚺����z�{��s�xt&O�P=�$��h}s�u�3�l����As#����J�]<���J�Ѝ��*[�[��"ұ�Ԫ��ͩ ,����"7�l��_~?��ģGv)�{N9hKe[���z��6\��}�_H<����#B=ܚtܣ*�7���%s�	��#���>s���=�k�6�=W��񸻬��H�D�iN�?&��Dy�<ȗN����"�9��O��NO?�wR�9���b-�Z�#�g��O�&��>��tY:G��v&����RÀ�J��ꋫ�JwS���� ��A���df�������$�P�i�3�4�Y�j͒u͒a�V5��t�O�(��T���`(��T���TU����c��Oe^r�ğ�,qt�P���
�ڛ|��𽮆���be<���ڐ-CFP;f⑊�h��Jx��!N�[�����D̼����u���*m�Xp�̆���c��ËO	��Z9�9��>��@���<�V�3C���0�n��Y��|�LC����Ie�/-�"tpN�K�B�Y��ǁ�=�1R��ŀ$�b��9��Å1]��z�G|��9{���劖(1&0E5��jcb�bI[$�MF�3�b�%�,�jۉ�rZ&�lc��-gv��W��a^:T�q{IiSųdC���#T��Tw ��j��}�W��&�6V�b[1�j.
���o�!y������nT��2T]����=����������(���6jf��"����Is�g�����fS��(��/sҐV<W�fZ�b9��AC{�!+���WӨS�)O �m5��-<�	�Q&F;�m��e+I�o�_4$�[��h?��Fe%�\�|��Wos�)�7��VS��`.��N��D;TVB㈶@����R(������!lW�=}��-��L(�sP��4�u���ߗ-�̻��g"PYQ�gߓBf.��������u��2�sŗ:yDD�}K6*���)Sژ4WI����9��hU�j<�P��R@T�i�M�e7`n��W� L�K�:����+1d�?�|nR7DUv>���P�KFe�g0�C�"V���]���m �C=RJ��7U"@:���\���@�m���FZ���s �P������#�XQ�+o̴���U�(��(��HgA���������*rԼ���E��5eW@K5�e^�E�Ӱ���#bl ���DJ�I�$�tW�k���um&/N��vv�ٶ����HĶ���&���W�^���� ^^x-t�%��N�	f��.�]�1C7�-s�aе� %'�6�\�Z�a\3zN#ȉx���1Qlr�r�vͼ�{��Դga�Ȑ�)� Is�ڡ%:������++~��gb��v7�'*=w�A���-�j!I��j��P�T��E 1�5��V�li'[�\PFG��D�V��g��32�,��޵�]��tsh��V�r\C��甛)�|E	�e3��yq��0ϱ�m�т����0bH	]���1�^2��<�F\<�&�Xh`_o���B�X��Y,�.��TQaZp���4�7���ЮD�rDn�P}ID�00�i�s�sp\��Ϙ��S9��ң��"�낺Jc8ω�j����R1)D7������s���@��W��i����d������Z�=F�Vb��o�>'}����0Hdn�<�8n/S���%%1����ۗ8+�O>��+ ӟ�X9-�I��	8Ɗ)��?��$K?M���i�ŋ���ñ�j�py'���%-���'f5���}��k:��&�s͉�Ī��u�|�����
x�>ǃ;�_�)��a��z��L������xI?+d;���s�MdE7����bP�0���-�Y���?�.��V=�����!U^g���dB�b5\�O��yV[��Gm�Qp�dG�f^�Ao�ΫE=���㳥�$3��P8�Mj$!-մ1�=�v�T��E���3w��oC�(�o 3)��A3ٯ��3/!�zޗ+c�����v?�AR���^ �*�b���R���n
�F�̚UbFT�A�����<Z�+�.ɢ��F��!k��(MO�З���0{R��^�o�ss,���|��x"7��n�^�|Е��wv��G�1�ZwǝuWd�L�Q�%�}K?&
�'��O$���,ч�t#�O��E��[�<��*�������˵�]����֍t�&�m���MњK�8�9�c��C}?A��7�y�ytS �*��5/�ǣ0U��5fg�硖ӹ��7����+�¡�����Aq��D�2~'��Z�_��p�<��$�MP�3Yڐ����1�A�x+i}�w4�a�D�ho�VwB��G4�+� U�*�1��;ړ���G��D��0L��U��ܴD������|�W1s�zD���U
�*�B�4��Kgt&�h@X	߀�&�ӗM�râ��e�uW&��,̒QI�lGD֑�#�*=w<�#N��iZ�c�£�w�oJ.��/����hN^]��yR�*H��%�|�	d�S�*Pl2.;`[s9�v�P�|�9�	Q�������G`"�+�Զ6>(.�U�&��v�����r,*�~y�����!�.��aź�,vy0��?�-�Vi�]�o,�iF޵օ�"���Ŕ��,�P��p��_�ʗ��]9��i��Y���#7N#+�*l�9w�$/�~g͸��z$x�oXLH���vaUxb��!���/2��껞���|y���� |ﴯU���m���H<蓌<H��Gۙ����D�HoS�sfCDuie1cY���<�_�������F�顊�l~��ß>/)I���+�������qo�Bz���e]G,S����M���ɛ�38��Lo�\5k�ì�4-dB4���n`s���eu2�F��Ɵ�D����*����2~���b�D��-g^9�(C��hhi��l	��"{�x�QQ�('�kޣ��.#�=.����h���F��|2$��dj/�o��b�U�F�W[�&�/��R�*:�,��ъ�
�0e�GTK�%�}a�_�vO�ހE/��i�/���m�(�}����l!�@Zi$J���L�����s��T&��eZC
�@<�kn.�_�8��|!h�R��Daq�!�P,ھ�e��!��J�B���ר����{��f��W�.%��f>_Ɖ<bͲb�t�865�"�c붕K��
r7���a���f��vX�5��Xط(ўAj���	�i���7��\�����vX�{��Ol��;��l�sE�+����1�� Mq|S� L-��b����j�w�p����_r�~�:CTu7k<��Xw�	Mo��Z�o���ԟ��� /��D�`H��;p�Z�� ���0�:�|�S�&qt���;�8��ׂdz�4���+�0�?��Q�s�X�5_���
#q��)&Ca4�.q�Y	�\�Ut�����*b�w���ϑ��o�I3�^;S3�B��F���4�/�d�R]�m���^�7�ϡ$�-Ж��=G��/R�)���o�~Hzp hх�����S)L)���qm
��W�Ps14��|ۣ�t�!�&����.��L�&���S~	/�&�	6X�!�'MH\���gDB�e:2�"0�w���L��W�\G��,����ތ�:M�j���o�֧r�bpw{�I��C_��_�����:́�Q7M����Í��~j7.gϹ�� Ng���W�`E4�!���{�ilC�����c�\`m	�4�7{b����$s�ɀ�Il]DP� 1�Q����t����/Q��w;�ㅸ%Yyh7�S�l�%+��'�Ҋ��]φ?�u�s��W��5W�'�u��@}b�ˠ�9�u.GQ�(��0�B��% l6�[4j�KK*�Ht�}�0tB:�2�t$�
j�?s�U<M*��Ͼ<����~�"��d�&ߔF���qZ�$���bD�q�����#T���Ҩ	k�|�بK�v�"G�7��q���8]I0a��L$�/�k-oQsRs*���T�Yv&<ޫA����6/(���C�7/����yB�5'[<�Y
���l�N� E��9�"}3N?{HbV0��e�0�|T�*b����G}�Y�	���QЙF[��jm�r�h�'7� �ifɴ��L�,��"*=�Я7���c\�)����(8�8����!~����\}��<0�u�����ѧ'�����ƨ·�<�tKN���V1�q�Z1A�[|	l�-܌���rmR�@�Q("���Qv��lE8��k�����۝��C�D�;߭y�B����m��-.���[c��d�-�@C���(q�8�.c�����D:&�o�K��Y�S��[m�K�.�r\�V�M?)v@���0P45�9E��h���J��;8��;ȇ���#���;�?'�j�����=O���,&*�,5 S���y!��]�Y��Y}��kv)C��$�D�T��u��E�յ�uF����x���趏a��.�a�c���1b[��yO��������to�����ML������$V9`��b�����U ;����O��X���9��3!NX���!�۪�����b>�{��D|?�9:�w�-z\-GbA��2l�.8��.e�н�O9UrEW�w(���v�ˑD��fxR"L��-H�#O��#�CM��I�iMi��-�i��eb!瞿��>��ͩ���$�?��R�iO��a��»��S_���Q��(��'h��S�Y�H�]��4~_!�8�M�<�teMUH�xU<�4��YI�yc���ǝ��ì���߯)xl)�)�8��td.�U_�1%�H��~>B;�
�ې�;�'p�ĝ�ޓ�<颉'A�#\5�o�6,��.'���P�0��}�9�M.�����@��9=Hu�Bo���OÖ��|����6����'�J[{y�QH"qq�x�����8d�-��<G:|$�Wb��r�U��w�k���
JQ��5��$�@ ��M�D��8r<�'��%�5�?�����(4O?�I|����#xX��b��$C�4��fs���D�?���S�yEt-��N<[�I3�K��UVN��̏�
�@[�`M��$�SL�~�1ɚ�)ը�'��s(��%OB���yܜ����GZ�mik�詐��ޯ�������PV��Պ)����%�w���z���*?���:^xL�e:�u0�J����ū�~@�V��IS{HX/�o���\o�P\ő�ٍR۔������>߀Ps[y��yg���d:���lR�M��y0{����V�i_�B�ϙ�S�u��1�g�������W����^����h���������$ߵ p�2����5!�<�x��g1��=�X��<�x;�	�aFC����`�l���
���B��F�?!6�I��ج���u���.�=e�(E�����8�La��ee��o �\aݰwQB�o5�_ه�ᄱ/�r�ᠬ[��Ƹ�4Z�ƣv	�:��a�h���H���g�f�I'�J��D�Ƹ�h���Kv3p��="@K�!�D=i�`����ᶋr��b���|f��[(��֧N�uӥF��150�7�d�t��H�c6���\VG�7[6;8�r�҈�8T�9�qH9���yc�9�.�����vU`���Ԍ�f!�=-eP�X\�����8߈�[UBU.U���>��X�y�<i0b�	�-������=�Y���.:hA��-��T�ڰ���6��.[�$<��9���Y� R_n�� *�H�U�2v>�YP��@�
?���5��H;5M��9YoE8�O6���P]K�~.zr|��T��V0�\�}�t���{�	�xh�J0��&�x�R%�m4��5R�;EWj��Q(KɰsO�����@*$��r�]$:+Z\����i򿨚	
��>D��D��r! n�s��~�Q\�A�K����A�%;D�((�~�����;��i{�*`���ڑPg�h<R�wqc;��ׇ`��h��N3��.�`f^�r�|�7�3B��n(^>=2���]��R�j�����gVhx�Ù�l�=j=�>�Rt+*?42�� �;`�;���Ock'�}�L�4��.Z_>?��*`H-Q����kcE��b��Dxu��yqav�������ۙ_�gw���z�(([�+�$�����xe�<���Q��
\���C��.��:��f�0E����r@��m���N_�DҎh�vY�L��~�0�f;)-���L��������� �-�������d����@���v168A�J����� �ցƊs�<�u�E��OLW�ۃ�����L +�c�e���P���%`H���G���^��Ҙ�s���3�����E����P ���%
/��������.H�B��@g+�������ϱ�=��c����:e�T]����F4ch����ټ�Tԫ�2Q?1���EU�
��l�@��4!j�6�{����[k.��}��	+�gɅ�s���'�����<�VZ����V�Q�Y�А�2J~/���`%f����ʙ,��i?�\fO�z�"1�ү:���Z�WK��������?=Ȟ�J�rt����
�e��-��BG�|�;cq��.���t�k[��p��@{>W+;l��,F�ԭV�s�+|�?ѝ�qr�4����E��˩���o�l2&��4q�
��_Q{Y��=X��?&w��6�"�w��9<)���3'{^^��q`�;�G`G�I\�n.검�B��qܤ.riʭ~�w	�O�q��k�4�I
V
���i���c��9 M������O� �立j����ʦ}��0��ru@ %wՍɩ�]����\�$����1�#��Q��`��S���^�/���F�X͉[*5����?�<��3�G<���Ʀ�w�Ζ��1bL-��9j,�����y���5�;07�a�D����6C�|ߍԹ�w���epy�56��������
]f���_���x��5أ"Sh�͸F���<�۴kj�<�JO��5��e]ǛZyg|㷙 �-c[�I��1�d�M���
����o9� s�L
�"C���.K�Vvv�����]�M 	��n �)���
|�&w�DIOh����[���/5���14+؝�w�� ���|�kMm�=�J3.��C��э&��WCqR�wj>PXhZp7��n>��q�cL���O&�tr��su�>X�"�Oܿ�~�GM��������`�*�	��c�GA� �AV5;ym��ְa����:Z\s�At���Xe%�<S!���m�V|:�)!�^��_���ۋ�����bI��oҙ6�w��xn,.L�`t��{S'|��3(�0�J<BC��ag��!�ix�M��4o�^���DЈ�Ny���j�"V���j�u��`���v��:G��@e�猑�v�!��-�IŔ�M'�ρ��JZ�%�'̔�zB�;����&��Z����%h5������ �=� ��çY���d�	��s{0�ަ5ڋ��5|	���������(���Ґ������n��B
n���btA�/m#�A0�N�0�9�ݙk0�����BK�b.�6�%���+����܊w~0��5��p� ^�Q��s6���;6�L*�#M�;h�a$m|����S�Z˳=�%x&�-��v�K�k�%#Q��NO����	Un:�����ؚ�.�1�XF�t����h$����������Ö�=ʠS��zs�,X�'%����%�'x+0�C6"�&'Y��$&�x��M=�]����J�DӼ/6�gǨgE\��6����=�Z�Af%��	/�N9�B4��&��Y��;��NEY�ћ3��,�U�RY��K^�:�aG�0�3߀��L�OrGX~���9�9,��H�3DRk���d0�ި-3�xH��z�a�:	pea�V"U&[+AH�;؞�[,�;����=#�z%���y������%�B���o���\e�FԪ�)^~h5����=����<J8�D��^��(՗�Ԭ~w�̲��i^�/�x�O�^5(�^����x�r�VJ�kAlk� �=�@���&������5���J����Za|�q�$�(R/n����z4@����<��_��4aǛ�w�Cƃ�%���FC�&�)�������]�ecwq(8���&~�x#��X�J(m��%�{
���\�[f��T�"w���}t�O�k�`�������ٺ�c��]��q���#����95�>0�����֊��K�B7��]ۼz�:R=Q�/g���w�h��WQ�6��/CY%�@���s��?�E-��f�����|7�y��>Н/>�T��W�DE��X��SN�� � o⹵s�,B�ԟ�f"D�J��c�g�M�q��5R2T�1~��#���}2|N`�<7aT�;�#X��p�f�.b�"��d�C�n���l�-���c+�7��^3AE��!���p|wN��S��LB����!m#�);W,(,������NV)� i\��qM!�j�Y�hOUmƃ�zP��/0౐�k������pD�Ve�ކ_p�Bϼ�,�#�Y��z���1vW����I-�m d��ǜԽ��(vݩS��xos!���B�ugJD��`k&���BciĎuZB���ƇR��,��4}�j=�$D/Tb7�=q�0	D��h`t�-��d#��~'`�fe���YF��H��0"'
�:-T���e��j��qVw3��&� ��a61һc��z27�aK�^���]�E����;��2\��냼	3i89ܻWCU��7�5��
+�B�K��	G�����V��x`�:(���2[�ys_��e�{_g�D�[�|��!yx ���n}J�>sU�?yg8�Ǔh��S�`�;�:ǡ��Sn�)i���N^�>*H�k�]�*u��T2�t�E��
�ڪ�P��D���pǳ��0A��FG�)��l�S��|���-��-"��*c��2�8D�ҝ��Y2�g�z��X��k$r�/�\���K���͌��3��Q{��2[��g�������I{�T�eC��Ñ�������B�ֹ�6�ٶ[����Y�iņ����IDc�]�t��ܪ����ϫ����O%��CRӼ6�D;��FgB:�M�p����2[ߛc�_+���;Y��_vyzm�	goI��R/hAoӄ@$`�����	IY3�6��!/E�m�G�Q��"��6�,l�i�f��L!���9w�j��	\�k�}E�MBuʆ���T�/���O� Z:��8H^�Ra���e�s��*��eWhך�&H���53��,ߩf<~fI']�]P��}�hg���|�T7����a���KL��ھXb���������{��X��M��c�G7|�Օ��V����v])���'!�]�)it
 
NtA�H!0�s��i�����"�T��ɼ�l1g�-��}?��ӳ�|�r��à5G��`�aܶ�w����Z�G�BBn��|2���"����o��F��e�xu2Sj
��5L���r[Tx>�x��Ud>�k��j����������]�(Q!��u�ӑ�I^���Y�E��{��`�WC��۾�T���Wb�r���\g�W`[�lb= .�ȟ���g6���w=E�8��*[�����*;�B3�xL߄3	4�E�.��C�N'*�#'eW���)?9����t��kf^r|��;+�PR/g�g��A+y���H�a�#WH�P$L{�Y�)s"b�v4$�e��z�8F��- ~W�Sx����p�����٨��b��v��	��#�o;�-4����"1��t�b�֤�9��?BL�p�pf�r��k펒Vn��Q�L��ix�;!*Z�C\1�6Y��i����ї��$d�w�ΞbJ?7GD��j|��d)s���"`���@���xp��1�h�	�9�G���9Hd:- �8a�ë�����(bЄ�� (���Π�L�=)+@�f������fXju:��T�eŰO��fE���tb��^�#�}{�Wy+5��y8�y$-�W|<&�9KS}��d�BS��h\PtQ5�/��o�'Rձ���C�?<��0��A`�+3~�p��4�X����~��;���d�2���k�g1��Wځ7����p>_RF&�u$�:k���[�b��_ݕS����~��j�I�j:}�jJ�jH�.7Y�A��M'pڳĭ���.6uZ �ԞrA$��AA$�T�2󇹖�m
;_��E��G�G�W]~%���'�)�X����?����2;`mwU��z�Hi���pH�'R}�*P�b ��^߰�����S�Bİ�]�	j���,���"`l��Q�_�vb��h��u����r#"1����py�ix�2K�=\�f�j��t+Lƣ�T5"<p�}���u����YK��L���J��������;G�+]���\�7�.+�k�����M�/�������pL�oD�xؼ�[룔���{�܄���6ǋz�<��Q��<���.�$�Z"n>���2hC	�+uڂx$�JO��}�����⺡[��R�`�=�M��V�n���� �oM4s}p�)�:��j[͖}�//?�y�s���	{����N 5�H���{/]�+;J0������`|�6ණ�@sit5-P������y��3��Y�*��%4ɝTh�0fS�=m�3RF����1����۝x>Zh[�GE}�o��+!�tB/۝��G��>�פ�X)�ԽRK�Ij��A>d�`b&�{ʍ�w�I���n�d�f٣8�dl��x�P�+T�F'����W�@e�$�ӜrF������<�=�I�1@�zM�;����tS]�B�Y�h�b�h�x��)'*�vU=�u��exT?g�9/juc����_k�γ��΂��Π9��m��2���.��S�nι��J�f��=�ꚫ�3��)�vd|�������-g�LhMz(z��~�〣���\F=OS�$��#���|5�ɪ=�$�j��Jx��^W�B^�k�9h/�3I��\J�+i	�PQ
v5��⦁�#sސ2�hu�:'mg;ǈ�����9���@�#3�s�����i�V��b���}l�M��:$��NM'%Ǐw')��>t�����kTO�eV����`�6��w���HKgNc� ��E2BJ4�>�vr�rۤ�e���g̾��6�p1ȇ't0׺|��S' �2�Q�[��Cvd�\��o�3`�,Z�S �S2��5�ߙ���u�J�y ^Ԍ�my[-��j����.E@g���cZ��K�[����8�Ze�p�D�����$���?�9@q]��!�,��X&�~��Wո(�.�d�1�U�-ԫ����ƻ�SM���N���f(��0��5��D��{��k˘"�)(��&���Z�!��U�g��sc���H���6B_u��	�^���EȘi�"q/��K`����c�t��z1�B��?����ZN:���]ZGⶊR!~ЍU|?r�1Z�m������#�P�fɩt�''u�2a�H�B��̏ZtW�~2��4�	͇ٞ�7�j�Τ{D��Ks0}����_D>hD�B~��}�?�)��O2��S# a�I��N�F~�Y���dW��1�]�`pJp����APh{ֻ��4��v���2��#N��RZC�>Ѣ3$-v:�=^Y+�8و�yEQ�3����.�m^|�.ɢ'���pA\����.��&2Kd�|݊$}i��bH_bq��݋����MX{vP�?��g��#���?z��͞�����������nP\ͻbǳ�h��Q����n(��փuxi�KXn-6Li,�Jl�r(H�E؝�4��������8��m���9l��oh�~���Ri�*��5�~��!�uۮH�!���7;�����.;��oo��(޻�<r T]�ET2B(�>:�H����<+��qB�^,t��� �B�!����6U��T��3S�-��v���E���Fp\�b���#�Ս����@c+�.7fj0�w���t)k*H��� |6k�(��%:SuM�=Q�/�>"����[��K�������/�Z���u��B��>&��)����^�t9>Q���(S�^�Ȅ1ϛ�MD�W$H?�|��U��ѩ�Cگ�c�J��,}�Μ q��ȅG��V�㬏#~*���D�}Ô#��R�I����߮U�ٓ�j��@RJ�FE�]R}fE$����>���=>bU������{��ݝ_l�V��9� �A��Ιbg�
�w*�=<�E�O�6~�nW�ˆPo���"���EԪu�"��IĠ������J��r-�51���źyh�i��^��O�l6f��Q���5ko�8�g�y�;r��ui�I��܊ْ��z2���,N�_?7�g�X��fN�Dj��*:��dK�љ�v�@��c,��7�d�+0Kc��ʊ���N-&K�d�� "4������1L"X���(T��4���^��F���fK�7�X��ib��=a	����r�Yс��Z�:]�MZ�=gIF��{f�Ǟ�7�a����;F��n�_;v��g��n���mr���� �V�l���$L6�z��h<��B(3�i~I蹎��D�L�N�8W�=7���-��(0�q��.cnH��ҢM̃e�c����)�szǁЎ���$K"��y��U1�Mf���(������u)ppn?U��i�a��b>��ha��yE<b���FB������O�m?��n7�9�fSy�\g8&@W~���/����L�{�F��a�gQ9ٽ._Kb������bvQ
�S��7��w��1�&��M5#�N;��V����4����)	uH��pK���suE��ྑ�O}/+~�Xr�B�
Gؒ%+�"J��� ��#�]�z�����4�%w��P$@� X�l.�}��X���9,��)G
O��A���1D�ǘ�fɰdT	��O�J��[�W�S�TW��"b�@��̸Mͬ{�A�؆<�ĉ��w��iHǢ�
�3���!�rd;P�$q�U�uok���X���%/���E���{UC��O�>`�T�ހM3/o�خ���-ѵ%0|�E��	��~�Ew�M�zV���ϳ�}z��.�9�3ﲣ��[��=��:�E��%�pEd�� �OK��>l����v����=�[�(�(�����-���-f��� `=�^y��ovz�`�q�ڱ�>:�1�O��ㄫZJ҇o����e ��@���2���*Ԃ�?EP�rP�n���J�%�8��Vld�ܲ�@���)"�ga��ɲ�B=������x�7GAf}���E��lj��>x~�3�q������X�)UW�}L`Z��5
���԰恆Π�%�u;��)%=���k{3��2�-�k�V�#�KS���q���YđwR�E����'/!���I6��5�V!lW��k+nD�	��,X�"ڴ�����I��3ۮ�]q�7�d��U��޷$!�+�ވحa�U�a>�����}x�L���IT�o�p��ռ+����)��d58a�8�OE�W�>��դP0S�H;������Mw���F�D�8��j�b�)�NM`���Лv�h�v��pݎ�����JtE]��j��$�T����c��CfWJ�6f��GM���&#fAc�yo����6���]���ޢ�7l�m1�*���c��1Gl�*�X`Xu���6�Η%�(^q��,���� .t�·����5$@s_l�e�ͷl�Α�Q��h������ʗ)*;Y��Qf��\��Lx�W�,D�E9��0�'��W�B/�e)T2KC���
I~�ǹq`C7�r-��@��9�_��	3Y���zDg3��h)�3��8V����x���_Y�رa<�&�N���N����~"F�����������"�w��Ӫ���E��x�EM��CQi�9ɑ=o5T|~'#�&)|�?�?t��h>~����b�m��\A�A�/Ȳ����M�Q!g)L��l�t��{*�:fJ���o�K�>00���'.���In����LXa7�z1��?�O�=J߈�[E��C�"m��V9��k9w��{�#����h%��?DS-Y��{��-$Q���5b��F����^2mV�SG�#�鈖?j8���`�!��7�A�T�|^�}\��ӋA�rZv\}��n��M�l����ɂ�N�R61~;�u�k���]����@�R���ZK��l�0h���Fk{:sD�j��:՗��NV����Ez�P��	�Bt�(�o�ZZF3�oҔSw�Q2r���d�����,�v4�Xt���SaM9��,�"�4�Gq�<��Ad`�*,O�%���e-;�__�^:�]�G��tcWlZ��i��
�qi ƫ�b�����;���=
�������jb�u�!��|��ډM���qL�2�՜y�ٽ1��y�qE$
A\�Ʒ:�}H����#��O=��	�Bw�` ��)A15�(���nd#��#�%o5���<8&�X��J���$�Z��!� �fC2(��mʌ�g]z3(+�Z�����!� P�!�,pmu�ԡ�e�m�X!qU��{>?�B��,.�qa��U^S:z*g��Fx�p}*+@a��#��KA2�<~�rQ� �0��Q���ڿ�q\��' �+�&ƌ��!j�6��
S�I�e�Y��C�l�QA���n�	��zF�1'q�
�A�X�S��ˎ.^��6=�SH�u>4�'��U,&���o�E�$��X�,*����t{S�jy�|a��06��:&��,�"l�b��Q�a���dy�����Cb�b�޺��f�4?$�>��<�H�� ��+��f`�Fv�7�J���9���J��d+���L��Ճ����W�����?VȦu��J٥��#�
�>�9������ΐ�[��z�rg�l�X���F\��[���M"��E���e��S2�(�&V���ʭ0��E!jhUg�6t�-g�,"�s��';|6�g�Al¨.H�N�^d4_:�Mo�gZ���z�لl7�Z����+d7[�v C_�vz~�mH"�Y�]��h�ˠ0z���>rt,��a��Ғ��$y�)�Op�V#��i (�sefEv���i}�)���;����ɨ��M�i��*��L��}�{�5����� ��n�b�C���BwDd#5Մ���g���z/z��1�2�㷄�Sy�|]�4� Ĳ;�v�H��*dA�YE��������"���3���=H���Ok�p+�+�L��\��Eu@�G"�N`}���n&�ޯ�����>e�o�[�f�Xwm�ɺE�B�g�i١���g�S�T�{�ȟ3��ʐO#��d�tӴ)*��j��iu���#�S	e8�x�q<�<�X��+���0[���ƃѿ�1�潪h���ms�{�о�-��I.&�A�A�,躥�����ߦ�����R�X���9�&Gw)HB �X�	��n���]q�c?m��/�矬�
s�v}Di�d<��@��+�CL���2��CUD.��`�W�ߝk@T�0\%(�S�w�Z%��������G��:�Ubb"�B��n��ɫ S��+_��\�
����.-l]%�$�n6�>�*P��΀�P.��v��Aģ�ˋ@����%iG4'x=�g���%�#��x�>�1%�	�Z��D��&Q�t����lM�8�\L?E�/�̓����i|��
�_���!b?�;ɩ@ӚE��[� cT؋�*K�ؑ$ز���y˓���C����^�d ��j����T��M�k�i,�F���+�[�w�� Y��q�n�Sю�v�;.1!+kT4M����	��ى���a��ܠ�3<���{|�2~��v���ד%�5��V����<P�׃��"�fM0����j�~C���I_3�#��L��f�B.jƝ��@����q��E0+9.��-S��Ǽ�!ؓ��!�%~�����&뮷gD�r(_\� !+���[���)/rg�=�GY�����U�z����$1w>��ڹ��T��>�ލ/[�����Z�O<��a��Ex����xE�zz7����,�������N�ԡ��ΐ7�Ԗ)�N2B��X\G�2T&���q��G��$4j��{����~���b�ҙS��K�7��G� ���]�(e_^��]��hC?%wS	{�'9f@)�J����ʵqt��+��
��IY���c�W�܃�_����Fb=�MTH��J�R>�닢�B'ְZXR̋�>�����(���*0z�E��?��!��l�e��c�r+p�M����"��.vw]�c�%dЦ/3�53D����`I%�"g�_dO���8�l�������#o#��Q�l�J3�Į�h;ʓ��ײl�-�!����,a�w�ZN�{�����9ZTz��T+�<�J�꒖�m�䟝���\�\��q�;n��"��H�M��+{䍏J/'K�Xs��l�$�9���n�a�+s����6Ϙ�o� ỏ�E��M�Z��b:��}�{�!����;c�Hݨl��5���D(cY�{=�~��Z�L�
���7wD%��R���#�x|.��߇���>�����
��i�ine�h�$�2�Z�"������1ʉ��|���G�

��Lw�Loc��$ѐ�Qê�1�X��w���0gOw�}���X��͏8v{#'�%�SE������,6i�@�	��^��_�����_����HpT^ۿB�����>�e�"1�^7K7[	���s��_S!���I���fȸQ:G���,���~�gJ�6�(����FZO_/%%$���}lw���, "�3W���v���R�,K�5a	�"�Չ�#>��*�%]ǵa,�Qg
\�C h}les(��S�H�b5Cg�j2#������0�=τ�"�>�&e莻X�����6�k����z��}�3Ot�+��$�����,XВż`�5��a��2�G����x)7���믓�b9��[T�����D�`��5S9����Q�V��ɿt�c!n�BП� q�ItɊŶӻ�lgTA��ǬkJ���%N�N
\}Vp���pӈo@����g�螡d�8���ӥ;-��m��C�V\P��0�nh�(�w���e$Z�x!�w�5��(n{�/95�\�QQ$��������gdۏe�Pe@����������A�O�b,��D_Mf	�BY�	�h���̸�?)s�ⸯ�
a�]�V���'��Vˁ����+D T���ψ��&���aÐ[ޮ7�n��͡�Q]�|�P������z���U����`7��O�6����m2u<ばT���јN.{P�+��̓Ξ0Qg;��٭����4f�0ħA�nR�'�|[z�wwh�z=_��B������:�,�8��MS$*���]M).ۃ�9�j���M�����\��:�`L�v譆�{Զ���CT50P�[;g�n���"g��"�&E��!՗NX��,����oC�o����^�yӞ'!��q�P����ɝv�#�]9p������Yy���f	}�����S��@��U}'$(dJ��j��ah6�`I�h��|��i�<�qڪ{���9D�0�%WE�`�o������*#D(%@L�%�Pm��QM�t?Ó�@�C
�~o!5���@��ߺ~O��]����p���!�smS4�B���8��O:Μű����8���*Χ�|��������+U�?X�$7��@��W`��Qᒷ>T���v��:��%i���z]�;s��T_Un�]���d�fܟ�h���Y�<��;�D;��wr�;3;�z nc�~k&*,3�fuYI�䢵�%�H 59��]Ĉz��fD���g�Kg4�*�������1ǌ�ʳ�V�zyH�����%2�������s���o6�P�	FA���e1mk���e������pVW��,��t���I������NǑ�ػ�a� �%v���r�Y�ހ�SM^2YZ��
�[c��_��ͷN��&�7�p\���ӮI����'	�ڳ�?�G s��p�uu�69�κ
�)d�"m@gBw$��mέ\��B� ؟f�����R�@p�,72}N�*��ڧ�`v8��0fF_��pi���6!!�#Tr�0������6��`"�������X=�]A����J��xH,+ߡBB)��X� �h�ˬ�
��t@��xX���kz+�Mv:7j���"3�t;G�A�5���;�:|��
��7�֤O��򧙴s�X%������C�H�2�Xi��d`����]4��P�wE+���Y����5HZ��4xY�+h���������;K���9�;yxWI��]�ˍ:����ڣ��3(��`�eן����O���3��,<��&���wL�Ī��L��Ƿ�v9���g([5���פM��Y��1Q��Ŷ�8��@��`�������Ϛ��i4���� ��ܩ�,8���~-mD��
.Bun�N����*�;D���!��f���O>vw%����L�"I[�3�hQ9����f�DnA(G|?��t�r�A��Lgխ�]>`��%k�介�7�	�=�zEI>�A��>aUcC0֣��-҈��C��1u��&`ѕw����k|9��D�G�;��{������4_����w`'B�_�xM.�6hu'�5B����ؓHn������� ��c[��,"{L�
n�V��J�-f����0��T��q�r�{UY�+c<3E��X�������a0fTG����=E��"�n��`FwG���t(ŏ�����慠�M�+��+��Ej�E�Y����4���!Md�q��7S|wq<�^<f(�g[(N��d�{�ϫ��͑H��*K�
��B�S$������Aߥ��Y��[9~;0��tĠ
��$Xș���g����Tn�[�YV�Z'�үOr��+�U�[�$�'��3s9ד�3����x�W��` ��|�ر�ޖ�#p�}0Ż�q��xk�-'6�8Z\��\I���[Ia����]7�9��Vty��''<��Wd!c�Uq!D��	�,�%��R�Z� #�!������$��!p[jT���F��>���Rfd'����L@q�R�1��?1V_�>��A�o�:ȶ�*W���zw}[�#N�$=�'�;ml�`6��k߽Z�ΊG�a����~���⭪%3>���ʶL����c�=�v��@�/K�#&�ީq 2�����P[X�X50��lqPkM��`\�C��p�h�fKSxXĦ��K�	l�u�6k}��������I����U�D)�����P��CnQq<<�׾��e�l\�Ѯ�(Xň��L�NhX�
3���w5.��|=���[UCA����3�Žp��S�p��*?S�8��0g$�%.�=�&�YA��{rb6E�����KX|A��~3��j:ɠ�1�R�<�rڡ�e=ܹ��dD��7��i�P�Z�܋��17�N|H.6T��I�p&�G�j��:�k�0,݈l{@�32snT=��R���A?��i ��;����ᭇ}��)��U���C!��c�������'��nl=64(1���>,�Q��l��|������s�Z�>�{Jb5� cA�ů4�`�a�x}ꡰ��5V��~�\`ݿe��,�vI�ˮ^+��ѝ�Z�*�������[���x~G��5[��Sv)TvBۜy�2}��-����L�������&ķ�R�|J��i^-#�Q+F���&(*�1��d}[s~w�vO"9�S����G��Хdťy��@�g��cJ4�-QuMp�V�GG8�;�����:���C��"	E��Z�b���h�H�Ǧ�D����_��5Ķ��I�#Y��V3�0�8�c�	9�H��(Q��M��ܬb��Au+;?��v���(�Mr�I�W�����zJ�0�F�	Ie�h�,��G3}�yX�)��K�(q��4�'ֻ|1`!i|;V�߲N6Z�x�[Qp���܈��~� �#��̷	(o�"��2�]��ܣ$�}|k������V��x���&[y��v��^��$_����J� �信rKvBG_�s��8����'��B�t-����l��%6 �?�>ef��аAS��T$Y���^d����uk�'�|�\k�Kc�E��oFC�w���+�XTe֒ߴ9��v}^ ��S���>���Gyׄ�i�����ʕ����P���ׯI�O���ՙ�ƞ�s#G4n�Z���jܪ1����A�=Ҽ�����у�w� Du��.�G����_n��,`x{��~e}^���w�?>:�������	M[	M�Im��.���L�N{�<��,�ɞ��i��Tk ���5�����]�ڟ��g� �L�o���3 �5v��	!.7��^�n�@�Ƌ���M-W�ۯ�dGq�H��1k��<! (��_��KEBe#)_�[�܇2)GA�*���"�ɋ���;.@h�M�Hܠ x1�D�2�����(�x���"+MArwT�d�����M��C�[Ի���b�K�e�M��wD�h��qV9|��J Y�kҥ����r���N��`��k���ď]����k����8�w0�<�|F}2��Or���#�&��[Zg"#&�ݸ;��Kt!*��/D;�y{��S]×J�;�+�,`��	H��JcX
���z}�]�%��~����QCI��6���}f�,w�����BF�RA��A��E���G`(��5�s��v��q��M�lHJ��s�ç�Kq��"|ĉt�R"M�0��4����dZ�,լߩ�<��E*S�+�F�`���@��H+Zy3�P=nR�Q1�ET[���qdC�N����f�}������>��OJ�V	@+�j-����$�Rt@6�A�!�F���� 1�� ���WJ����0Q��Yp�����|\̀ŇI6�����ȧ����)8�$�R�ϭt��_.D�i�Y2?��Q�-�4m^
N'��nk�{�z�x�	�Y�	N�؍(M|F�ˁ�L飝����,�n�!��*��ڙ��_�c�L�)7�#Ӱ��a�^��\������}�h��+�:��)$���*��Vl�Bix�S$aq-Du	�ڴ׶�#Z�p�:NЬ�B����U%�*be���G5~�a7��Go�*�G�? ��� ����#B�� �&��ҩ��/�5��9�P�B9$���������/�@cx�L��|A��\��f�%�{h=jG!;PBD��z�7/I�E������1}MU7b��p�Ȕ��;��
4��
�5�%M��&�LBYH�O��C��j��m �_�	.���UK�F!"����	���ڞ��6`�	���֬c�*l�|m�WI��.� �Lf�I�R�D��7��k��@����
�~]�J]8�1�+J�]<5�����d�B}\��N��t��*�Eߦ�;�5��_o�vSITnC���c��=mw7�2��6��d��Yv��M�ܞ��$B���e˲f �X�x͒�"[7�R��<��6�|�Whڜ���=�~\ZΒ+ޒ���n���~Z�L�,�V�2XQM�C���F��XW�Ya� �S1��{O����p���a��ߌ��]!�8���j��Z����z����G~�6`�:�|7���j�8"���P���@a��/�q{\��
��j��ʌ���<�7K�89B5T��Nr����o��9-��#W�3A��9-)��"Jh��
.}��`��9ӽ�E;�Z����S^��6�N ��}٫�}ӥ�0��-�K���׆�'�瓡ȵ�0z��H���qM/4ЪpM���z�j[b�R���l�l���3N����ZQ+v��@NDQq�I͐�a�H8���*�z��>����} A�^��N%W);I�P����p�YxiXf�?8v��͈�kh�0���EX.J&is�E�P,��Ť%1Z��,~*��dSES�W鎋̃���=7�1ț7�8�ױ���K��Ԕ(��j�Dv*�J���[;���.��
��Gܽ�L���}�� �N2
�J��Ȗ9Ǻ�ޮ�ˡ.�C�09��!�	^A|q�uˎ���6Mt��Y�}%�b|�d���3/�Ss2��C��%.�Vh�[H291�r�D�v�f���c�/�e�U�w�l�9Q�3�[��=V�.Y��_���d9��!{8���\�%��A������W̩�Of���A)R? ���V�	`����	٤�k>Y�Q��\���T�I!� �H@-k��nϋ0��a{�^]4�qnR�C���2�lz��.O�T�	l���C��'@V�,,^����k.���١V����]�{B��G+7(��0NP�r��P�� 	xi�{����=Q�.�-^�^��'�� e�!P����f��yw��1=z_���+���� m1'#�H�	F �KZ(��ͣn������@{�P��ٴ�� �"
,��p����@Ѵ�HЎ�����W�G�Δ�Јc�!�1�F�7�sR,�h�f��[����Ĳ�'�`���a�Qԋ�qA�'�/  L��xR�j��qבY��U0�
�4R�'B��� d����.A����c�$u�U��e��ع�qs�~��bB�]���o�|�j�%E��2��\�
��s�bՓ���X��ۓ�ʝ8j4�������C�|�F����@���ç�5��r
B����bĸ��7m���1x���p�����|�VtfG������F��>�� 1����t>ff����Co�(��nI/��j*0�q�-��ԅ���>m(���W�ޣ2�����=�<<�W���1\����z�>�ӡ��w%�Io�dP�]�N����m�ezV����� �S�(�"���gR��u�Q��=�%���|3�ᘇ=-��7���38�ٍ�ݘ���^p��&&���	�Q��۰8��%���|`Ou���R)Z#Zt/��"*��14�]bЬ��q�l����L�GKtŚ_(�;��Ue��X�5�Qh����A���J|�87�`N�$�)y9Nt4D��vUA�!�r��J;׋����':�k$�h�V���6`5п����Ee�\-��yaڍ�d��5
�7z�����#�W<��)}A�V�_#׬�6��wY�I�p��*�j+�8��O�e�	�h���H2�vծ�qu�I�7n8*�5&�$%�N��I���AfW榐v�D�{2I8�R�8�� ��8����5xU"��OLʹ�Q }�n	�@L��� �H[���������mי������\�h܍���?��'�[��2�KQ��q�r;�f�8������#3D��v`�S&�+�*vR}�����_�1y:	G�(���N���d?�m8vr��c�a��Q�1BJ �=�-��1[���[���tH�d��l��d�,D=Jd,u`sd��=���i:�7�|��Q��A�*%�#�W���QE��ư�@���f�xӟ3�`����Hd�Z��A�J��:��YR�g{[����F?��k��s��K��Wl�dǶ @t���<@��#��\�>V���E�cN�E��0�?��gE�̈́m6V��]��,$0B����n�𰌻\m9Y-t�?����B�L)g��b�Be�E@e�/�Kј��:����(0�[D ���,P�Ѵk�N7�����n��s7T⁘��Qd�ȉ��E�SG�5�+@/����n���-!GH^$�?�N�o��
�9f4]LT/���q���1[��q�`��Mb�Μ& ���qv%;C'�3��GV#R�q��~��y�Зz�u�ӛ�"�o��<�K�-@��!�S C�@����1��@�c�픅��������Ն��8����T�=#�H�0���pl���\�[4�>Q�­�:C�]��@ݦ��i�m���`+��qS%�huh����M�?q�V���*�.Ơ)���([�U��-_�'��P�Oܴ��nC��:�@#E�wWh��H��Y`��� �A�8��!/����)2t[aX��G��f��m˪�_#Ÿ#
~�p�*xjɁH���S�6�w$�� ��H�'������k��R�Q��̶o��s�V��㞅��2j���xǒ���\L�f"^�BF��|�C+*:���9�nu�{N+#R�sW�w��y�2%��� x�M���'�'���,���CA��Q����5�l)y!m6k��юf��وh��6F�?��������]�1���ظ:�g���E�wɮ��3��@@8�n���"EI�z��m�	�c�[an�?�m�ܢ'/���|r��=H�!웍��n�t���������$�j{�B*|�Z9��41`IN�hSU"H�3��\ix�]ڼ�܊���1YA�T��6�J��_�8k_�	4-`���o:
�'�zQ�V8�������'��7�A�I�"޵�/�H<ͻ��?�f*h��T�l{tA8�賺���͘�A�=�o�v�ۅ��6�2n3��e�`{�w�S
྿Xo�z�����-��A_�*67~�6����F���N���W�.��rT�#���\�ɕ�kn�)�-�j� :9+;W����p�*��ʓ��@�7?nRǈe��Z���5���mf��A�_��U�"?J	�*��P=ѩ(�u{�f0����_X���t+d*[ ~��������CQ�d[�v&��?�7S����%8�#�@
KL����жAsk���������h�%q�[��=
�ݠL�d���3�J͙Zn	X�� Xg�sG aQ�D���CC⌋�j��3��_'�,��Ř�#�R

��
N�[&�ס��,��W��ie�Fxmu�)c���N(Q�Q�R��+6q��a6|����#�J�i˴<*�,P�o7�u���h�1�_oG]xNO�a?���w �}��ӝAc�
B�8|_|�!�'/�����_O��x��fCm��M���Ś�C�Ը�]�KFV�+I12/��t�]��N�9��?w�];��:�AT��7a���9T�MƵ���8g��r;�	vX�Fg�OZ[S�`b:��ig%��H`ȶ��;���J��,��*|��e�7WT�
0�m��,*��E�5`J�>kl�F8	�8�����&���kS߶�0W��n����,g����}:�?��cx��Ζ6W-��a/D�񎰬��{��q$Q0��[�q���{�L׏ u��@̹/H�IqI�����inz��S��\]���CP?jW��H*���~���h�I�[&Sf�]Ժ�o�r����_Ci�eq�N��z�:&���S8F}Đ%�B�������m���a��0E6ۻ8�	��UK��FN�J,w��uL�X[#���+REe�,)h���P�,���<��,P=X9�~}�&l(c
�sɃ:L$:�f�Ա2��PZ�dh��:�S���j��w9��&�ڑ�}�D�2��pP�޾4�էC���_;k4��n�ж�W��`�x�U�}��d~͸�� ���A���`����<�ŤN]N�.Zͬ�ԳF؉f�a�=�;%����br��
������FH���ec�����;�^��I�v�@�ؽ���q�&{nD�N����Y@���]s)�{�i��~���vmyPH+�� �,t�L�,�hy^B�"=���<T](�����d()|6�v��c`�;m��/���y3K]���y�3��W�Z)Y5����!�­וg7�$K��ٷC�d�%�����>�ǥ:�a}�f�Y���^��=��ORM�nI�g�%�ZY�ڌ@���Q��4.	�� (S-����PJ����	��.��&a���:
[w�C�hGr�ԩŋ�x�:�߅p��\�
B8��xd�A�`돮YÀ�ř	��~}�
-|u�A+��
'eJa��&�'��Z�?��>� ��f�vq��l.13bڈ�{GqL��G�U�u����'4~\zd0#����ڥaq��c(ڧ�2{{µ�+�~i״Q��t�'m���ٍ&y�òs17�ٸ�>��֭PʻHq����ݯ����ٿF6\y�)ND�`<e����+ʹ�a�)BF�=$�]��ûtp�J��S@oQ�?���D�Ӛ����� TR�F��E�AS��O$p\��4J-KpL� ����-f�b�oz�=��6���A���}����t�W�9-���a+�'$f��^�<ڟG��^�1��pI������ˌy�7X8��Z��e�@�-W*��yQ�x��v���;_�t�����'K��U�,\EN�=�m��
��NI��$���Q!�ȝ��b�a��� .�ϰ�KZ�V�k��ӯ푍.~mn����&��������u��XA�Ǽt/�;︀V~��K��>+�oͯ�`e�+���k�J+�~EH�(t��<�M
u�-�;�g���a�*܂�'T��$|*^> D���rqER�u��1��VHg����7^�	�Y,$ '�Q�p�/�q�0R�a0�|#�Q��2;/�A�4ؗ�Y�y^��s�NL�ض�RZ�<�ʇ��®`	�����x +��'����}���Q�l���eT�������u��d��_@}�tbu����4�0�C(<nzȀ�:��HD�=H����s@k�1��T6�9x�?ʡ��i�"���fO�H��:�j�F�=����n�����"�w%��/���&������箔琑� ]0�8����W9+���Լ�`���.UA���3�>ٵ/��� �Ջ�{�Gۥ[�O&�SN�|�h�v���2���؎�+W������F(T�B��d!����(x�!�oG!d���A?�KY���h��?�}�����a�@
o���-���C�:���jUh����tRP�e�k�FQz_L�U�;�WO�98��������<
[��q������`�p���-=���&��pQ}�6�����t�W�(������]��p�Bew������6�����ԀR�\�67v]@�Ia6��9-�"�Z����KK��P!��T2f˿8��}�2)���їR�����aJ~ܳ��I#.�Ň0�^�e��<$���2��viEe��\N����{ �����T1��I�b^c�}��~�/��e �u���O����@�5-M|��/�;m�Ǵ�|�i��-G�<>:�Q�ܯ��N�3��U�A"��A˚1H�F#f�M�QjZ����0�抧}sA{h�,��؀L]jkᝰ��j���;����	����:�Hޭ��_�e�V��N��5*�+g�F���?��9MʎY���,��>�駘`�t�J��c��-�)i�~ vT4ۙ\/\Kd�n��E�\��b�n3s�'=��ī�L�Da{0$nm7�����S���a;��z��H3{�7J��h���ӥS�������.{���(;U�A�/ҙ�X�$�0��ct����AI$�,5�߾9Sd��,N��WNFť���T�^�����Ex�`D`hn �|kш;A����2C
��G�pZ�݀s�g�;�*�(�)�P�&��:��Tý�N�a��X׿�24��wߑ[��X2`C"��-�
��Ȗ��'���n���#�GV��|3pך�3_�\N�
�b��ӯ��z������W9Xy�h$Q���Ϝ���J�q��N�<G��dE �"�兼�Ԗ7�ѵ9�I�����r
)U�*9�8��m� �_2Oa���_�G�uso���Ơ҂��|��oK�`R�<*�bU���O5��/����*�˄=�������)�c� �v��où��|9G�P�Z��/�i��e�_��g��dLk�#��"���ha� �F�V�ι'k�2��Bx��nj@F�\�ﮕ,���ҳ~n}�7`�9K���������iA2
	=�Q\̟�=�r�M��F�Zg?%�k�'��7��Ϭ@&K��a_�Gru�����'�%�C_; 4�ȹ�1w�����;"���L1�$9�*����D�<N$M��ש���0�r.��|���C&�=Pp�c�˥J`�-�����<����yDӯZ�:%
�*ic��۲�^#��sr�P�p��U�{h}i=�(}s�X���� ''n��+��v�g��"u�4U���*$�����[R�*�e��П�8��b�\[�X�p��(��@Ǥ��ȓh8V�����n��N��Q��@��q�M��7����@�Q��x�}A��D֬Y��*S�'��Ǯ��ܮ�I`�mP��V�t;u`Z������`@�,i�9����/P��8�x/��ZV���:��l�!��l���]ȝ���*;S�����Dqi�3�Ii�s6��c�lv�#�nN	��%��P|���AN��#{y�D�d'E�n�����N� �9ɰ1�� ��*4l�ɨ��[�C���t|0K�!���ߏ�#��9���+��M�t��\>G��y�c��"O���곒D��Y�@8��V���cME�`z�dw�o��7�]Tc�׫Dߝ�- ?~�j����h��L�1�}Ϩ�Y:��/2�'�{!�=�{a~�ܤ����5u+yBB���n�A�qr���U-B��u�k�w��݋���t&����@_4P8��}��vj_B�����V����f��~c莚Gd.~<>8��?ij�,���S��7��{�����aIk+�t�zX�U�P�zR��T�mf01l����@V5	T*9�w��ub8��+�y,ʜ�'dKn��ham�i�6���H�챑���
��eS`A��ʞ�w(M�:�^e�ғ��{Qm��ܑ�Q �l�c�#e*�-Y
5=�U����6�d��wC߲���u��9���Ր.�)�U��mi#ϲ�_a���6��.�b�?�N"I��s�m�,_O�N�+ڄd �Ȼ��3U�L���7F�Aq|V����#|����L���-$OE�1��f1GN_�������#i1��}�#�0�W;t��Lb>:�]و>l�0�/��w�s|y��x6�U���C��r�`!����e�k%.��G��Cog,����R.V�"��xSw�{����+���[� 0ֆ�?� V��%z��'�KД�[{& ׻���������Z:p<�,��Q�h$D�TSGV�i���Vm��'w�c�&1�T* %��?h~';G���9��Ͱm⿆oK;���J��Y��o޾l���Ut�B5`0�o��}Db|/�=��"��$t�靠� ~�5�ej��Wa�D�+��ijjv3&�,�0\^�ٔS�����S�[�����8�ǟ�������sj�A�:zgu#C ��n[A��"y7�w��dTgى-��-����~.�_��x��0%���\I��LxH���ә�E<�E
�^��@�敹{�p{��xU��p`{Zy���4���VX�	ӓ0y���͎&3� o�+O����k��+{��ؑ0�rf���'�7�!He�2�I��67�'�������ܐ^��(r+���>X��������Y�s,�=$�7�3`�c���;`�?��s	)���f���Wd��B�4�.�-˕��+C�݇�W�ŵ�TF�S-_�����]K���`3�O�ey�*�b��a��$T��^�I��WD�<���a�ɗ�{��Ybz��I��xX_\��X\I܉��<� A��`NBQ�2컍
��W׃��9ex��G	m>\��5$�Pd�yǎ�a쓑��iK��$`�U��I1;��}u������l�  KIwK����Ma���J�<�vVښ�xk��0���=�qĮ�v�E�xG��3�$�_c)�:h�a�y.2_0�)�ٮ���:xP�������%�9���G%i�S�d=J+
a�ܳǧI;��V��.&��ó�˹;�-���؍�/�Փ(9z��˶d��?�I�a��m9M��e�0X��
r+��KeSޤv�Ud�<dć��;2m�����C���Q!�c~��tP�k��F�zXJ�S>6��=�}6�kX��9۵˘0uuW��OI �>M��.;;���Tjx?�����T32i����\	Y������Y���=C�&;R���F@M���
d�@HԳ��L �s�x����S;�)6���:Lqf��'w8�ӎ��a�C�R���I��� ��K@�_�{6�u�\�\i;z�����@�eJ!˟��,� ��-�����E�m��t�[z��^TEx��
�޻ߡ�/,�>�"���#�{�\�J}q������z�5��t�Y&�s����y7��\p��-��z�a��Q��ѢE�]��:o���[$��A<bu��b�'�{�,�	B����
qδ»�0��j��Pd�b�c�UV_��g��"1����>�e��
���n>�@6��ʿlؔV�CJF��e5թ�1"'��~��c�<ð)��N��?��׷>j<�8^u�9<��K4��b�2���e��,l��v�S���(9�U���[��0�������K���H\�DZ��I�6N��WDv-�Y��&;������h�#B83��;P���S��jχ�߾���0�gN��4A65H��
N�eX0ӫ�lت��5ഖc�Ɂmk��yK���"H�Zj�?jMy�A|~;,�ɆeS=GV�U^��	�y��mL.>h��M4y��<G��W;�����k*��KC��47���ޟ�C��')�A��	���j�=�z�I9"�J�Ȱ�,5���qY��[$| �@�Q�*q`o���u�r盍��V��¿���
lHg�,��䧾�V(��C�6Hst��#��������H��/�<@��q���D-	�z3�р�E�הKq��G���*x`Я>�n�2:�,[�����f���s"�d��[ҖY��&�]t���Ed�ϭY����a���N)��|�eZJ�S�[�-�����^ѓm��
���D��z�8���D`�V���͔ծ	�K�|�4����5��l�%�zohcY��A�8��'?�7����챾	i� ���U+��%Ke3�%�s�Aޠ�����֏ւJ�=�
��d#}���R뙜�57��u����Z��]��*�7%I�_���X�=�G�x;T��5�fY+-؛Nԧ��<�ߪϿtJ�,]t��Z�jV�e�x�^(�*�/�\�HS�zi+�]X �}�f}ȁ�����޻֛(h������5]w$<"t�D���!%��#C�haco�rѷ�?A�}�"�!��H�]�?2�.�L����
� 84>�ݔr@lD�V:#�<;��-n�p142g��eFv��*�5n�V9!��^V�\�3u����1��ѝ���9CJ74��|" ^���ʾ�L�j��PɆy�(&�С5c8߁����m���u{J7E2�=]�Q���B�IעT���d�~��^@K��+�8'	���}~��yc/ K�-����.s�NL&VC��_g���:��A$K���Qŀ6�Wե8�a8
nI����^��.�$�
���G�jƥ�����uM�5K��mY$�:�G�Zǌ��+t��$`���tE�}��-;VBP
el^V2�ʽP�;��˫0�YD��yq��)���Ԫ�Я����Wo���)�-ɵnx��p�.��$�w
R�6�5�'˛`P��I�s�s��'���u>�+F�<e�Ao��%��ǲ���n���n���Sr�ö�;/Գ6��.1���y����H�P��$ߌ�x�1�"� Ε$Ol�'�d�F�!�
p}uٲ����ر�"E�A����v�Q�5nx��*��U���~8�69H/.��m��5]  k��A�NB݁�M���P�-������Ѭ��Y�wA���f��(v�M�a�R+�gsy��~�N����b�r���.��W�J[PD�K�~���su���q;5>Ȣh��l'~
���_Ȯ���Ŧ�DRaG�+�4<~�$��Z�V��T���
�"A��.?.��fB�~J^
�����]��w���I/X�h``����2�R*�\�_H�̔�9���M��10b�.�[ΈƖ|�*�d�PB+��(j��$.�#h�B$G���zq5Uc�0nst'���v�H'{��c�S�Ma5Qi�r�>07�S�z޳a���P�L����rt��wIX���eIC�k/�����7�:Z�3��Y�m�
q����\�G�I�Dw��^c�Ae�&�>b�ԲƺZ�����j0Xm��������5Oà��#�Ǎ쫜`kw�����"�m�c�G�k�팝� Ɇ��7n��`�v�3c/��0���د=�[�'�_}Z���o�`䓛z���1^�&B�}�W}������J;�N��\6ܛ78г h%��I��y��Z�f�ō�y����-X��~������ߦ��x���8@�¦�"�.�����=5k�"q��Ɋ�si���eXT\,�Rͽas/�/���O��|� �L�� �h�jO!c7��������m=imN$/��1bՄTJZE�.�r�@m�TR�H���U�����n}BpDR+ �E�ؖ����
����8s��%��j���^T����eR�����YSbч���^v\�ZAX���,)��3�)�M�a[|4���2�7�ۘ���L%���N�3��D��_�����,�lґ�� v3.,�lR��p�]s��O�eU� V܄ئ):��|�*�rO�I�+[���U��f��h��y/��|=@l���Fn��<Cm�'})���ڗB%'�C�@�TND��xxc��$��2����T��A�$��`)ُ�i0#�D ����g�󪤘җ��&�"ێ�7�U���zPDS/N��0Hz?��F���S�3,�ѠK̀#��%0���T�J}|�5��z�
,�:\���Yo���|���l&ni=謳،�8`����p���(v��
�EƔ�^��z8A�h�Z�-��$���<o��c�!�hk.1�����J����U�O�.&�i
�����(朸d={����K�k@��y�by��H�_F+_7%3Ro��-;AK&��ka7�a�To9?s��I�8���Ƕf�F���%1W��P\2	��+�5�!>��c2�=�#I�Gc'~�XQ��i��'�_q�X���noTz�`'`�
z�*�ߐƊ,I�w
n���ů"|<p�:������v��pR�, 6%^4���D������!U�9�YPYѾ=��aNj�\(Yr$���>d� ��������xNެL#�*N�ގ�DV�*�{�;r�
�����Z��(wv�=Uͭs��9	^R/�VE28��n�ލa%��J�|`+��!-�eA&�#�A$V�)�p��9���0+�G��id`���CN�f�*֚9��	YG�)	�a������=|GE�� n�*������?!���WD�B�PK��)A|��*�翾
쌕��4{swD1K~EM;����ڳT�k#ǞK����eN��5ʕ ��]Yk��i���zί��u"x{��vĞFM�,�g	O�~�����H�	��_dY �x�oC4ygZv�,��W���(��g4}�X���	�I�v�.\��V�g���S� �+���Sf�$��>�(6�qt���n\9$]�PK�g�m�ҥ۱0� ã�*tu��;i�����5�����6��p-jf!���n������GyM����
����^Y"q�oWU�U�￮��v'��+�V���
��1O{y��'���e���A��.�kdRf0�H�G�t��3�ݸw	�t1����[�G?Y-%(F�.[��.2Q`/Xw�gn�b)�}�&	��dr�FF6:e䎻�r+h�O(�vUWO��n,'u�N�;rh\�J@W1�1�3�*��a�9WM���z�g�������B�Z\�����2R��.:�K�˼�D��C�L7p��lު��<���B�ֿ?�vbT�<gAq@ȯ=��Ƿ3i��-�!�;[^Yں����AZ�N�yM�A��0�Z̧n7��jrQ�� �7f�0��o̐�ф'w]�+5� �QQ�R6�"���V%�N�n�(a�2Œ��é<���t퉏/ETf-=�0�4�_n6(T�}*a�ƎʖiK9�2]�1G����y�ղJ}uqH�`����V
��ﶛ��ܶ �m��Q���*��b������`���,	�3Ӗġ���a Y���b\���� �s�pd��wɛ.����Hy��F��]�-l�C�$	����0�b|�6� M!�׌�Xl���{�Y��0V<Z?1��y���E�A�A�H�1�'�S��~7��� 
���"���s�o��W��ھ�^7�x��.��d�������+k_�t`�{�ʕy�a����J��\w.��_�����h�B� �҆ڪ�nv�����;}�� ��#�-�+n�klP����q
CR컏�` ���sC�sf�r\�{������e x8h�KIFWF�2y޾/#;݅y�ּ��u�74JF�8;�c�t�*]����j�<��y�F�9z���:B<Ȇ�{s�0��>�IVQT�4�z�=ޔ2�m%7ݴ5�O��(�	��v3���l��KT~��4A�-���W m��?�����e�
T솪�9��b�v�nb�Î��!�z�߆	J����%E�J:ۚ�Z2�(�����SUm,��+Fx�)~�����P��bY	w�e��d7\SA�f���[Q���PX�B���\d�9���X����Q���*�M[�ӆ�
&ֺs[a W��j�8֮������A�	��\�!OD�\] m�L�P�\�=�;�˱�K��S.)�MS��c�z@��*�p��菕TX*^�~y@���A�����Лujy{��ٙ�}�90�7�`���b?0����³�~!�BY-98AV�7V��^٠%��!)�&�]�v_�tn\������R�(0���=�������)u�\���xo�;�=�b��B�O� ^/�%3�%���EO��Tc7�`G0: ��酠ۆ�q���d�OnwF�u�<�U��-��p8Ǭ�=��@PJ�7�Ql5{x6|0�0��w'�����w��,��z�`��2��F��^��_C�>	J߭��`�>��Z��9����7�/x�а�_��-���/��s��mp5��6.(�� ��k� W"����q����^Fa�EgA����d<qbgh���d}�Lrm���Ee�2��Y&;]�[!��A����M�&5��5)�����<�RP0���4�FC'{x�+C�>�'�1���f�6
{�@}Γ���^N(�� �±��zto������D�M̹�����/`��7������~tAr���Lڒ�4��K���LUi" *���[���%/����}�a�2��ьt�P��W!8��x%e�dC� 	�y lO���rȡ���QZE�7bWa���6)~�6W����h޵��_�d*�x%K�\Ҷ��#�}�����:~���&K�Ex&2��)˛D���4��X���͡-���|�Y�>��4��5v����V�H���A����^0��KS��_���e ��'m�옆��+*�ZK1�Bơ1# f���b�
R�mEz�Ŷ	7*	�u�4��ENuhd�����/X�Y"�)U|	W��S�M>��(��2'Zyj�� ����T�>�N�A~d��!m�B���;!�_����kmF��
m��;�ō���2*�>�I06]x�[#�*�WlS���	�#&}Y���JIq�9"�ҡ�	VE̓TmSƹx�E[�q�"Z<#ph���ه�?��L�_��	�����I�W�2��ē��C�p�Jzk>U��Xdi��Z�������Ls��1	a�"Q�84u�nѱ8�N�Ss� 6zV�ㆥ�F��o�nrSF�I�P�I��M_;��Ȋ��$�u<i�6�����Qh;,�դ9��l͛8E�t��R��Fet.r�\��4�6{�'�~�];�����-A�l�ˇ\��>�@��v��HH����MۓPK��%��2V��'�=���Χ�) fR̂�P?�ݗ#A�U@�v[h�G�D�<�}�a�l?V�Ӎ��^V�%�t�����ϤW�^���۬�KT���p��m��HBBT^5�6�@���8�l/���l���wI����k[�<��2E�э� ��N�b�kk˹ߋS���'&ߌq�Ğ�۩������U�f���ź��"��TU�(�}���_��x$&Z�T�6��}&C�}�=^�Y�P֑�l��p��(���73�g�~2���b�$!�PE<ˢ�BR�w�3���A���M��@�h�}��R�'a�@NZ��H��q�c�<��C`k�[�Ѳ{P��W#v�̲}w�f�yXuH��p��/�<���vvj��M	<��T�נ�eJ0�� �B���D~"�K�@�*��G�Xn6�z���yT�
�u^����,0H�8!��z��T��!8/\L<�\v��h�;�;�$��=f�[���˽�C<m��,f#ES�_��/ˠ���jƜ:�<̐���.1��7���t��Q�M/�|R!�W���.Vcq�G[������l��W�I?%���I����$��y>�[? 5X:���t^��	R��s��d岨I��?���V=��vr�	�͵N�����@"@��]{�	؋w9�m|�2R�J6�ٌ��Jq�#n�@F��*?��!�U�_�7p�o(bVI6ֈ߻���i�Tڐ<}��V�Mi`n0Z�i��p���^��I�$ܲ�7^{{.�q���!r�B~<��AUH5���7��Ʈ�J��1��oem�q'���
_����Ҭ���+���X�Z�Q:�yso8Ő|����K��Ks���?߫5�h4rk�Ec� �����S^������׿�����9��{ZYޝ��nb����1@<�������f�T����%�!�nRh�Ջ���I�^��,\	�9�L��q+n���؍Z���O��'�yȜ�X�t���!@�'~��^bLf��^�w_k6�D�J�i(VtV�Ҷ�x������p#��r��<�![Jt+0)_�������^ݫG��7�]f��81Ĝ+�I���A�� v���ML}�%��`�'�|��ɞ��<V��Ğ���\�wJlI��ȼ�3t��V��@��\�]�"�M�h	e�_�c�E����@���E�x,��;;�SkV8�F0�X|���1�q�O��em7����	c�;�d�P��;�+�D<���i"��J����:�P�Ki�\�7m�d���M6�/;�ͦ2��
�� v�K}+��_�t�B�q�6�2�W�p%�� �>�!��c��7*:�rb;��~��v� l��8��U��.x�o�x�y�'�VI���+��HU"�*��q}�Eň9L��{���[c��|v�W��K�o�!@XZ���3\2^���%6�~�b�.a�:��F�`�œ��)_�9���E�i!^'� ���6�xL��y<YV
@h�@��"a�}�l��E t��J�/���l��'ي�?��E�i���-������9����U�Y_�#���޲�{�["�/�촚k��l�4�+ϊ��t �e�� �_z���:��#b�	�� ̂�g�#Y���Idb��3��a����}/*�9"��0�S
Y�F#�e�>�Il~�d��CF��K"G3����)X5��G	��S�R�\\	>�c���^���p%U�'"�橛`��A�ҟX�a,��M���Z$���C�F��|i��c��doｶ��zQb���|�p�Dk/0��s���0����^DHp��4�ܛ.�ݞ�̒i��Ɩ#q�R�Oe�u���t	�\�IX걨.�&y���>�SȚ�����\�ј-��Nt�7_�A���W�nN7�:�h>Q���䯅�y+͇_)ߏ�-I�m�|�������S��u�uKRvw/T��x@���U�Z9�O=WZ�z���7O�Ntƣ��t�d]�v� �b�l�*K7�R��.�c<stiԁ��!�M3����N.��M�V��qU�ML��-!e��-E%@����� �y�֭�!�C�+��/�lf��FA�Y�P�UM��5�M5g�{|�����jb^��T�1��%�j���A7�O��b��8���y'*J���9�?h��T�*V�¥��@��&8츼g����Q��X������(�4���H��E�.݈�V��jnt¦VLa�}��u{�Q���1�Rs�`߽Y��xӶ�&�bU�M��#AmF���b �ct] �?q�d�1���U�tv����b)	�@�=�e[$_ U�����J�E��PS5ٙ����0pfE>-Ԫ���aҞ��%sk@�"$EQ[ߍZ_�J6�.˿�5�W�7P�:�4���'o�qf���&5(�Ӂ�:Fx�Q�d)��3��ML�F����G����O �T$E�q�oj�T�j7{���0Id��+]��s�j_ �=�I�N�]K��Xh�Ԛ���<^=	' �}�7�$�+\_�L�e���N9��uh���^���y$���F��YUe��pślC��r�a�TTf�n��T�N&8�A�/OÆT F&e�(!����>��p`��(����I����F����k�0��zh�eQ����1������.T���{���$k|	�?�sh |VSSz�uH�g�Kq����Srxnl�/�~�ܤɃ �r�D?5!߭�a\��,쥀D���nm�A*�_S�(�(U7�6��(P�Z��(�T�����a6��D����!��/<נE�=��1B�������"o��Sbb�+1ͱ����ϰ���i��j��#W>��Y���J�v�x[�1l�L��B��{�'��2[vC������*�=��/�V�!�/��XL����!��5�����o?� ����&#yU�����@�4f+:��r�Z	�m���6F�w��C>,�yiLp�>qc����c�]~A����W/�g�݆R��b�5$����<����F>򵉪�"B�Az���t,��X5�S�ކ�����h�1Pk@���[0|ǔ�GVZ��	l;��'k���
���=c�n$:�Λ]���YH��-q�a��$��k����;�P��u$�|��/�,h<�"������Q���nA���+[�Lf��3(=�N���X���Qk��"7� ��6�Wxb�����ְ\���p����;���W%��"R&��eU��y>��
�C�����+�x�����p�gQ7D����g��N7�!Γݽ��^����� 6�0���g����4�f���S}���H��δ	z!n�ܑ��c��exU��Īj�Ȇ�X���/�y�=*l��#��н�f!�SY��v�u���$s�
fZX�2c�˥ʹ^�����5,d�q��3�����x�K�p����ǐ
Li�;d�e��Ĉ4��HG=��ƣ��غo!c��;
?r��vD+��:�ht���5����)��5�����MI���w�@�ژ���^��'3k�`b��z�[��R��,ƒj�K��89�������3m;�,�b�5��	�ٱ��a[wG�1�6'��w����T���	��{j��q '���]c��<��_I;���T���`�2џ��vr  �uI�C?�kX�ʢ�s��R\���^Qlo�z�_�:�h�Ƃ�t�K`b��ҿ	+UM��;�%���)����-���u�\���>[~���ZL��Itu4U�����G8m��AT�rL��:�ɭ�o,��_P2 �LYq��C��;~*��C �ً>�<5̋�\H�*S(�/�\@W��/L��T�n�u�d��A{m����g��k!����y�o*��&ޅJN'�j���x�l~�"�a �^ሹ^/v̪���ƀb�H�z���Y�%x���z�fYʞb�Z�g��3�<.2�5�6�`2���W�O�kE�1�P(͔�r�I<mֽ����e�_y��We��c8��V��	H���`[����&Iו<Wx~M�i"d��p���R)NRq��N5m�x���8�JN�v(��I�� ƞ:�R�I���8��+�4�������:��������w��A��
�#_~�5zR�#�d{�����ooX���ݰ��|��^b�
�����:i�@��^�7Xr��*���!{��s�i�SBt�ρ���뿳K7s`I��p�D.���b�Y �xh�;��[[��	�[�x��]U��ME��]�5=.�vJv��
b����HV?�~v�9=��@���Kz��ͨ�.�5S���PH�+yL+i\��B?#IN%���ip��ݩ��r����E�V�f�B-�wu�:��]���n��t�묔��C^kK&�����/c@b8�#ǙOa����\�E�-����g�����۪���6�(D^�@�^�ȊPS�j�]�㞢��MI\`�� Nf��A�4�j'�ۚ�)��??+���C�: l��^��qz�oz��q��4��Zڰ��.�F-}d?/����c����27��������;$�[��r��h'�>������yϗfl3ur��L����9��hCf�q^�G1�������ӱܗ�����M�1�4����'�:�.�N�a�ESt���wLaD�,�����E�^8z�V��S:���=�+j6�P�{O}P�ONa��[G5�5�W|��3s��m�΍[���!��gJ`G���A6W91�'�W��e�7yE�pj9�!ĉ�wGi���u���E�ر���T�t>�����/�^�>�#L��`��Be�y�M�3{�����`n�{7�&��w
���Wrٰ۠�[��A]��Ǜ��2�S��uC,�o=E��L�|�
�oQ*R����Z)���c^Y-�����:�r��/����:��ZW�y5�Bx5pk�j�'I��_��ٱ%jK�jL�CP^����7��Χ��|����o�~L����zN'+7�/�܂��Xg��Њ��JRL�S.�����i.���Y=�44������9vD���Z������c��fő�v(��G@7��:���zT>Y���Kgƀr�K��[t���	�~�.�x� �3�{QUY|�V(z���K��= #F�Щ��������m2[.W�o�)��j���cS;|6[8��_�s�T��Y�%��|BJ�e ��>|�.��b
"����F����ּ�����L�yuO�p���o�0�rs�FT`pP��q���,�3�hfٱƚ��q;Z˝$���uz��툳�fq�|�σr���q��f�Y���1E6!�mė��J6�ӽ2�����63)�:�:���������3u�a?��_|�҂S���?�-ț��a�B� ����s�]�rF/]�#\f���6^
�'g(�?��N)R�-��̶c,��5��a1%�����C���٥9w��Ⱦ�K@Z�X5h܀)�;��2�u��Go�{���j�1�:��k87 )ԏE��N��_sc
�#p�-֙R#�d��ޝL�ɯ-����{���>��.�{g��-X;L5��0;�UϨ�O��Ksn�A���P)��6��^��i$;��`v�B�-�ކ�GL��4$l�f�y4#f�qNU���X�c��T}<�)��57�>�oVç��n�X'U�j)�^�f��/,���7a��BPdLN,��QD�=�_HL}���S{��9��3b��
��g>= ��^��@�p)B��Ϭ:6i������� "����D<_
m#Īe�0��	sq(#�����~aP����8��5�}����{�y�1k��I�3S@ VZ�=ۦ����s8'���݅C�'������7�eu'J�D6�5�oؐ��@��*���b��щ��f�蜫-��5�>B��]�_�w��x}�5�Ӟ����A�����U�5�/O�ڔ<��T
�U�]�2d�Tt3	�C�dϕ���J��S�v�=E;H���ц�AZzl܊����������L$�K�U�Ü9�u���:�ܷ��F��toKմ6������"��T�ۇ΍Y�i�n���hB
:J(T��\�+K]���C7�1>���f�b(���$U�EO��/.�xQ.��䲼��(��*+�a�b�~}y�7�|8(�&�I_ߞ�{'q�W^
��b`z��O�~ w+Qţ4�g5���%����"��Q)	��ȷx�..�NE�cjh<��������U:��r[�ySG��I|ͫϓ#� �@�έ�72�2A��J�]�8�{AV!���J0J٩=F��לa�V�܅ыJ�iU��X+^�!W|�u�l�<4؅�Ϯ#g�d����D�Z��P�\Nd:�+k��%�/��0�_z��`$��GR#�q�44jt���Q��_���O����
�(Q�Tj�����j�ց'�*-���cao�O<���#��2��Z%s"w���,tS�Z�2)���$�g5@*&3·=�+���S\���F���3�o��N���E4}�j$s����b�N[,�f��A*��Ӏ�xX�-acg����������!+���r�fE7��U@����o���X�8�,��b��ij�2΍U�������I
y���*i�,��x��%jN�*i��059�橲�T8dY��P�E�4P�: Kگ�_N�����q�
hj��
Y: Vcw�l�dj�u� `�R�4,��ۆJ:���J��S�:c�\/ѡ��i��Q �@8��bYZ�B��q��6I.�,ْp(�'"\��d	��v�dE�-Zٍ.r�@�i����ǣe�5�� �����2rp�Q��å��.(T�i/3�db���Wz��Q� ���uՔ���e ߉;�Wq�[�m�I��^������p��fP���n�����}�J�;����"����;���^Fs���FB�A��J�ȩ#���)rOݤ����u>fN������y웬�AȅI��P�"*�F��k��~q=D�N�8�|�l���J�`�@=[2���������!P�̈́n��Wme�j��7���[�L�o�����my���g�@�f��Z���+���+xb�?�&���q�S}4;}� b�M�Nb�_kƣٶ��
�mi�d+N~�]")��:FD�X����jKd�`��\*տ�[�0�12O�:�3����me���3��Sk�@fY-�/7A�=���gho�b�w�{��Ia'Y.o��	�𷏸�4G\�7��z&�S7�Е���Ԕl3�6�{
�'�Yu��Lžʮ�+矍�c`prRq�[g4��w�U����?5�d�����{� ��G�9^��e)�m��i5��'��e�~�n� X`č�t��<�g�)c>3\G���jwe�:��W_�;Y=�F��<~�tㆎI $�w�l�PVɼ�Z"��ݹ����>�����F ��=h� ��9MZP�㹚c=Q����5<�]�Ǣ��Gd��Yl�
#4||+�ͼ���oq�?��6���)�S~�f�P�Ck��D�Lw'W�k�`���!�"�g����fD)5���䔂#�s��ZO���1�n���:J7f��]"Օ�A6#�3O�м{�(A��Өʺ���u;��S�ƶ9�o�O�#Fg(哧��7�e!6�|	�� Z����q/��T���/)F��i��/�hnO���CR��&�V$Q��҈��g

T�C�@���I~G��,/l�|���7|�a���嗼@OdĳOh��nQq��k�<�f�K�HY@鱃g�G��;��ُz�
}j�4+%<M���[��U!a�G���A�s��ӟ~ɜ� �n��e:l��n�)��˙���" }�Twi�练�r� �� ;|^��n��#�z��zI�M���A%��]�l�@�s��&�$�ƈѧr��mY�4�ƹ���v���	��Ꝕ]�_{W��I&��o����A�Y_(g�7Q-�8�=�y6\�;z2�z������,"��i~!�$F7']Q᫙C��;o�{�=���>��ABA�X���\�%���z�r?�����Y���c��#�|�+9Ŧ3����\E��U�*��}�ː�6i��:S \�`��;R0��t��;z���üx���wT����c��J�0�_Qu��!�3A�J������|j�'��v�?DL���K>��,9��C�}�y�؎g㒖Tޜ�Z�������%��dO I~�N�=U�ud�lFH�P_:��D�O����)��!�rø�Μ��{�~�J�z��o�
8���z���/����ȅUH�-����'�x�e���T��c!������K �:b)m��+��ߪ��t᪴�'�/NH�4QVv���y��)���ՠ��I�R���z�^���'�AZ���}��{�i{�	.g�����_r�n��$LxWJ��߱�H��o�Je2���]�����G���_w_+��Ewh�r'9pp�4.,�7
&G+c�r@b=�P{yb�_�Ez>C�qS_��s"��0��w�h����<8�%��%�;QL�G��O}/�����0d�.e�*��&������ә��X�ÙH:����]���P��k�F;�2mL=�=��NM6\%�5���h����$K`���o�ę�a	�Γ)��E����d(nc.��	k��?���M�S���YR������0�-���WF�K.��s���'�~3h2�9?<:�〳��%	�A$5�@�WR�p֭�WP���+>%�[¥��PKN'\D��f��*�Y��:��f��ե���fzNK�����<A�)4���]z���= ��Ћ3g"��]3&1;F�V���i�Xd�h���D�J���M�!��.�(���z�U�1T7!*D����t�W	v�p]�ȵ���+�G�)�jC\�����)>A=���� �uS��4Z�.��V���~x�f۷�V��{{��ӹ.�7�+s�(@D�{.5H~�ٍ�ܙ�Ut����;H�)��l࿩�:�֨��d3|����6�x����y�9y�;A.�n3:S���Oc���l{�[
,쯪��bꉜ&��v�;��&w�d���ơ����ac�
DlA�-jlπ�\U�h�=C!��~f�*�wR(i=��-y:�1q	o�:t�m�l��Gs+�(Iɸi</�Y��t��,����B���4�$���=�&L�����<�X��-�q��]4����Ɖ�Z��)����X5ؾ�&�"@(e!OB�$�KZ"�J��:l��G3��E���ŭDb�LN��V'�0"A�����:!��IG��VL�2��8��a1���{o!�L,X�z�wؒN�)��Y�2طi�
[K���~����.6�B�.j�/�� �Ų�	�J��+%h�ք��s��d�Kf����� u?�p�3��4����B�5b��3\Td�
�"sHuѹ҆5���̫���\N����n핵�C�"K��\���
�"_��y����kW�Y)���m�X���3G&z��ėC@̽�⎸�Kn�r�p]`��:�&Kpo�Kp�H(�D3	_� :o��K� �i��QC0�����3F�%I?]���O�]E?U�w��@L��
�M��xk�-�(���?#ݡ��#��4��KP�#�O�����k�^E��#��Yt^oZ(ҝg�NW	1*��5��)F0*-�tQI^���x
?�m����-m7�i��m�I�2d�8T)6���`�(#g۳I�v��w��麧jG��&��2��O�/�ǂr_��!~Q�]3x˅5�"@��ڃ�~L�l� λ�W.��p��ʷP��	��61�E����-��Y���]6q��K3�t3�D
���x�C.�,��h1�t������qc�+��V$���Q=��^��,�����i�<LĮ��т�+���_�t��{�K��n�H7� ��4�0����i�.�?�oAB�a� v�X�I�nۺ�{��A�1xujg��c
tU3�6?Vׁ����g�%��#�&|Ux('��#v]qaTs���Yx /ȏD����rFg��s7���C1���(�ݑ���S�/�7Ϙ��v$�o<?ru66�P�����U�}c��r��&i�b�����1 ?	�_�f\y�5e�a�rE).����GZ�e&���hK�1��YJ�\`�gD���z�D(^P�{�����B�t���%�0D���kr�W>_J�}�co�
̗�	׈(�)L��?��I�0fgi�A�꺯0̚���='��qV�Q~�k�z�!QƲfR�) %��7�3�^�)#��$O1�O�x?���..�I\95�1�VG�$M饳Sd%�Ƚ�&�̅�ƕ*���>c@=-����zz������g�r$djAg�#gd&a����nÅ�����=�:r�v2.�����΢����88W�5V������q!p���E����l�j�JҐ�qz��L�����L����등�� �B�9����o�`NQ!̳��
�N�>���fQ_�θˢ���z���_�AT1e�� �H��|�}��NH^ɣ�!����j�J��i&ؐ���|�-�;
v˭Ҁ7 ӝ�?wH�M�1}�Z�\�o����h�U�s���]��xŨ�⩼䐽k,Gr���ݽ�0�nT)=L��y<�M�= ��DFd�)O}��T�����X�5�67^1��1BA;�&�o��ǓⓖW. �zG��+����r7�G�H�>�8��v�dTlqV����\�dw�)C�q��� S�%Cq��f*����
�3���sѲ�*�3e���Ut�{���рJ��m��q�S���h�j�s#�,iG���Xb� K|�n0�ꊶtj/�N��Y����T@P��CQ]���$^���86��.త�f�d,|��n�NJv���?b�³�����G��l	��p7�Ɋ՘�~�v�]�"T�g5esʪMr��y絥+Q��8tc?�͘V"���i�M��O ���;	.tbuW��y)&{�� ��v�B�ߟ�b�L&�-�F�7>�� FQ^�����a���� ��]�щ=���-Φ=:�z���6[�qHBP�
�
B�X#���ԕ~�iZ�1� �:{t�v��z�U����h<_��"��ȷ�f�֑	ձt���_Q�K��͞8H	�Q誂�	<�5��F�0Z�r'	�(��8�J��/5�k�9����d���󵘼���U5��y^N��	-j"������:O7 _v�:bRG��v�*����;����j�έ��u����jۋEV*�B���iED��G��D	mrW~0E_�Ah[ �[���"�l�#�!�>���)b������sz������,1oH^Կ��&C�R����I=��dsj�\�]߭��KɒuԏZ{d�ӭ�T]`Y�	����PK��z�C������z38�+��e��"(	7�e������	qhw4sN+�I)�$�
��D�kg$�4����O�i!��:�|vK|��>��y"�r VP���F������Q�R�"��E"n;�dz�j�B�J[�T��ti���X����p5���a�5�hFH[�ܟ�NB]�����e��nUC;���qY�=���ظ��������c ��e�-�Ĵe���_�+i=�>�Uȑ�$B�ϫ�� 4��� +h�m_�RO�Ŭ��,��
�ɞV�^��&~���&G*T���$+�;G@�oOHP�����le�v�Iv����
�.\̿�C��FTЕ�[|;O�p����Jb���l�@d�����Z$BR4�^U9�rc��0��5��$��Է��lX���Xh�C!���i�\H[��+�e�b�h4�W�b>�ŵCK���E�CC�j���׾��xԦ��Li�tb�1n�h�6r;d��cжTˮ�o��3fck]8�^]+����<�1���e�˴�B��� ��^�D7�x|.���©L�z������j�>y��3�!��<������
5�����ӑ�A�����3D>ڹ�FZ��w��/3GV�@+lX;�S@�;��9L���H6!
�ϖ���LRkcIiH��
�а�n��ATr0Bٶ�{#7�ю0���y� +�5 Q�_�YYz�3
dt������s���	?�o
�u��Ș�8p��r1���
�fCЋ��xkb��Z���- ��+�����7�2�xA�Y|P�'���3����^�}Pt&�3
�hߒi���5-���+oIh��cwA'�q@��>��#{�A+lĨ*i]�}� $$T���U9m���kӏL]���v]`�1;�B<��[���߁RP:��,��, �4�r�7��}�����I�T+KP�~��	�!6{�L�`���0�����h2h�uy��I�NTz0"@�����}b��*�菤�}e���`�]n?T;��Mk�ߛ��]�����:8AW��,gs�S�K���D�U�7�ϰ��<�Fyr�zL�ɋ�<:�̖1o�/�x�6�B^���=zB�d=�__���S�$}m+�c��x탬���|no���BOa��]�����G�?pf?��Hhqޑ���]׮E�﷡��R_K��n@Ku���Y��:_é��H����;b�,r0S]�'�b���S�b|��"��&��3G���&�0�Ҫ5���T�4d%�k�=cN��(��]H1� ֕��m��e	wz*`bN����}�U�u;�=+�����G��������E����5��Ge|�9�5~��xd�5h@VhV�	�13ʱ�sy�J�8�d:�X����;zLJŽ��2G�o��6
e��=�lY0mߛǪ©(Z\$u�B��6n c�H-CY���-( �Ո��Anf觋-U3�O�W:PW{}䢌��t��O�޳s�dE[U�GB�+��ؒ5&��p,6�߾��\��{��%?Y--$ܡ|�D���r�%�"��o�0I3(��+~�a����Ć����g���7�rGȱ�wPV�˟
����
��3p��	�W)��j��Oz�$��=t�@w8��
��`t`UC�zc�ɢ�=8�	x�@:����dt����*2en��l��h�,�2W�qmJ�*+�g9�,����YT��/��`���mŇ��L:��H`�n��K)R�w~����w�d�^��ߩ�"#}��ේ��/��3�o�Gu5�ݾ�f��t82�/�����z
�n�s)z���9�(SsH8A��U����F�� 2*��KW�r��X�n�B�۪<_�e��x�`���z��&i,T|�F�a�[�����?5f*,1�6��?�������fo��Uc�H#��(��=��%㗨"�y��8i�L�z>�D�
t�u敨��R�	{-�m`F�!�W5&���=�LSk��;�;�iU���0Q_�cx~��n�$d_&��6�"R�̔��LuM$*�O4����P�$�Jj����1� *oxo#�k&�Jz�����L�yY,��-��ޖ�@�!�]��e(5����^cp6s.�'�C�oøӍr��퐃L&l�m���<��~��9��?�7:ٌ G�}��MեI&��W�%�Ђ	-�gEw�?-�O����Uf�PA�U@�Th�V�/8"�Ol���<�?�PF�V	�CU��>�ǴEoE��6��'��o�݃�x���Q�P�ъ}�s���{��`]���h��0w��s�����58��􏼲MD�����E%4C]���z����8#����X������� n�A�)7�ht��m���0�NJ��B}$��=G�ձ�Ų��`|�������M,������:u5L��a���g�S�KHQf�p�J6��a���ʔ�A�v�2�2q��>u	8,��A�0��M�"#�wy�5��Ĕ��kx�q�S���hƝ̠�"�e�x	RM��+��g��5Ȅ�i�3�P��c��a�r@� ��IB�#����, ��K���37� d�+i[e
�\�B��7i;n�q��Gva(��o�t��d�m�E����5�����$i��8c ������s�'���V�?��a��/�r�Lʌ�v���f��1���.+b���'��s�n�:4c��{LK�I;�Eu}�������6	"�[w*g4�Ƹ�/]�S����$M��W��b8�ê�@=�@ʝX'˫�B�1�Y�,���h;��YbK�8���M\]c� ����wy. ��69?��j����y.TVy���Y��_/5h��+��9�R�/��H];���4� �H򀥗VkTJ�|��;?�J��@�~�ݫ���&���5T��`�>���<�H�`��R�sg���6e9A��A����K��h�f�y�)s���q9�s�Q���O�D_|l^C���1# �ôXG|�j���W�EG��v3]᷒~b�!�:RW?,��헌�E�����ښ�Hn�Rpt�9l�<G�^�10	��8�K�xe���u��l����?���!9˽����K�\�#��M���Q�4����?�U�&�ݰ 0�9:���X8*�]~�Z��;��[ce��N�����g�c���I�9Xi#�=��%�[��>���XG���4s\c�(Σ�(z���!���`c�����gv\+T�q�Ɣ�����c�k
d�)�3�?�@�Gj�s�m����֩��WO�^��щ7�z��S�2sB@��sv��n�%k�n�u2��jQ59p�6:Sxe\��l�2�r�ᆒ�t��S���A*'���5�Z.��|���9��H���U�*��Ϛӓ0��	��e��:{\j�qc'GmŅ&��45�����Ab���]B�~�D�TV]؁hcꭍ�p���|��6���+QH4ZrV7��G�d���f�
��j��`	@C�:���%���鷨�z�/�9�M��_�o�`�nޣ�]~�4Fm1�����<��n�����_�ӣR{
�ތ�(f����yʪ��TS��f���Y_��oe�"a�VL�5$|�H$d��X��$Z���L=Q1|"��	��F�@/M����۞���ߜmo;'=/ӝ/��W$���kr8�I����<�g4LA�x!�V�=R/�C]�>��$�����un�����v:%���?h'�G����y��j������ݙ������陰�|�E��V�� Q������K8U�i��H��%Bܡ�e
�Hm0
^d?x5���c}\5�F1>�b<"���OE]¨���4�̈$,|>�@� ��e�*�f�;+��*�	�IP+�pu$;���������x��-��p��m�}Q�w�$ѵ^�E�q�X�M0j�i�q��fǚ���/�@Z~f'�r`�#�$���#�\j�iO��	����q뾏���猟�c��|c��3����U1��a2+>Qk��ި�:��N�-�5�p?d�ȯ�:e~�(��;��͹|eȱf�V��"�+'p��%�t&xC���]�U?�)u=�$���l����MT��
�5;m����N��Dd��`�}��a�KU������:�Œ��%��Eَ3��!6�ã�eu�e��gW;|K�8��^&�����k�a�coC����g��o�|������JD��{� wk�%�魳��w���g7�I�CQ�s���=Q�i�e�n�,u^0�31E��U2/Uq�$)��ٳ����S�5x^��r?RY;�l`�P�����G0>͊5/�,5ė�u�w��	���ONV粼L����8����m��7$��F�؂�=�i=�t{�3���?��qT��w������i��c�����*}D=7�j-�m�C�om��?�9�{d?��p�����v��� �r�c94����Yd�����\@��?O���-?�={z��NvA=%��A�ޣ���9Y����jꍥ���0t�؅#��z���_���t��������6���QL��f�x�1�ҩ2r���Vj=���� �������G�Z,v�X��Z�P�1�phʹd�LG��s	��"�:pCj'�=ޝ@�A�BX"��ߕѷD�#&\�&�g;Ç7��.���F,�N3�� {{Ͻ�h ��J:�3]���p��������w�>��#���բ��=����u.:��v�,�oD4�	=��1�`������z��g5�E����Zm��"o�q��B��_>�Y�ǩ��OuOr������^�~�l��Si4��NϾ�'���H��,�Q*ز����x���Z=�Wl!�K0�S]�]°��;�BXf��h/���Wֳ�FSr�W3�+�����fH��r簙ĝ'Ě!�<��V7���3#��#�(�7m�\@���Ϥ7���P�,����mh�5ʰ��(K�a����.�2]�4
oHN��(�d�~(q߆a�VRT�v�\8�X���ˡȹN�4��ix.���B�w��u�E�ȿۂ�:[8����h�B�S)�6�3�5�1^Q�s��of��HT�%�T����.-��nWp��n������<m��od�L�H�����fKŉtH��t�)�ծ���E�ٞ��)綌����퐦
|�o1�;~���t*h@��x?�o�5`!�.�R^�4�Ǚ��dZ��e<�n���?\2�A��o�]��\��*@u�sZ[������Ձ7��tO�8��#�+3IC�v�r?�1wN�/"���6��O ��#=J l:߮��9.�C�H�,��bC�z�:�DKv] 9��	m|�8_������+��lF���ަ;�qX��ZI~�j^�Dn�@5VU�+��L��M�{�~,j�i��*�ة�Q���;�)~�v�4�#k�y���^��S%T���7�K����n��~�S��bf��v�BlI����{�^<{����?���yYb*r�|,�Ϛ���|_��n���x�l�I�n�P�'-���'=�C�(�Ց��8�|V6�v�&{�O�iZ�\�Pyvvnd`�M���h��y�N�UL�Kʙ5V�����k�m
p��ܳ�'d��t1ͬ�JN��/h���T	'O������,^p���s�-�R��ͤ\��G�6���L�i1p�Q˥9}�yq34,�%�_��_�D�g�hLX��;?�4�<�AR�a� }�q=-��z�F�3I�9��\�yr��L�E ��ʍ�꾸ɻ�*ဝb#^.��w?*!b�'\���r��5A��Q�j��4��BH�Hf�Z�%�u���F�E�Z�x�i���B��o���z��w�1��v�����I�k�s���+�D=u�gɭKB�#�$��Y�y]#�%8E��'�`�C��sg:�h����`Wo?�m![1KS9��;�Rd������a���N�þ_����G����ly&ߡ��d����P�"�ґ��v��C�qI;�1F1���:�MK;yy��e������?Ǩ�6�0��R�G��v�"���q��e5�����@�Y�h��G� ~�h��ρ���o2D�gO��3�)�59����F ��&TR��M
6-TCܡ�cܜ��l㧽�I��ҫ��h�	�>#�qQ���0䍜UD��=����(�a�f�_�|���CԈ�|��!1����+yuú���^��C ��ؿ�5J&�-��T7���cJ|����M�nK���҈���!�zpV`�ksύ"	�äi����I1B3��Q<>Y�V�����M�dK_����(e�������L�+g���ʬ?SJ�K;��h�X�O��5K}!�������g���.�Oz�>��NQ�~B'2I�iK������ޗ��_{�n��k	�QV�t�BLR=�`[��3a���!�,g�����3�ҥ`h:�PHBG��� 6��Q���as���o�%�O�������f%�j����]�	3Ǥ+�W��'1:6�fg
�q����y����ܙ=����n|��7"!!4Ӎ�b��f��Ү�W�?W\*G!�.������[��an|U���aP��5�"�q°n;K�����1�b܊[|s;m�xw�
��m�q"���i{�M���^�P��"-�	�]���6������\�3,���8/ �����*���1��q���5����f��up���'��l�����L?R�=�m�9X�ă�`R�Ĩv��Rՙ�Sf�0��tz���A;�$#��dW��V�hV�F\E�m�� ���?b�(/?�(kg(E����q]:oK�)��|O�Z�E����=�j�.�T�����u}��4l��7do�d�����&û �e����p��	������"�͗����o���WB4�U�@��i�LJ:�Dd]_����'H%��7�Ҫ�u��ΊvY�����|8'�H�����>}��Ƕ-�4��\�D@�kcǋ�UWM0`6��|!�����'u4�������^(M%M�v=��k/��#�'"��o�YK��j�Pkc�Sa׀;�P��wWD[6%X�
]=�8=��B6��%͢�+�S?B��CZ��.�������|;!� �8|$B��Lc���T���>�c��;�b��M��XeX�O��l��ˤ��L?~h���1[�c��iX�~	5D�oX�v�3��� �u�W|�>����DH�l�܅���"�ِ� �7�`F��KQEM�9�ԫ��c�May���:�p�����Y&�x9U̵0=wu5��@��Ws��_5��J."೧��M��L19�un�K�x4��w��%��6@���������������b�ܗ8�1�8��7���]�gx�/�/������7_ mޚ�+~�������3T��A��Ap�#�i�*"@�����[�h�����k�B�[�8�XAR���s�A�;%W�L&/"�E8��C'���A��ϱ�!�r�	�#T��l8_�T� �����w7<\wZp�u��7�>�*[�5a�1�!�qv{�C�NR�D�\I�_�B�ᨽ�l�C��)(�p-�j��8C�v�菤Z:��m�����q0^���K�[�s6�$������+^��K�Mg&yh��_�9=Yj	C�n���Θ�i���NGZ�@ު\����Zġn)�p#��w�C��h �	|���r�a�gf�1��x����?����F�jUM��s�J��;s��n8�fS�+����; ֻ0"�iռ3G��D�%�^D��Yˠ�;�L2ރ,�ftR�4�a�pzt�E����oe�D�P�xs�Q�[V�C�z��g���ˇr�gul�P~TaP］�5mD�N;5,b�9#�)�|nP�#�7����(i��~����Ϊ�~�1q.���f��ʲ��&��x��PP����&1
5e�޻�����B._Uݟp���o��4�# Ӗ�s]N���Dt՟O�������N�n^a=�b��� z3�K�l��ՂB�?��uh�>ڻA�0N�`�3q�7�D�6`�'ZBJ �P�t��gn�}�ߔ�*�4��A�P��dH�!w=:p/d6��0J7_������ U�V

��K������Μ!Ū���u�Oy��)�Y'۞��}u�lJWod�\�vx.<˟B���ɞB<�z���7�zݬ��B6W�"�ͨ�>��*�A>�'�����5����Q�놴��V�ߊP�L<$e�����D���F-�!���|`��d�+��c��8��ԔW�efHlV�'���p�Y~��`�{Ivo���)�l�4|�希U�)���X�b��43s/��?��s�g��T&�����:#Ɔ��m�M��H���:ߝm+��B��'�į�������>N����Aiԝ��'�`%�i�ͻR�k�j�@��d"p�� >�m��n�U��r�̀�#� j�E<r�l������+0��. ��'���]���C�y�`�w�J�=�AL�z�p���!�m��@�f�-�L����C3Yܴx���5ɿ*�T@@l�(���I�h���qUG����U���ӬV
jӉ+�o�?K{{�Uq�	��cǹ9^�Q�2'ZX�W�]��൱dNG�*�{����k;w;>�T�r��Tai����vN�t���Ă��㋋wC�+
��w����ݵ�Ƨr~���,e����w�Dؿ����]�r_�Tl�n��C�R�iEzb��������,�/�/ʌ/��@ͱ�[�
�¹�7�i���*�d�LƆxDq'�������r3n��;���hn<�͡&�Ai|���U>Ҳ��,;��(C3��u@N��tC�:UJ ^��|����W+�]�l{q.¥j��'_rV�(������Cxjv~&��ƅ�Xzb� ?�L4�2E�<v�cATt���,y���o��=kJ?P�%�d\��������u%�M#'��7�̪N�h�T��$�j͑w�3@bOK�O58iuM
�L�`E����5�!��
R
�%�*[V���.B��=�yR��,U���K��h������&{Kq��$y��d�՘�@&��/��l�j��7eaz`s��??�x����z�������<�&|Q����}�,&��PΈ�3�IDڰ�,�_ن��ˣ#�Ey������,u�n�}d���2 ���]Ttܐ4�r���D�L������%��
�p���1�6F���qv���M�H�|՟΅���p�t)���vd�����p��.��"���Pf��9s�ћ/U��m�̛6 �m�͜8��Q�w�U��n�RVOۮ�V�	���P���% �ך��V�G�@��ԗ�)hɄ�5s�O�s���}�WnG�Z��z0�UR�諠��k�H}�Ys�R���7|H�9o�ZZ�9��6��vS%����������r������Q
6&b��;�x.$k�+��o�HR
�h���W[���ro�İ�X�G6�'��Cl 5ޮ?١"�T�x�d�b!���C�����#����2�#9&�R�G�,7y2x�Up��7:q������M��^O�=/��2�D��n������P0��_&���^`F����`S���s��U/c'E%����Pu_z#�ܓ�-�K}� ��	����):�gA�I�|��N�5)�wyQ��	M�d���I:h��)�IY�}o�Z�<�8��'1��Sf��(t&���W��]���5�&5�E����k.��7;	m�hi����w���xYR�w�<�O&+{x�կ������xc���V��6I&�kX�6Ma����Fܸ�0Ao�l���
q��˔�lF�cr
����.�0y�jg��ΑU�@��y��2�LQ2I�����
�z�]X}L�<��.YX�� �Ծ"�c6@�|�-����(�N��q0���.�5��R��C�4?O��O���&�h��S�C��؞p_��e_R-c��w���IE[j�m>4��ܑ�V�h�2��( &	|�Y�Lg6�l�v��g"n���!h��<��>�;����%�-	���x�b�0�0G��������������.�����q
�����-@�2���|����Ǣ�H����{�	�3$;�A9���t�(��M��j��A�X3���/)J���ϡ�|Z C�s�lO��奉�J�uj�z��9�д�][�W�����q�Bk�5��׊��Sԩ�����6��w���>̉���7N�Hti��p���H���tH���4<թ�` lCO��1�������*E�����8"�Ą:1(s����Bl,��Y�$��v�ǖ&Y ���D��KZ��҇���o�8�*�;�A&��m2Mh�Ǒ�(���o�E"Y�I�'��7�B+¸~����!	9U5�;o�*?���yn}=!��Jt�W+�_R�0�}�͕D" 2ˤp5�P�aC| ۿ�mM�d��Ly�:	��."���8Q�;�m֢q���m�GG2�0B�@"}�r�Gq�,��&�ņ�	ɜ�{�r�s�����^C��P;�Yi�-KR|kt��Ϙ^܇yQϴ�u���n��WT���v��P��z��}���h��2��'=�-���������/�'��Hr��0�	��W��
�B�Y�ti��R|��j�@>~��3�8�N�^�=���!�7b�R�^��zG E��q��4J�V���#c��vPWo�0.��Y��W9���`+Y�b��-��N!)����O�9��z#�{-�!��-����Q����[�6���k+��ϣP�=k�P�ʋ�$1�����#�#��"���z�[	�������\2�!����}�y�֏:$	t��|2�/��������
�Nu�3��s]:��>q�`�4��M��5�)5�z�ږ��"�!Z���YM�������]��pq#�v�Y�����뎟�?��q�T
�t�%nxʲ�� $�[�-��կ)��3�v��F.��4���� �cի���q��\Fi%a���7�����I$�yׄ������?1�h�V%�!h���n��6\c�7����cO5�r���,��>��낱��[C�MH�NI�l4P�&k�P�ĞT��itR��L$]��rS*��dk�1%�w��^ΰ�r�4��O)$����lB�x[+�� �kN�G��?4(�[v��ǔW��p�Pek-����ʈ��(��@��:^�g��89>�ӣE��'q��+B��ħ:�W��N�q��h�3�e�C�QR��t�N��-(�~`=���X�O���e�O���\Bl��U��L���ѕ��$Q���<��P��U'�������C�-�>�k� �� r]�Wxt�rL�Y�[9֌s�O!���@/1(��)::�����+A��	yU���·��>6�@���?��y�m�CNh7�#��=�|��ԏԖQ؉��Ī���4������D9��t�tn�&�_";�B�.�>���'�,��x�<�(�[·�t�,!���
�7����ٝ�ʋCx����9&H��A�H!Rw�`/��L�Bw�:0[���Jv@%D�n�I?U&�sB�Ƽ��Q� �G9|�V_?��~`$�Ȳ~T[���|0��u>�{�:iQ�NC����Ճbr$/M3G���_�,Fr�%�{�z�ћ�b����G�9
LEVH�����&;�y��Z�Fk���lؘ���X�� ����N�U�M�>����h��`���v2_�a��i�+��v-u�Ĵ�}�������E;�$w�P	&�g̙n���+���t0���,������^7|t���e����pꛐoM��h��9;��f'�0KvAҚN ��~.C���rh��C�pԮ�!Ls�q"L����G���_��209������aL��
�kW��e{�ԫAP�<��Z�>���Op��������W�]�<;�V>0��0vYXY� �������ެFl�Gı�n�I#�t�'Jp2�T�L��䇆T'�On.b�B�n�@|���M�xy>Zm�2�2�:$�4-�h`��֫Iվ2�jW��p�uh�;[��3?:��Odȡ,�4,�%��o�I��S��`��)�$q�2�*�4c%(N�Yߔ�R
P4��Tr�d7��Bf�����ruݰ+X��b"A`)��y�VF�އ2ؘ��S��!yu@���'S�;�B&6� ��0�+)R�
�8;�.6.cHK�.]p���Mr�X^�Q�V�%���]H��m\�\��~Ǧ� a����Ǆ�����JK�O���_����$��L��p������w�#p��dHs�!�66Y�f�.�ѿO�U��mɝ}�Dj�M�M����q�9����J��V0��z���&�	t�ru�`ZAi�n�б<�?�뎴�X����x��
n`&y�o��@2GN]��u-����g��r)���?${�2����7b^*Wf�&X��Qj�f�I�M&@��JY��ȇ��ߤK	�	�vX�ST����V�ɔQ���^��}`A��:��gz��l�'��m��u�\��!-�R���	���eX5��p�)�~o�=qQ�#��p�Q��д��;�T�l�̡�0F�[�]�'H[L����`�1cf�l�L翘���6!I��x�9�I]�^Wu�����e�С�)��
F!u�xP��+�����$�����FM���/>tE2p~4�)���L��ʝs����5F��B��hE��X�O 思J�ϕ��*J�e!����ڲ���f���܊wp@~`Ԍ��K71��-�m�|3���n���.L�t8Z�:�@�T-��y�����ۇ Rl����ѵ�ց���ݵ�_���_�~(*��~�� gк֘�8�7����4c: �����mT����x����3륹Ь�m�>yϦ�T
�$��5c�P�)I��~gK�����0ѩ�ΥK"��}Tܳՙxz��h%���i�e	�"ud	@���PG�l(3��r̷ T5�2�nFz�^Y ��^�z�=�n�����C��=_��=�6�Y����©2{l��
-o�d�:� �'��`��Ƌ��30L�;>�s���KQ�z����I������7��#(���3������\w6�9p�Ȉ}�5D)7����V�K�d)\	� 3�z���.�q�ݾ[��+ö��~G��#����\� r|ǲ�́>�A@p<�����p�jF����6H�P�����Uk�U��+��S�$�.�`U�F�u!��"�0����r�?���q���B� �sM{4[%z��G���|�y�nw%��V�{��i$�! 5KV���q�*V�D(��A�Ml�aTGj��lS7�Cw���a��.�>�u���7�t#i~u ǧclQ/,6/��[���I�&jFu��L�������xa�)�!�z*���0%����������`H 5>�l{�y�	��
Nݿo��zF�K���]�.q+��F%�hapr���չ�����"���R�9
6����/ǫpv$�g�C�\��Ǖz���3u��J3~/Vڔ�"c�)�����쾹��1:�'�zw����;2RY�;`L�)l�Q́�4�1�2��	�q��(����{b2�j�<t�����2|mm�+�v��œ-���b�"��/�ѓgp�D���b�"�yXw`�cW8���I��5��@�ϬU���|ʖ��h�-�r��eպ\��?��w�}C�,��ZJ/��Vv'`���D>;|��mǜ��w�<��m/��u�M�эn0[	���p|��1����GAlܓw_������R6�΄��&W�L	A���j5̞i���H�������\:	�7 �_S��4>ѝ�\�����sn
�s������NR:�����Fs�w�/��GtN���iA�5��"7`�ncC��X�@ 0�Y��j(> �O�	�.��߽�7��*V0S���0�m��+}�Pw�L{�2iQWkJ��8.���W�����Wv� �CY!��0qua�T�JgXI�<ѿq�¨6��eG�`)�QsN�VdZ���-#N�Nl�O���4��0;��/2���o�b}���=ݯ`�H��W*�~-c�GRy�|��M`d�S֛����c��>9ߑ�l�NT�a�����l��x
R�#�X~z��>gv���ǆ{>�P�"�tE��]�
><qL�k�8�4�h &�Tb��Y��9V���J�T�����I# �������lb��
)<��3�ޞj������}�@1b4k�>�:����)6A��ѦD����	�
>��r^h�-���u c�C�Ȯ�4��>�B��6b�x�]��XR+IW�C�����	�"|^�b~�uȵ�Rc���i��D�1���Dn���hlGgi�sJI	cZ�Ks?el��x��G��2äzeK�Tg�\�����xޯ[ЭY�M��J�����I��Ғi,%t�`�/yc���{5�94��u��~ۆl�a�+���5�~�x捲�SKG�C7���SZ%L4P7"!�ݒ]xڧ9P�:��(3ܣ|����U�Sh���G�B��};��>͚���?���SY�����>3�	ơ���	lz��IT��L�C���cA�9��4{���^���]�3x�]?`��=�f7!�Q�u�(�U��-;�:-�x8|�Ri8�9V�a���ε�H��D��:�B��R&��z ��������3&��b���	���tA�����M��S� }��"ha�6���F�N��"���)���4v�D���I�M���1��������N?���%^ͽ�}$Kߓ���%pL��ꐃs�� <)�M�����D��/��aH�T�5"
�0�(�I]���E[��ʶ�����q������z��`T�?��R�4��<ю6�e�d>\��;���i��[k���c,�+�T:u����7�W�j#A�`�<�I]7�ǟb�J3��^�B��꧴��[I�ct���l��v������$��c�@��kn647M\���Ȗ���nhv�ѧ��i(�.�2��&�tL��8߯'%6<��O��W�nrA��/e�f }*j��R��,�"n��Ѧ��9߰�IܓL�>Sc�J��_X@0��9���L�au��v�{��`b��ˮ�c���d� �q��H�N�� oS����
��j�f���2��^Ϭ�-�/=V~��J�xK�k�Ŝ%���ށn�"2�&�x���<d������q�	L��/E��H��d���iQ�h|f(���0�5���+�h��ll�ډ�
*mз-��c�O_b�m���f>¨F�\�� o�r�5�^���g`�v�w���(�,��(�L,Iy�O�Xqo5�<�X�����]t�x˷��SYɝ��M����3�W3��%^#$`���\���Z=I�5���ϼ�n����%s;��:��FA��}q��?/�	8	T��}�$���Fc$�\�B�|.��mc�iB��iPȧ�����V���&����J�������7*c��;���D��DN:y
!q�h*��r�-�o���zk�������f+~9��~�	�W~��e�\����;V�+,�ju�����3�	z�1[�Ǧ�BBׂn\{oa����y�X���+�����Ms��=�L���p��lw�XR�X'��
H�%��h,ei�')������&�i�\�S�s�p��@�?.kL�D�#��t�D����8��k�-�ئ9{��[˄>��Da�M��)�8�R�"�4mez���|#������X	6[�6����U�w�d�*bP���LD�t�0���uÕ:jV�Q?���pN,Շ���������]y���4�ȿD�MJ�y;-��^Xc_�ᷜ�TK5ڀؙ��!=P�<�m����s���l��}��Hw�`OI\^� �/�m�(�RA,+8n�L����;�A�#y1��Ɓ��H
&u��[����^�������v<�	�"�9�����`~��>'�C	�	V�=[�3<|����<�="H	��Wһu_�|�6�Z9A�3��~�����T4�?x���W�[P�X�E�:�\q�A����c!-�n.#7��j��μ�T�M�Yt��+�P�~�f�-E�=G[�\��pA#t��Y�d�>F��9gO��u1w�U������'['�1��FWN� �Q��T���F�Tu��;r۳B͵a��<�' ��pL��<���s�iok��T֓-��lKu�x�A�v h�V� �A4�㏀¬0�d�/O���@�4��z�o|�<���p��i¶�*����Ǭ$�x���iC=BO�}�y��s�1�b��I����Q��6��G�� ����4��ǹo��M��A�j*]�=��<��g�*b��j�)?��I���*A'�K{��g��o����9�����O�"@�Fh3��:�Xr���t�7���Z�P��8�x6�YG��E�g���q�gG�Or��7��H@�W����L����V�d�ۜ-�R礎 ���*֖,� z���*w\L�%�6�O*�@�w�Eq
��T�j>Qോ����\��i1^��_>�R��J��ޥ'�y	]ݺ��z'x�������Ϻ�ʆo��}H�{�������ݔ7���.`ָv��}|����Ca�N��^v|{R�H��b>���MbbtU���&��l)ӆ"w5�� �	�K$�=]�ҋp�T�\e�"r꼿�_x��]���|l��
ƛ�P��mKjb�?{t�|���PU���_+<9�cO��|�?�6�2pB��$�&|~��(U&�[����iQ4�8f�cj|��7:ix[IHB�9��(��{_����{�i�k��"�*m���>�>k�!9>�)�N�t�	}��U��i'�m�����Ӎ�]Y��*ن����F���
�	�(|jZ�-��U���S�a��;������D:�tw`i���)A����D$�wN�Yq�t?�����5��M��1�4TE�6�%u,ߩ(;"jM���_r3��L�GdA�M��_4�������cz��ص����ql���=�����>d����9MDiE�,G�@-6���T�����0o��~�����;D'��u���a�;��)������\�1
O��C6F>ఈ�Y���C��S�fH��!0�LN�S���,EVhh��`�,����Q�΍:-�GdG�%��qD9�{dζ��l�W��E���Wj.y[����b��dY�g����(J4ؚj�������_uIG�(��Kn�z��=�5��2 �\(X �M֯��0c	�k������&�����̈́%Ɍ�u*��P�
(�g���1C�!&�}���L:��<�nȊ�$���p�Z���o��V4�G5�����0w:q��0�Bo8&�?��	�x<EkH�+�����=��(	qJ��OZL&Ћ|��S�D���kj+�%�:�%就�T���%\�5��H���m�)ɪ��a`��J!��/�T��AS�z�@�F\U����v��K#���C,.߻��W�x}�&E1uv�r�T�P��J�(/�kU���aC�"jpq�\0�Q��\ ���x>�Un&Gt���x�1j���e�B��L�n���X7>Y�r���f�؋6�9GQyP�3����jX�^kiF��u�r��D�fxs�pQJ`�'�8ٽ �+|1��\��;�O���/{��B�	�Cӎ n�I�z��#�!����k ȗ*$�~B+w�ܠ5�^D;!ս�+�_<R�l�ټ�f��4hR�.�;-j2����ͷ�z�)	�4ݰ�D_�q9��)��d��e��a\��m���7v���Ctʴ��K�S9���t�
e��4���e�;d����X$]���1R�i>��̝��\�ѼX1A O
��]��8]��*Ԅ.}TEe�[~C�H!��9�*X�XZM_eS���0��OƾU�H"]rMqB��M�	Q+[����){��q��G/u�ԦM�?���\�dTZ�hZ2��d8o�[|5���"�r/��i�t~D��j���_ �`#�v~QK}4�/�Äi��l�n��b� �ͫ����G� ��`�VDQ@/(����0܃}�`62t��gY�|�ɛ��(��j��̓�u��B@3�˯yy�Y_"�q��2sy�C��[�h��NRv^�����G/��x��ip����:���Pk`�1	Tc��_�T��F����+�Q�g�nr���(����%�+1(��v�K�F���ڦv�HX_����K�z�*�)���[)q|n�*H!����E!�xI��޵�EvL�_��x�Qib�E���v�C�
��v�L�dd-�{���e����'4ݺ�����+�t9���P(��L�Y^�i	�D�6��f�>wup�kNEzi֪G�0��Y�7J��n���&�%.� b�%��Ӆ���(���՘(B1rT��a!@u�!O�|Ҁ:�ݱ�0�0]
����\y&V'h+���_��"��A��U��W_�Q���Y�c� ZM�[��v�	I�=(Pݢnf�ŉ�*��PqZn�&c�t�F����O��linrĴ����8ǟ�P����^�@g<�Lϼ��l[h�
4�a�x8�#*O�W��>J����*�Gv��(9�&����$����?��r+��y٤�N5�jJjjCo]�-�:��e�%�%yO�u��)��5�r�!1���ܳ�gb"A�urTq1��-!"��'�q8��p���`�BJ��+a���/?�߼������\�UF#\�yXp��ziB�>���uYU�GZ)�әc�bV�GsԮ���@ü��Ҩ��Ign{C(I}7,�π%>�J1�&)C4����Mm�� g�B�a�X�C,%�4*ޅ��R��-
��52^��~ |P�W/;C5$�y,WP�;����5��岄*	$L���j���=�sS�
�P�J���\Ek�2����k�o�1 p�� �9X���>�b�(�lM�zF3v�<�~{MeI�U��惶�Zjv�&W���d:�����u^�#? Y��Ub2���X����ܝ�C;	+`j{��3wL�(�<�0;��}Η|]���|-ú���0�����nhp���26ίwKE$�$ڂ,kӂ�V�����OWk�]2f��Wn*H�]�I�(.�F����ֺ���F���e����������q�����1V�;'A���͍�!�r��I�5}j&Z��oU�>?~�' �G��&B���؝XL���7�u�J����^sGl�l ��Z\Q��EK��Y�R�[YԵuu�,���Z�3?��&��[�.ÏT;��+�*��ɐlP�w��Ժ߫y�˭��)���BR����#�R#W��x�C��mnz�~x����VqJ 0�b+����`u�pA�{��]d�$�_�[>͐����В%kL	?�3yLsD%����B��m
����{E�녀�)n�yA�9x�ε�����D�����R������kUu�-U���v4�����~Fv6�fDa�ܠ0�Y�����{�����
 #6���T�)����q��ʓ_�[L���|$�W;|B4�T���CT|9.�o�S5���,��g��E�1�9Z� �z�.�YF�[��D�qm��̄��V����^�N ����@�� Y�eӈ>Ø����:nr^�Y)ǎ2�HM��9R�dI��[� B�gsN�+v���>��0�:ɜ3�(��/t+"��(_�!�Ewa���K�=�'�C���mƀo�gi�
����U��Q0:a㖢|y��D�g��$T�a�Z��l�͢r*}�kD�^pFr��m@�ɋv�O��#�
B��nD�Wȯ�F�(�b(0[=+���8�L���p�;�<�V����W�ף��#`��6޵&��ϸ��atҌ� ��
�Y�LM�C�ɼ��|�Cf70������c)�v��iad��`p� ���ZM��L���y��nr��ܚ�zq0>]��O���رG�X��>$��"�Gr�:Ry�J*�7b@���QU2�����3�!O,��\U7*�Cr��%f��b��{9n,^��U`x8rs���6�L�V��Ml4����f�aј����D��t�.�D?qwH��nR�f��*�k�c�5��!,���7̗������ҋ�6��kT}7� 珺U��������l~6{-����c�_�|�k���@�6&������VTD���MC�ab���* ���ɚ�]�"�;D�I�:���P���@m���5.-,6ܪ���&N���cw��/>�����{��L�[h��?�nZ	�<\� -�:SD��>�ю�j�d�Bj�|Y�TG�M����t��M��~������p�"KlO���[����R=)*�W�@<K�P��@�����$J��V^���f�`���ٷ[A�j���|q��q��Y���(�Q��o�T6�_�]L����V�����\I�9�4����}>���H�d��G*KlkUc�G�jKp�۽�=�������/���w|�L�>,��+�
^��g�����>x?%��tis���;J	���{j�Xʕ�e��K^�+#��LV���PŴ�Ƣ�i4�S1�l�]?��gw$p^g
m��i�t{o��>*cINu�G"P���$���lp�E\=)�iKv*7}��T"O����IZ�os�u�|ϊ�݈�ݸL�l���ȱu�c9��V���;�*��~I���C���)�����LK�t:++!f4�ǗS�͌;y�