��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȠ�>q+��q�N.�T}�:\K�%�"ԒŖ�9�ha%:���$bfrO_ �,K��q���X|�����_{[���U����{)��*��I]<�֭`���[�ɖ��c�G�`���Gu��*����eS�GiE�ԋ�@�h����3�y����.م������κX�&����;c�]��q�'���S_�ϼ�KI�"�Q��G��8�<Q�6���؉��'���ke���0���
#,l#��cYd�;��1�&a�1P�D7��@a!�8y�L
Jo(�TF�Y�-(����D�����8��t���-
�(]�� GV;f��m�!\��b{B�_��l~���9��Zu���B�}��У��"���˩-���p?u1�Yl�Us hk�RtHfW�:�ޡ
�^����&��y�����������:]+"vS1��y�Ig�$Q��=������'�`���.���o�6�੨1���ѵ��a_.��g_asʝ�g�4��3��D���F�Ѭi�L�$�X^�	��FP�f1O�9�'"n����v(b��������0+��㙘�s�́K&���G�ֳ;n զn�r���Jy7��nƛ�J���Z���VܐG�Xi��xMB���o?�aQA�Z+�D��\No��Z&��jk�d���{U<�\�U`G���)3�s^Ǥ<�8 ��	��|���8d��`��9n��Ϫ�S�N�e�1 ���`��S�0.΁O�5-��"zW����=�ռ�^���G�D�//�P�X�d� ��
�F�L�R���d�՞��MtN��� ���$�w��D����FԌ�B��� ���g��a������Dk4�f���{�����6_�.>zH��A5nI��V����q{��}?D3��b4;i��*�vݴn�м�z���F�m��m��zDG�GP�#����&��q�����ӖC�ӾC< �hӈ�a�����q�౯��rF���շ9���w��j��+}&/��W�٩ W5�p�g�Q�?����>ԗ384�c���`	����'^���6�e�m�"5�gԨ���rٳ�Fڃ�@w]w� c��iP�)?��y�{��Q�F��$������Q5��;�'�a.��e�'��ܛ���S�~=����S���F�-4b��GZB������E&Ơn��A�6ǁ��.��8�2"�������4k���@�8�Ħ��B�<o�ǲ"�1����p���C�ԭuCԲ��:�7'r���ǦH߮/.Y���FCd���؞f]3��0̌��lx�[�Ze�f�O�&����n�Vî��K��YX�N�,����C�;�Y�A(��O/�<���BZ5�N%-��r���R0��l�[��~o*G�n��ձ�
y�5�x^���Y����|{LT}&�
��4�xE�[Z�\�@��9~�}�G���d1c��3PW�.�E���������=/��@�d!o�����т�g-���eY֪U����H����!�Ť|�sG'1������T?�;mY�K������H����e���/P�y�DS�[}��ASy��v�$*�TRZ��O�����]R��Y��ٹ�g�!�[ji��;�zs�a�a��(���K�K�azS2{�%�������;�<��ϓ��c}�Ȕ���/=��A@'3*֓�%�"ڧ����
���$-���j�m�b�Ƙ�"��������j��Z�o���B,9��UK��!c���G� �_-�����}�����3Q ��jm���If�-=�iۈ�$mM��>���u�C���4�6�*�H"(�D�24���Kv9߬�>ુ~�֓��vʡ5�ﯗw>��$&�-k�y�}d�E�Kg�S5�n�C���� ����<�c����Sa<L1�C=����z���]��p5�V�qg�l;~�es��)af� 0�5,�)�V�藠�'�����-�rǇ���œX�ID�يʮ���.��Pu[B��X�h�9�5<	q�Q���c)X$f3d�h��`����c��I��I�S�j���: \��́�3�@ѻH+9-~E��8PC��\&9���8�P���@�W��H~���]{Obb��+2��%�rOá�Ά��P�m5�CR��h$�M���n6��>���y��#ź�>ѹ�N ���q�}K�P�8��w����Վi_T�bP��Dqc����#++���:�כ�Ae��/��|�tI�e��U�d��Z�Nx���ˋ���/|�P9�ӗWB4��C�[nL��IB���4F
}	��H8Ss� I$�~���=��0���8u���s�ih�f6�3GHl������I���!�x�>K[*c�Y��.+����� �	����� �����s�ټh71��\P6:=���;&�+ݭ*]:�d���W7��"H�15p�GQ���*���/!��c#L�O.��$Lk��x���1h�$��,�+�����7�kj�|�$0�܁졟�Eֆ���އ��^��:��L�Mo�[o�^R��?�@E�o���[/�`L����h����
Тl
��e���oV]�=�kl��WWc���x�Y�e�R����eD�mbBq�E'�/�Fn�?�|��EW{ᅏv��p{��lYhC3���.zt�ܿ����L��'�7��@�����(Y��V沀Ȏ���jvG(syg�\W��s��Ys\��8�
÷�1]g'���~�e�9�d�Ѽh�tڅ[ -���?��_��x�zgִI��r_��<9�=�mj��:Y�Β�7P!(���pLtJ1���<[.?@}���p�w}�������k-��i,o?�R�-�0~�[hL��ɸ�'ft)E\���Qp ż�.��������P��[BlG_����Q ���|�,��<gD����p.0 ��>�~���<D���R���>sB�Ă�y��
"旺��,�O����Wܼ<+?"�yE���w�ʙm�-rP�����v��Odnp$�-��R�|k.��^4��p��M�xKf�:b4��=@Y����li3*Tj�=��Y�M��&i��՟/$�;�j�g��ò&�'�ԝ
3ڒh����x^�p�����ۥ8'���5��,L�%�؏]�*5����yk
p=�}���KlIf��]���)$G�MB-�`U��"!�s���Z�&�R|��#�)��s� ��ܒ��ܾ�6� �u�B)ӌT��i��Ϙ��|�� ������-a�a$KL�x�^�ՈxE�� ��L�fk���r1-~1��`�c������f![��cu�Pgx�h'��A�0 ����"��-ѵ;�ۋ`��H|��!�B�;���S�����S�Z��6��Bb�:�{�t m@,�bޞ)���@�4���z�8�J��f!�BTKh<�n���d���M������Q+,�s��ɽ���`S̞���/Y���%Z;����
��!G�i�"jĹ���kv0,v%DA����n͢Ad4�!�?ϵ�7����i\�rKu� Փ�(��%�昲}.h�<�A!����Yϊ{�R�XUK������Pp󹼡��f*f�0_8�EǢ��Y >�R���8L�~5|:W���y� vj_錍^2P����u��eT$�BH��T'T�uL}��� ��pGU��9��W����
kp&��GZ�M�Ab8���R1Id��X#��}��*�i'eM ��n$F�ę�jr�f��e��'�a*Aγ�	�I�a!�L�nrH����`
L��6M�m��� آ�4���M%� �a% �Qm�@_��"脬C����sU��@�	4rW�"��欒wKق��y!k �L�v	E�V�����W��R�]�ғ
����)T�Ȫ8F6>�sb�X��D�}[\7m����O�m�R^י�ݑ���4��VY��5�G�zD�^<��B� �I%j�Z�w�p� pͧ+�P9�[�4+�g����^��t���=q�����*����CV��U�g7 {W�.' ��!67/�b���/	�ξ����ڀ[~�4�QU�k9��a���y�����+��E���(��A�Տ��Sܦ��i�͐�Iz��@��#fc��F�����Ww=e��L�!�o0�P�H��w��D!m�����k�]��*\�­-���j�!su3�����++�Z�rEa;��Q����<gw����O]@횟��[:��E�]x�;#(����cpK��L�{�]xG��r��>��<;Ƥd��jEr. �S��쟞��$�=��C�1*�|�.�i��/g�����@�.��'��GZ9�-T��z�:�P��.N�I�G%���=���9S6̿$�hj�в�������{�����g0*~c@&N�[OJ_x���_E�Kp���?��_�3}
��wz��߲���3~����Z�G��c���������M�ɇb��O���+V�z��4���j11�.�{&��I-g?���m����%P�%q�j��;M��h�c��g�T�Etg;"eb�$C��q	H2c�3�U&W��.3�xL�f���]�d�M�	�.�I�c�s��F�w�۴!�Lӆ��Oq��N�:ia���R!��ݱ�kQ�.��=��%��M�dΥ`{(w-URց��S�R��,���Sh�����[�Y�tXŢ��،�:I�9ڌ��gcĐp9R�\�D�cK�Y��[~�����M%Ь�����.6ir��4#:�]�Y�(>9�A	�h�����B{����	��!D�]�]!�]���@��@�-�Q��K?r4�(zP��嫚���p ��G�rt����%��	�$��$tl�9�����T�u��;J=�N�����S���Xk�G+T������R4:�ܬ�!j�H����1W�Q��-yX��+vƆ
�
����<������t$(6>��"�n�D�zX@O�7���V���
��d�B�R�{E_�r&�L�Fc4��ߦC��p������Ε� 99������t��.ң�xL�$����W|(C����J���;C�;�����i�0���@��'o�{�<�=�fH���v��Zû_�6.JYtg��I@
�)˝�"�e�\��rjY�7	��	�
7l���e��5qW�x+)a����U��M�A7��g����S	����;��i�0�L�˭[y�E\�A�1�Ug��a%NX)kQp��2fo�-*U�2�z�w�i՚��)�[��w�2|�k��\[>gmﻧ[V��E,�����W�h�l��C3�8�'�Q�1O�f�>��lc������-����`�­��p�X�QT�\�b��x���)@E�ed�l@q/'�P�)�bͤy����Ο��Dz�ѣ�-���$�y3�N���>{�
{��ܥ���r]���|��,�x��u�l����r��H�i����n�(>�Q4)�1Su\l6)�1�N��D��]��!�L�T]�8�����1�E�
xh�9�h��37B#�H���ơ�1Ú,lhC$3�A���t��F��W��qɀ��^4���S�~�����Jr�
=~�2���?\�Ay�*�S��"����a�Xʇ�dg�ظ����zpGkQv�G�<8�KWzwW�D��������D�t���If�y�0�ۛ��#@ɝ�����C��8~s��y��H�����0_\OU�����n���ώ�E�Hr߰D#���
L�WfX�'�)����t"qt:D:�A����ߟ�%�t�ao�ZRR
��`�b�ɶc1P��)��EZ��c�95�Yw�|�Y	f�ğbc�Ѳ�A����׾%�KT�� �_���&�ύW���n�/O��V�V1�.�O2���BD[ ᮃ��I	Wr�b4X�ė�S��.����������̱���G�"D�`�j�g��c�n�q}Tq�缳���p�	lã6�(R�����PaH�
c�ʰ�'�с�u�"�=Ƈ�'qQ��_0�Y���J��)`�zږ�D�*w�!��@.�>����SJ�T�@��[�Yi/>��UN�:
]��+s�L2E�PV��SP���As֨�hbq���/!T���3P
7_�$L��y%��ކFb�\Nu�7��s�h�x�F8+�-B�1��,�����H%r\s�<̡�&��m���"�q�T&���Gud��OS�z�H�mu�+��b/]�x��:yz2 w�8Q�h�ހ0�2�)Z�E��]�~(d�]�a&�wt_p���.�d)�l#͋�g�(�t�Sn�*���!�����'O�^���eY�Q�]�WI�qt&iP�j�/��/2���
V�e<�K5#njx�k�2�{E��xF�st��H=�U �̪O�s+xW3�j8
�Fȹ��  i�	��B�.!$��x7�	КH
�r4��iV�%eܰ�R���.�Ţh��6�`����*�,/M��p�fp��C���q���[K��<��=a0�7��~�RY{�C�q�տ����/�P<��PXL�ޛ��N����o *�QY˶��R�&�'z]X���6�BS���aՕu
�3p뤷v�ub��JK��i&�]@�{%ᅒi�� �i�nD�7�Q���x���XO@�m��^�x&I�#�O�Zo��tyt��Z����np��x��3����	n��J�ާa!�r�0�[> ����rj�����Xg����N���Im1ԣ*�e(/�,���"_�bhs$�s,<��^P���~��F&C�(�X褉�q�)��
�4�C:-����CP#���j)Jܲa\[Bg7�IWa �,��j����*r�d�����jdə�.�!D'2L��q���0����)�a�祡+x�����?�J�7m\F�.�E��o�l���8��hГJ���_y4g��8�R��HT4��U>�Eњ������7��B3��tԒdף�j�u�)8Q�a1	�E=6A�xf�^<H^��i���z/��n�,C�r�7"�6�\���vR�LE�72���>ڵ����[�"? �.�AK�-çO�yV�?��m����zD���T�&�Ñg#�L�l���6v�ЅB-�S��ή�rddRG��ڜu������I�v���mC���S+��7�i�q�ըh��ɱ�n��5���^Y��U�,,�5��6��w�7��)ø����k�>��|�5U�`���{3�1��c������v_��+���aD��=�O�� b�9�a���@h��
��P��� 5�0%� ���*Sd�KƏ4�v�Zm�[_���ޅ<F5�/���&�Ο������v�t��m��&�TuO��ŝ��?�a�I��MH��3�B}x�9���&$A�5l"�`n��GD�j�&�m��&�k�v�K�?��򟼊KG���
�%X�s�ѻ?ˈ�1��K�f�:(,2>��82y��.�tL� ��~�Þ�ӡ G���i�{�(�}trO�_�[��E��Q���Ðrp#-('�).j ��WC��ʰPTt��"�;��i���>'t��a�������3)�H%��	Y`�A���s8J.�l��Rm���=K.`�u�hQǨ�'P���y�_o�{g�N�H�sm5�Q���*1��q���b/?N��\=���f�s_QQ�^�f�v&�r>z����nDj[E�#�3�~/�&�ֻ���+@���4���K�~1?4����r��8w �~����o2���9k�QAz�#ʏKʰ����B�:'.�尔�
��C(�b^Cl해�_b�v��i���c;��( �O��W�Q��Q��L�F_Ti��0ƅ`����R�
Mp�"\Y��AO�&4�>��FlbJ��	"�O�������B!���\�i���N��X$&��B����^������ ��/�2���u���ꑙ�����7��gF�ߺ-��'�y<���;j��XM����g>��$^0����S�h;rn�]¸{��<N ��DJAӮd�:F�����]d��Yh�#�mfQ���S/��$�U�\W���v�	�-�����V���e�W�$5��8IQW�A6�S�� kz&
�����e��E���)��J�՜�H􎩫�[�y����F�n4o����ެ�ڒ�I���w5���rY�֦N��p�7�d^k1�����q)y(�Rg��Y�t���Z��R�/�1+���oLJQ���]�H���9�5��ÄH?���}E[��,D9�e~;���+�\�^{���Rs8���T{�w��8�,* r��;k�<��{j�q)�*�=)h��B�CCkN; �O��6efjK�-,:<^�LI8ofS3d��=5A  �I��q�%���	���ߘ̋�Il3�3֛����!$a#̎?<���@U�}.�aG�"�z�2��(�����,	h����i?�	?n/��+wGɒԲe�.�L�KU�m��#u�e��ӱz�����6�h+XZ�<c�5�
�%fe�`��~ͬWwL��z���j����,���D�N ���������䒮ѐ+�4��k���օm���A����
u,���O���z��j�@��"}8#���n�|˜[����鍂%��}@�h�{��"�`AF������mgB����h��=(E��NPO-���c5��RX��MU��4Y
�wWdl��(4�1]V#�r��=������uk�2#�	 Nq��u΅�L��>Im��('vx"�\Yz8�^�Qv��Cښ�M[�L��;���e��w����NwMd�ռ�/r�M�b%�0�cdtN=_�s�5��V�A��e�mM5n�\��.H���	�M�5��YY�-��
�k�Gi�f�WEXZN��͗ �'z� ]���e��ks��	ݸ5R���5O�w<����5K�lt������6�_v� ����x Λoc++Q��t/ �6�¼�t�7�����a����� �W�����l�r,:��f�����c��Jՠ�9���o-��b)JX_���{ap*Iл�*��!�&���%f��[�U�lx7��Oa�
}3�vl���MH�@�N��~0�w�<����.�C��v§���AE�e���L���L5����16IohK�s�:���~�G�m�&F���1H"�! s,F�I��#��òV�a(��5Vɕ�2�.ctB9�:�SM^������
�cP4�7`�B�'�
_��0`}@a?�E:H�ڐ�l
����?q���S4#}��79��*�E�����?����̿$LT��O�ƓP3u�|�X}r�A���uDK��b������2�8�-a�'������{���@$?��$,�C�S��J�/�$_z��ZM"�W/�Ú^�
��{��=�G����?�8��:C0�s��P��2�H$����3���P�
I��BR����U9��S���ow�}���_��C:J���*R<�ut� %�"9}c�6�?K����ż̠"y8��rb�r�FH���]醱Oaxs��'�&I�My�T��}��QΟ��hޓ ������Al�a� ��L�qžeȡ�O����%;�\/���vf�T�]"F\�	i%��b�Q�TB��D?���En�6����d.���ޙ��qG*���!�Yx(��#]n
���Q�Ь�v`~���''eL2��+�,_N�s���S3g5��/bu3�Y$g!��y�jcl��й-/2�h4��O�:,��ƶD=pј�dIǀ��`�{i�}}fp�֏�eޓ�'#�\�ᩑ�ia����2����	�N�-����p���j_�1�k��	 ��r,�YM�;L�UP��ܨr�#Dtqda�K�+�-ע�ŵ��	0��?=U9x���n����S�0�F�������A��$���mA����H���%�y��X�D��Dȴs���g��su*�ш�I�����!����Z�7v�S��^Y�(���?���i��`�M�L��y}��^v���ڙ6�Ł�8�hb��p����{y��I��hM�!�۾^ַ=�s��XhZ6���Y��F�8$��@;��irȌv�g���M~��dRM�M��[�e,)K�+z{�-0��ϾȪK/5(�i��`P��l�W �.�jϱ4\����c�m,�r�Le��?�2�@����:�R<���Z�UP��Fx�i�m���Fp����� t�gKJ�恦qo:!�%1粐�P8	���n�֛F@F/�XI�A�izP�bK���v$d�UW
�uQ~!�8��>��sX�җcj�X���}r��Dz3�TS6mx����a9l�_5a]�q���n�+�.�!��U����U*y1�<RB8��X�Z^h���;X�%e�������N/�c�0�/��pe�PN��JB��(�+M�j+]�7�w�|g���t��R�CD&�>Ѧ�+`ÂL�{h� �H-�3Bn�q��OV�H�lB;�8��!�b�QA�]s�|�6x�h&�t��\'w7w%�J9y.|oH۵&� ��b&1���&�fXc��)P���Ӝ��tk1��N�]���nNMI�PJ̖a�*i'��͕�R_�1�	ȃ7�T����ZWm��
	�Ѭ\�� �SW�o�rјR�����6�/�<��8�G���{���#�6�� �<� �|�����/��֭_��[|`T3I,7����}\���5:]!��$ 6__y�ٜ��{4z����������5xA�u�
��x��$*��M7'�2��rA�6_� ~�'�D95�^_�`��kW��}B�M��4U��Vn��ǒ0 ��)z ��b1�.Ӄz�w�&�{.��(�"�w��L��M��di����*4|;һ>��dP���V��!XCK��4$�K�>�� ��B�-�p��id������(9�Z.c@���XM�2�y�'���"k�����79}��d����&���kJ�)M/FLh��~��	2�I�;�w��nV!�<�!t��ݬ�� �+���|����_�f�-��2& ���JZ����6�um�ott��|�r���6ϐ"t�(O��o�ͬ'S�4-�`N��C�@IO��<����탘؝�m7���-uӸ�u��G�
k��몶ϔ�M8I���Ph�/0m�ji�8?����z��4r��`�q�7��r=9�{��]N��Ī�O�[�l:�X&�B"BǽئYo8�\��D�[We?���FQ��_I��:X�c!sF�T��v�CҘ�[+�RM3ʮU�޴R���?)�+S-@��i�i�|-�������jx����h}h&��t�ߕz��I:[��S[�EX�Xu5�T\SK�Z�5$��u�#nY�-�����!�m���=�մ�xB�BG��C'����V� Π��}�u2������MIF;x��(�c��^�v��Gf���)�;�L��מ�Ϛ3;��}�h9�Ʀ1��q��u�i��9��|�9Bq�%�$�� ��A����;mT�C���S� oI�3L�M����Ʀ��.�@��t��|7��Uȉ;���O,O��d�dn���!j�`$��а�"�$<�J5g/
Y��߅��?1�ᛤ�X�����p)����R$F2˽��ű�q�B_��8�v5����4�9䶟YP6�V�R3����%���*����O6�xo5'�7A���!�3���<#3օ��B7�.�y�c��:a��9X�7�|K��S�9��?��#��I��Xڀ�b���ʱdϰ��&����rt��ٞ
�W�L�]�ḋ��s+� `VilB��@#�ȾQ�}�\���	G��!C�艃�Z+�if�ٗ�{~"w!�>�<#�T�8��\=�q���j-#ڏ����%(��$+��)]������y�}��X��W���:Q����MH�͞?��&����QX�K�V�}i�!��������h�Y�2K5"z>�9��?���-�B|���~%�W73�H Y"�6uQ����G�V&���%��7Xt��_�7�c�k9��__{y9t:1t���|����1�{�7�(�W�P	�c?���׉��)5��{�T�j�J��@tp�g�ɡ%��M����dh���|oG�g��.^�+WR��3�;c%�5���$}�N�2#���RV8Y�S{��d[D�����ķ��0�:�ҁ�p����3è��S30b�ф1~-<�?m�s&"�c��+g�f�0H=�\W�C���l�4�N+}"TC�q��?*��#��y��L�?��ɣ���f*SKq&�����G,�x0�.��(�oL^2J���h	�V�h�5��7)�]-�+�\Gw��{�
�(7XĮ8N\��w��2]�b���!�=����Z[�q����ek���	��Z���)ٳj����Mʇo�5�Q�%H�e0N���,b��B�o	x�8'�c`�@k��4�G�ԺG|,p�ZzoCLx�~ONi߆��E���H�	Լ�L÷@��#�B�ﰅ)W�b��q�E��2��U�<U)H�ū���)IW��lhي����'u�������C��W�l�d�MZ�k١c��z��:5�+��������1��p�QAѦ���&A���1�E�QnN����!02i��i��K{wt�����~���8���I��	>TiX������-��]k3�}a6�IGHzN��!�9��r������e㐲��`2,?�@6�#4铥MVo�R�hJ�˪�����	�)(�Z+�;$��|34D7���s�%cH �/��]�K�u�v��0�w¼HH�L�՛�]������Y�{n�+�q����64,>����ݕ����ѭOﳰ����5�e�q�����@��	6��:�vn�5��O�Mp�RQ1LK�4#C<P��^f�-Ζ��=v��`=�e�M�ޒ���:�W#�9��D�𸽴�~Ubimk��Vc2�Α�+~�"��=�w�+��u�� Ϙ��!m�1�d��i!H�b�(c�D����r�E�Y7q�p_\��p�QR@J��V�Rx�s�c�O�SS_��T�O��\��2HpFCP����V�>�N얋Ӫ#��=�wck5�lʁ4�a��n�H�Tx�_R�%��	�]�4�@E��@����R>9�x#6���_��Q+�v����&d�_�?��������uZ�'/��"]�{K�![��2?>6M0���Α*����b�eKd�1g�1��nᘶ��F<;d��J�T��m]2q�rn����ȟ�{f=H&�d�a���9�r�J:uAˤ`DI�4��b��ܭ����k=�
6�&��=�eҧ�n�w$�JT1��0�DR7߬�Q3pH0&-BI&�4�6����������@T >��_ؽWNte�y�1!j��X?yA �'�r/��bMLcZr��-���a?�0FJ?�G&�'��A(�?�u!�S�ܝ�,����n�N���p��J��i'N���z��F��L��㥝�k )Ew��++0��/�P�5���BF��"��Xq�h�~�.��!�����<Pk��T�� 3י����P���R>��N�k#Ѧ$���t���ѹ���w��ҬX㦡�}��bv�(��5��{�N������ŵp[�ʳ6�e2̄�]�j�Ȳ'=m��$�����v�'��&{M�1�T�>Ff�Ż��YO��HC�"���$����08\z�0�����A8TD͈g\YO�Q#��悦@�&$��p�4�dO��ڔ� �	���vwԕ�e���	 &�%�ȟ]|VVD!K���a��AWnw��Y��y��Vj�c�ܩv#Ij���޼�lm\�X�H�v���Q�F����k{�|1�}]�cև�SHz>p���@ӭ0H%Z1Q�S���O�p�W!&v�iK���X�f&��� -f0{�.oYM���������[tǗ,�sZ0�c̐0\U|�b����׶�J:-u�)	R{0ᳵEX��d����r�6)�9�tUqF�.{����j$�͢�"�5��\���ޅ++��DՑ���q��h�����A���h}�zK��G�T@Ebg���W%�>�]J�Dx���*s~�O���B)]�Y�t0���VS�%�`#6#)��K߽��ߚ�Z�����s� ����dڦ,��۸c�S5O��\us �Ԟ�q�9*��r�V-��C恕��&���i��]��T�Q\�G��tA
%c�7���8���~�,���M�Uζ6���C���-��B� �����`(��@B㽐J��s((�.�{Y����#��%�E�ll8K���:v12�I.�\���͍����z�T�1���[
����h�TV��Y�r9t��m�$'�ҋ�����e������������/|��3��E���%��z�-��y�U�'Y����,���*�v���5��J\�`��j�*eDr0�,u_EC�_�\5f�,����P8c��V+�a7ʍ�͝N���l �X���Iz-�Z�?���ez5O�l�5�:�ݧ����G��Rǀ������ll�A�\T�x\�n`�3�뷖�.�,=�!b6���H��Y��3�R֬A��Ӹc�n�&D*�}-��/��VD�b.yc����%��W8,���ҷfh�z��|���J��=��C��#6̎����R�ǽ=�Bm�\%��͚�Jv�����_���r湇��T������U=��`��� ��RMd+���ɮw���g�c�*�ߣ3a���3�=z����	LI]�WQ����\�qH[�bB��<o~����4�bd
�7��0��wO@*z�Ͽn��J�P�S��=�=�3PfD���9��"Q���b�8ӎ�A�Z�9��՚����!�2��/�/m'A��8�������H�/	-�gG���T�m��_�u�t��}$�ѯ���{�Z"��<W�,������#�x���#3���{Ⴇ�r��������#n�!D��ҮqxUWu���"�.�Ur��������c$H���z�MNm� �r���)6�Z];&7���8PĀ��{ޗE8�I4��ZM���ޡJl �|�K:�o���/��)�,����u�ͅ��7�?
J��!�������$�nF��%qBM����
��n�眔R�h���+�^8^�}wĳV��,�~�0�՜�|s��¹VƫH��B{�ITt4u�ҙ5���XC�0[7X�4A��F�(�p¾��f�֡�L�˵���j�-XK-a�Ӟ���tY�X��r$�&�KЪ5SD�����)����$�^ ��-շ������*8�͛HU8f���R�ON�����6��t��h�ic�{��\��ۚ�ҹ��
 �#��R�쀖^ta�����}-���Fi�eة��´����<.��������hQ�Q@e��%�!��w�O¸f
��Y��E0ϟ�c%i�H�T ���%�F&	N�NR���/G��t�(�p\�E*��A8�W�[p߶P� Q�1W��Ҙ`�����������$:��YnX5T�ʝ`�,�2'ci'k^֋�3݊V�G�K�$���ϕh��� ���mt��e�д4ln�a+�/��~Aǻ���"�d`/��w�k;���>ɯ"���{S�z��"���j:R㑴�T$�3Z�;o>�OC;]�p��w�B�6���turO��pJ��-|�G�Ov��n�Ma���l$凕0Ǔ��s���4#�yC�-\��W��Ċ��Mp�_8��L-{��p���=q��̋�PDGH�C=�zSs��u��L�q�������w�q&�W��I��Y��Lb��T4���~����ʜFD ��i![�=�?<�*��x;���ڬj�irk'!R�c/�&��hP��R�P�-}i�j	K��N�V�@Ĝ~�a��è��a�Չ�����gTWh�=�G�\�żhW�B� ��U&��n�u��M��!<<��'(4p1d�1�K�Dm�t�'͖���^�x���]�O�r��qR���?g�b
jҥ�Ͻ��Fe�Œ�WNǼdE�_=�_u綠"?f�(��"��(���^���)��\$�<Y�4�𷼾�|a�R�xȬ�ޜВ;[��Qu(Ew�	7���O	��� �OY7�{�|�M�"x�3��GX�gB�Hr�K2����-x��Ndo�����g���ʟ�[j���dUB��|�������{-[��<}�����m�� t�(�
+��@�nr}��Wi�.����U��3�!�Bs?�t�AL�������s��_z�N����R�2"@%Z�g;�����^�wt����iRHG�O�e�H�P�Z=YUkl+ �pY�[�d���"S&~��<����g]gP����� ��_���`wMUy�>5R�?*r(f.�6t���'�DVW-Bi� Ҳ��P0R�������}��3��
�ɗLkh�@��"���w�z{4�� h��'X.�c�R��itHS8!G!ݒ*V��L�k4Q �'���;�Xt/���9X�3;W��U�����3�1�����`*�"��t���7��P�3�<��
���Y����H�����# +Ȅ�6&{�Wy){�v�{����A|�9�B� ��N�f� 7V��y�AL�h��; �X���^�(�"�n�>��jq�A%h*�����>p5Z_��Nw��
S�9 0R���m��@�q�A�#�߳t�'ϸD�瓮�t�7}�����!�k�]a��+�$�.�^5bѢ��� ��5IĊ�mQF�@h\���r�Qe��ؒ��S�����h"4CEA��y��s�UΡ����{�[l�=D�ٮ�g��?�%Ӯ��& {ϙ��xW�{������;K�of� �ȳH၏�n��7$|JQ��y�r���Ĩ���� ��Y2��00��D�K>�����g6�D,=/�[d��5׌�u��{ ��:����÷�#_Z�9�M�� �,/�&�k��>i@�X<aB���P#<���p�˃USh��l��2��J����n�8�Y�¨yg�T�[��������c�(lv��!)T�䝷��1y���ra����YT��3{�Q���T\K��@�q������-��5�Q�#N��S#N���z�S��i�Ux%�OD: ��!�^��~����s���W|o�g���E����7����D��g��|���������X+ڠ0�Y��Ɍ}0�>A����灁sW v4Y��	��P�waԞF�T��iԨM�����2S�%�k^��[���X!=f��)�k��������',�C�j�Q%5��?w}�]�o�ULD��RfT�f����紾Rim���w @J"^�L#]�w����RWs����Y��sN���_D��6*�&x�Ĉ}������^��[x���Zȹ��FW]n����ŗ��T�W#{����i���2�`�ϩtfZ�����mC�� ¹�./�4*�P]��ʍ������lh�(��iFh��I�^���a��ga�S���^S>M�Fѽ���_����c,f�R{A��Ƕ�/�:6�+�+>���Գ�D{h%�I{��V�N�Y���ftB����	?�O1��š��nu��o�>]U��9/�q�`nڬ��[K|��Fb��9,����~����z{"���a�4�1�?����s+�9�M���,��d��mA�B�J�����;��=L��&.��*8<�+Dp�J�KA��ǐzJ�9�Y�~�!�<Ϋ9����E�|QG?eh�!N��/n�2��?�o�I ��h�- T"�[�8�0����-�͸&{�,�?K�T��c�a�Cm2����՗:��~rE�v�h	9���F�:����#6�J~p�V�K闟6�<LF�X�8;)���S�6�>+���8+�
�x��^Vcm��ǤkǮ_�m�~u���wzH@NU+m��^� 2\�����������6��1��o�ݪO����@x�\�Kځ�S!� ��F�Ƨ)sϢӿ�}|� 7|`G9G�Gw��E�إ�SZ�f�<3�SqV����(b�,�;IᤶA��}��M��˨�+�^��:��JN�3��}��ݧ�G��\����g����-���-�=�L�[�J}3��{&���;���[)�����߭PO�µ�Zq�ou+���g�<��7a��x�?��j~P/}u�1KE�v��(0����"C�'��lK��iJs��Rl�N�u�/tO�\�!��^5�C3�+�/|��4�̨����֘bhf����SS!2�'��Ša�z�̢��!b��|�q����a�\���q6�����.\+��sh!�~tbA8b�w�+�T���Z��a�����<!m5�+�v'y'���E��8XF��@����H}�n��s�$.n�1���ϵ��W��UT��`/�_�:Q4�U3	���l>Slt��-CN�XeF���r�+
�8Z=��0R�2{���Ͷxq��yrx�ŀd�����e�����\c=0P�^D���<������ ��&�aβ��0BE���Cf@T�I�v~ǃ��F��+�R�l�)�{���z����HK)���r3���?��C�UGdK�;���ܞ$��z�)�> ��|k��U���G��{��[����?T�D�:��	<S`lK/ռ/� �s�cS	��'�|�{_��|��s��H�DK����X�!��2�������p�"w^����R�Sd��BS%)~C�M"|�y���s$W���@+�9p\���ج�d��o�1���ߤ�Zoq,. H�$��Qm�M_���ˍw�$Y�錀�W�g;�c�!�4�d%A�--m1��#`-۵�ܫ%�=��,����Ȋ�0g�lS��L}�Z5_(�G*��vڪaN%%m?��S��hUd��V�̶��lW�@���̈�{��豺:[�q-�#�� �n3ޠ�±�[Fpx�Ε����y%-�PYcO%l��Xz�6J0��I�|i���﹏*�0�^����HEkkŖ̜�e��E��i��h%?�rAn��j�c� ]l�~;�1y�Q]
8�3��qU�2F� 
��u�x�2�1�Lά2J�e��3K��\������Gi�f��� '�3���	���*{u��Z!��z�sIVBy�U�8�0�=������ճyW=K{�4Μ�fx��(cLK����ܟ�ހ���g���c��`��O�{㻪�'����.����咈�n�V�&)���}��{��%�Wy�hǳ����xr?#�T^�k3>\�Oְ���Q�*���Ĵ_@���5~�to
Ik@U��d̒��F��'����v(� x��Y��D�?��q���Q�9rұ��Υ��jGk`��5�#�(�H�`%�(zX�K�'�޺�l�'�ᔖ�}몶���3���06A���/H�t+���rg��6�jQ6A��M�_]�,U(B���G�$�(���@��,�:��T"S��"�_��F��.� ɐnf�C�9�5��5�#ؿ5K�K^�o��rF�Rx _�H�Kr����%c�{'eJ�(d��=CZ}0^��K��L��G z��i<S�4q��A��G&7\���[��7e>��ٛ�-�c�W�J���-����}:�R��Bk�ȏ}��Y�m��f~��Y��ȭ4�[2�td+\�i�P�,�1��3��_[9��֍��%4N���&�>�GIy�� �+���o܃�]���R��=Ⅵ0�QU)Ӗa3ez�b�c�ː�/S�4����Ӷ�K����Д�F�B��e}�e���'�i{���U�_)l뿚!; q�fXa���)i�nl�r����"7 v'}_g�qPEK�����h1A1��,�w�I����C�.��H�|�y�_�<�y��<�:�c�3)�\K��d�Y�;~�l
Q�s�#��P �3��M�1sg�H�0< �m�}�Q����w�:�.�}+'�(%/Ⱦ1��<��ߺ��ˉN����t"�qp�#��3�XX&���C������W��x�KD�`��#�PvnZ�l�)�F�+�L#�/�oU�E̔���$ͼ�߂
�{�=���w&�ĩp�n�[�pΏJ�ˤWB���h�RT������i��M�����*+b��F�o�r^�������������/����0��.?ǿ�P����<����H��ަq��/� �w_tVkҼ��M��ف��lF��㭓�Y���r�.�uW�4����1+.�޴A�#k86;hf,-�t@Uq�a��w734&�W�S4|p�plc��
�*ca-�>�z��c������藋�TG��Z]�^V��	J6�`��n%�4���_�5I�vs&Ly���T�yD���1�BK֘7�Y��P,C?�ټ{O�����Y���\PJ����r�,���$ӎn�Z�:}����w*�Xn�$��9?�*��pd��h^85cq�t��x��&t�b:8����1I���ϳN�����n�E1�N�r.�+�/�퉨KG�O���o��l����\!K�Y�z�C�2gQEf�Xw���s1�3��y@�3�UE(c(�2	_�*�9 �"�8��m��i�%8�v�E�t�$�,�CAnۧ�.��ٸ�[��3�_97������E궉H_����/q��L��,����7;����$:��CU��ϯ��#�]���M��mqP��WY=�x��,}��;va��B ����J��[u촅�F�u��IF�K�VTvc&��~'{
�����;j#͋L�9o����:O���d]�f��<���/�qX����0��
\�6+��l��p�Y����s��R"xT{^EN��1G=�=���S>+�(����Z#��Wb��r<��&̈�-*}ctg%��R߸�$sTϢ�)a`b ~4�xa7��'�K����?ĥ��*�{=3O}zM���Y�I�5�n�%8V���+>m��J{�� `'�\��I�G���daD?ce/\VK��ضh��+�2'h���C1N��>��i��7�J!�r�e�sb���9��{
��1��}T�zfƬ�ТI�6��w4�K6O�U�M]��Ѩ676Һs�י��?����P�C�G��W'�ӎ9�L�|�I���ʽ{�)P
�cu�˘�]��\2S\`����hzc�}�oC�cޱAG��8�X1�k�gjx�NCsZG�������î��$g��O�qF�����G�Ih��?9���`3Qӝk*�1��9Itu��v�B��Ys��K����4�Z� �2�ߍ!7 b��X2m$���~4mN�A��U�'O��_�=tB�"�����h�&=���K®
(2$dw$�uBmZg��.��U��v��"�{���V�]Y�eJ>%M' �%����C�:��5a/7FIt������ֶ���.X�/�+��W���]_�#$�k���#�U��'�5��<��h��J�rZ���Y��!��������<�C��F��5�7�+&vI�8�Ϗ ;���+��@P
d��������eD`��/�
���ω�}ޞ��pZaώ��`������5�AN|�I�.9�~�J�w7Kj �0x]�?�oA$�mf@����})l�I��2��uIA/Wsq1�q+��"�㫬��w��������N	�X�z"���	A������Q�?��u��Ah��>�@1;�J�[�����*:�/�@���N�*�Կx�c�O_�Q���+o���m�ߧ�ݥ�Z��;�L#LD������)<+%b1n�T�=���3��ٹ�܈�ݠ��c��������8�"���j�I�N�f���|�S�"�_�!��ڴ�����5��o��W�RƇ{c��x`�[l��eC��w���SH�`�o@��]��g�-���*	j��&�'���aɤ!\�YxҺ��ڏॹ�B�+�1���r� 6�\�*���sM02�Ia.�䨮�+�GJ�?*�(����V�ĥ��@�S��S���aJ�d��ɻ�'a�¹{�G�K`���/B���@I�p��=���k���{��q'�&�oYy�%^���W���u�I`UR{"�y���`�N��B���f�
���I×|#�u������`5��C"�������z�3�=U��6U�
�I�=H�B�
��k��9
p����&�^q�bR�M��-.���J����Q(����"�<\���c6e$	�4d�h/%$ƈ��ʅz^[��b'��O����67��'z���Ƌm/R����K��俫)!w֕� :�R	݇lTnr��uק]>3���2�	�t��G�i?f5]M�������(����m�'��=W�RN9I��g��h��N(���8������a�!�`~t��$�Uv��50e(ե�e�q>I>b�yuF b���_x#���8Ο5�[��-ٽ�5j^W�E;(*iDZ-���h-�݆ub2�3tf3]�[#D�n}!2�H�V�E�sDE��|^���^��k��$�N�L�Y.m�\+�!:��[���"D%(��+X��HC~O���h�p1>��J��0D�TE�i�f
�+N}����s�K��uyl�{0U�0�-�H�T��m�O�<)�k&?��0g�ˈ����[��=�ʈb�Q�j~��Jx�ښ�X���4
�q�@�2~��&�z�o�%C����zY��p�t��� c���
۝ �SL(��(n��c1.�]�_5䶑49�B@�g��%I��sQi��7v}_J���=�Ktα"9����zGUF�q�Ǡ���O�����5)�g~��&!�82 c��Ā*���D1A�
��R��s���Ts�f�s�{Zr��Ϭ[@�(j� 2Ё^a��9����mu�g�^�S����J�9��
�F��Y.YS�h������xc7��J��}H��$^F���A"gvA��M+�Ŋ%
ʚaF��+s��K�t��]�8���4xʵGq?|��� �uC�~E�6�v��!ZV�����n�AUrH�*���rDRO�:.�|G�(X�4k�3³{��ڤcX��0����g�ASO��
�CV z~Ļ� ��}�1~ޔXKd �|�,%���ˠpW�C�M_�8���&����)�$�g���UB�b4$��jE_�����{���l�w)6�C:S�B�}�.5�S����d�K�c��}��V��6+\]Q+`��p�n�)�_�,�d�S'R4�T�6]sC#�Vb��&���/Zl�!�4* ���F�@9$�,뛪P�mwc��}��3yS���ou����m+d�������������ӿ���_z�BS��${L���䘘c{�+�Ľ�:��\��y�:�sy�j�s�r3%x4��d�U��T4�d{g�6�'�az:�{ߥ �����W'��������	���0v4LF�V�'S�Tax���;��&i����Q�;_��}Oh� ���C:��Y�n-	� P?�D5��]M��[~��&kK�4��ί"����~�����s䴜�tZ��0�6U_��w>��N�X�`���� �� y64詄$��Behq6������l_6B� ��U��ҮF�6�64�m���0��qK2C 6���Bdم/�~A���7.���y���:� �A���"amK���P�}>�	9�6��4��K������G_y��5���Yr��&酇=N���7�\�.���*��$��27�*Z�~�c5��L���>�G��KUd�8�tsi���f�ٌ�ل|�1D�?��uڧ�{#cw���yV�(�ڠ�ƛ-����p�'���@M�����SQͻЛ:@6B2@ �s��C��Ú�Bk2��SMHޫ#N� ��5G[_�J����z���� �:�U�|t���U�-�b�.2�5������ۏ��[���z`Za d>�Z���b��u`�4|,�/M5����f�Q��,�����\p8vSKiE��u��B�[���4{�#�A����«ʃC�x�BF�syo�i�C��'4�)^�7�+Eicv���EAB����߳F���Q���I��ׇ�6
j�l�s��M��b����״v-
G�(]�gJ�780'N���=�I���&���_�����o��* �B��O+���̈)X��B��,��1�m�z	I���H�jo����� x3�-�2o����^m�:�5�뛷�H������3�67�يU���|���yj>�wS�7�o�}7G���;{tx!z�t]h�a=0��oL���H_�t,���,:7��xHXH:,99�<-��l���x��, .Tr�����y�U	�HvkW�=��=�-SG�Tn��`o�PP��Ĳaľ�c���b�i���50� ��m�juL F(��a�ϧ m�1���J��@Z��F��	AX%ް搎��t�绩Aq���ajշr;Hrbn#H�	�s�K%k�r���b�D*6�3î���|��9�J=��>�K��Lv��/(D!��2�0���N%z�{�f��
����p|��!�*����.[E-;IX8��p��	������+�u	�Nk덷�������$��	q��Y�P㖨(J�n+Z2:����Ϝ����!��좠K1�w� rFa�az��<փ��G�s�^�҉��&�"�Mk(�)K�:֩�ŀ{ae�{*&z��l�~���t0QT�=K)ܢt�W�u��lۤRpJ�e�'���Ϟᤚ${}���ˈ	,m�ӓސ�O5`��G�Z4u�l��
�Z��E\��V(-;O�ĵ�sà4J�,��x Th�~r�*I2���ƫN�NEйl~�b�n���U�hiQZ�KLF��Bb��Z�/Q���s�D�x)t2��t��#$�KO&tm�ބ��'�la�>|�-��O(������a�����%���za�_��7�Gv��f�K}�L��印}A6���ze���}�[��(�۳�1)�g��sFʍ�͌DH{`0B(���4}9y������
��\Oٰ���{8��i�<ǳ��DMo���:e�Rut��h��OPO �r8꼄��F�7��e*OJ�m���j�ͳ9z^.�
x$�&X@�
U�ފ9��<�N�����_m&��X�:C�)PI@$1^\4U��7���N�����zuʣ!�{M7��nF7ݭ��M�|i�	:ڶ��˥��b������S6^]EŌ�.���&)��{A�i����P�<B���;�F�&���j=0� �l���;��vs������BАaԜ�)���$ܼ�<:v�k|m��&�6��7ŧ�y��~��F�o�2�:>�M�
5:q��$/��d�[o�M��z���i�ܥ�-�S�7B�1:��32Gu�`v;m^V��D��Ɲ���c���b��Aљ�}���5^�*��50�?��&�\���fJ�`"**�4��$�gSK�����������2�<Dmuǳ��z��+|J�s�ꋈ�_|Ri>8��XCnK����z��Q����ߧVR���i����'��¸����kW)�"��o��4�h	��|䁛.g|h��N�x��IZ����>,�7�m9�vB;�~��hם�?���-Mx:%��|a�,�N]Z4g� ㍥W,��[`B��6��W��˕�V1��@�0 �������3�`�yF�JUq4/0P45O�$=�U��B�pg2YF�t�
s�1����	.#����I��(劼�
r�;���5/؁|h����9:��n���U�`kD?�x&��i���S�E@��s&Ns���V ��Pr����>'�	���2���̄j�Q��bsy[n�LUl��}����`y�(D�'�PK����2����_�
%ed�����E�"�q�Pím�as.é6�-q~o�������a�DN��w|�훝�Ŕ���q���h���7��I�՘F�*HS��z9X�<��n(x�q��l?ږ4�
`'���������]�D߿%��v��Ŧ[1�<��N�o����W�Da�dX
��b�6�a��<RO �_S�(AT2m.�m-��%K�ߖ������y0M�6�ѻ4\T*79)8S1��P�����!8d{�ad1���u|����ABY�z�*>*Y�Ю�WQ	�Ol6)��� V�%a�N츫+�YĽ��{���կ:��&V���^O��MQ����e�V"XO��?�p"yM�h�G)��_d�ǘs�`9{�j��p̪� G[�Dn��R��Rӓ�=����tto�m/)z�B���5L
$�tцۀ��M��5biW���t���G���=��ڵEg_��.�EV���ur$1������Xѳ�x~P%5�@��k�� )KtI>Ϩ���v�M%@�q��U�MRa���U��F�3�iv�]�v��I ��ORw��h�jn��:��e�Að��̸d�ݔ�z��������o���X�K���\8a+ߴ���Bz�e9���W�[U���x4}涕�n$�e:_lx����Q��K9�)p̷xd|�B���|Dohh�,9�����#������#���^��*��=>�^.vU�̡P���s/֛3��%U�ڝ���d�8W���;��`����lϘ6�^l_L]! q����pG��T7��踾D2w�µ�@��ߐXa;�$���J�L�J�FW���t1[r���IS^�s:�!�{����M������E�P�b]�'7�l�8B��x\L��f�4c�w�06ӎWb��@�<�w���vvl�������RV�zg6��h��G����v��).���=���-��^�ݨ?��˵H�p@]��'YDf�p ��˵9��:w�3�[�@����&�憹��mQ�B���i���z�U��92Ȭ1)��|�\��d3n��o���?m���~�R�x4�cH��y�d4�N��J�����̲�qP�9hrQ��W�T��Ki���m��ͦQ�|�t�۶���}f���gs���^"2M�(f-��Bo��d���y�f���k�ُ�8U,L*�ɛT����,��C�:�q�?���`M&r�y�]�V���gqk�{�����&���2���N}�6*�����J߾�7�NoA�`_�<��q.��D瑁=܇�r2�]0���R�ys�˪������X��!֮�m��ϋ�2�ui�"'��H��tU���w��B���:�qT�o��ngVJ �9�A������ڮ���D��?�]v�{��A��|U��Kd�!�{���M|��탃B�����W�N36�5쏌��q�X�q����0�/3��j���h��]"�<ylЊW�U���}��i6��n�ƋDL��ϻ�n���\��$�~�8�7�7�f �����4�Ԗϲ)1z�/��ѧ�b�!�x��#���h����� �*�x6.�z�8�|�52�򡈴�<Rv`�~��k��y�H��D�L��dO��6�:�1 YST2��o�+��㛁� ��0�ݱ�I�Ԉse#��|Yܸ�I��O}� �,?Ɂ�~��k��T�-�$��劂� v�r�Î�[�ڮ����@gNb��{��M����n����<L�<$�;�I��Yb�e����\
 �i�^�)�3�N^w�b�%�=����{��Vy���ü��sá�����L}+u��Q����^��Zt�1��و���XLᲯ��˰�B4�&]�,��)��W�ͩWy��UB�U��M�0H/����g	��Oa7r!��IukJ� �х7<�Iy��?���rA��� �ZM��k������99)焬#<'��NF���^w�Y�b���揲��on41*a���Y�Z[���[;�7a�!kWڣ�g��s�C$�'���R��a�H$/�r�ΓD�k��K�b}dA|�7�n�Q�m�u3��;<�HVt��$�j��NU��(C/�Mʬ�Abqv*�t9�$�Y$�"uBS���p������U�h�WylzȐY�*`C�/��@��zV�� ,��Q|]���L9X�ǍF�$���"�80t�qmnz���1K��ZC�k�xB���6������#�o��{j84k ��3s��M*�zr&K���#�!Q�����f`�{�7���H�y�/;8H+A!�]�
�vF�h�op`�Ƃr���������9H�-�Ȋ�Y4h�(Y�ù���n"����2c2�:8��g6iŕ���=�b�,��=��<��
�_�XD7�/�����|̯���7)2��(�N+���0�~W/��wg0�'��fm]Mf��Ʀ�0���F{�ʐ�.@��� klHS���Qp:��ɱC\恍�	 N�V=��Ja�+)M-&&�^�@�ɓ�!A�uѓܘ�����NB1��ْI�%�&E�V�a�l����E޳U|�TK�M�`aZI��L}�b�Huh
��Fun֨&'R�Q�;Q����K���{�M�b�&��qp6�ƔM	��uR͸�L��N���zT��mtj��ڈOm@&)1��� %blao�BkIA��c�BC�r���{�z�f�&����۲�� ��U��]_��_�L�֙n�����![5@!��U����Г�wݤf?<�,Lu��Oj\Cв�p+�����U���Ḃ��͗��u�R=�x��o��OU*>�B�\)ܻ8<�b[|MĤ����L	뤈t>犒9�X������F��ʯĨ7�8��G��G(��õ�Sq����f��`.k���b�	�*�,�x��<9h�aH�D���]Mq�ʙ�~��';R`��O�|�;���ӌ&�6]��p�|,�œ|I0�M�4RI񁳧Xf[�/b�잁߲"��p��z2�����nI͡1R�}Ǵ�F�k���)D2`��CTփ�x� ��׃�tΛ�
߼w>�⬤A0���J�����ou�V��9g�����f
D��[.P8V5VH��ź���]hp�\G��t����^|��ą��7�����S������^�M�U��?�${���ܪ2�D�9wR����C�:'��z���ƣ`Hy���9)�H�˦!Lbn�j��jѳ �L��̨&��(r������,C�k�5��? k��Y>�~9|*Y[��Y�?}�����h�-�����܊���p����[�ȗk�����B��g�/���H �<�A�G����^c��Uȑ�E��r~�2�5�+��>������c��1Lp�Jٝ�EN�͛�BӂP���r��$�{!����^�}�i~����CO�&r����f윏����7�{�i�W����V~�$2��+��Jt#�0���M��'&PR��������B�����$3��V���{j]�g�"�Q�UGy�lݦ �k҂�����|@�s�3���R!.#���l~���4��]��M�;�W������}�;�>�^S�yֽ</>U�9��f����w�"����)��9�{5e�@�)%jz��&�y�씋v���Ec�d��:�QĞ���ȡK�G�{����#��J�y�~���d&��2>�s��w��I�����g\�&�K��4C9�B�&� Fu���턾(��飛/���;��9�%Ů56��k\M~'i�MO��~mK�4��i>����}:��hy_�X��S�����=$݀s��C)����H8��������;��_��q�uw�{8&��c,���5���Nu\kw�hF����OE�	z�Zz���y%Q;�*�R~��'�MG�}���~ꊙ�k��VVR1���z.�C�V��$��Wn�K�s�	��|� ŰМֻ4�����Q���nĥ�9��I�j�dz_;}nG$��5-V�ɅU��sIY(n��oQ��Q��;�K� �S�v�e�u��@+&n��*�"a�<��w7�r�Ah��+�	xcb�J+��_nf���*;�G۶�H������3�˂
$���
8
�F
h����^Of��F��0��~�'�ژ������3Eh����ȀW�@���"b����mc�FG�?��{�S����y�M��ʣ�����-�D2�x�'� �� 佴E���LvȾ�5t؜+Y~�VE��I]����%�fL���k�%z'�lm2��Ӯ1d��b���-.)7�&gu#x�d��=�J���~�2#Rt�i��,Π&����%e(f�׎�����OZ�R�4��D�o��E�:H��oo�+S�h��]��H�B�ǿt���l�ʝ���<M"m�?�U7x����<�?k�SR{�ts��x�V�Wyb˴*-5�p���Pi{�z����=[�������r�q&<�
�x>�1��A��Ƀ�Y��̩1��A,碮(B�z؈3B��T���?������1�`�c��f���={A���"y�3��c�t0I����x����H���E��\u	�`�R���(V���JjM��	�*���~O������V<��F���49)�7��]���~9�����,��8��M]�z�X�tT���6��� ^w���	�r��wXv��Û��Π���eH�}��L��ن�@ê^P�f�<D½ޝ��pB�t�F9o��x���bqQ�Z��i�;��R*d�H��[|�8������wN=���[�Љ�	,/����5�憥yoll�|�ORr�t ֈ�_�����h���W�pC���))p {��eL8�����C"��#�����T骚��7�4��9K�Nб�DF<U\�� ������*�np�����^h���@������3f����O�N��I�p���(E�I�+�$�)��H�c5�~{�!S�/�i�wiG�0ie��;�<�G7[jO*c��H9c��=�e
�z��1�� �|���+WU/^0(������\��o�!{kTar�Q�\#|����{�/ܓ�+?��>̳�;j+�l�멝���,v\�
�X�T�����~�xo6�{
F
����v�U�t�ocjU�K�&�\V|WpK�Q�?4|1�8ևw��6���J��n�˨� ���*�qA�w;5��F��Va��S�bil<���q�f1����QK�(r��ؗ�!�ϊ̃���צ��!l�:Z:�O�.�r!~R;L�n�u���������%������}>����	KJ���_T?��+�!���e0bر� yO�	�k��6��n��-��'�\����`Z�l"��6ƣ��.���n"�j��]GT"';b�P�In�|GV��Kˌ^A#"��E!Q_���+���o�\�/�J+򕽡.A��p����� �:߀����s�1H�c� ������b(P�W)����	qE"�LtYt:�%���L��C�7f�㝭i����ep',N�>L)"h����1B��)(�����ܰ�s�s�S;�k9�%�����zqn���(�)�oCh��3�*�����wEZ@�Y���6k='�_�!�v�i~K�dH���@,�DZ?�ؙ @���Vߧ���*7k0��9흱M��jYu�=6'�1>g>��
-`�z�T�I{ӛy�)�luD�R�3=\����w��ze��V�����9���z�q��h�ج�Uma�ۭ �a{�w�;a4%N�W��`�M	��Dv�;T��
�qE�"���H	v-/W����̬��9�	g�:n��o1eG����@u�ث�}���on���V$��f9�(_��������o�E�!:ڜ���8�Uי�Ԣn�1�P"b��Aa����Ц�����׋���ldJ!��n�����L�
]�K��VR��I��Kbz��跄3-�'�o��-����Y��U��(�΋UuJ��џy-9��7���I�.��-�M�7$��R�Z,�����6x�/$�O
֤g�\�0y ��YC.�>�]?~�'�u{�#���.0��Dv\׷�g\e�v��5����O���{@��Ub������=0Ru���Gq�W����k�@g���U�o�a���s�?1�� �q�_�y��dG0�2%8�*|E�ݹMf���҂Ώ1�q�����@i�9�l��$*k�ȕx���<?�N �Q��0�
iQ?u�t:" ��w����I��M0�
���{��b����x&�do�k�O�϶H�4��w� z�Ț���M�H2��.I�9�Z,�ǣ2����Z�B�!a�G�~O�����sezxd�Ŕ�辊���L�nT��c��n>�,|�*�V�8�c�<�n���&��ʾ�U�LZA��0\xꕻ��;y�`�d|���ԭ�}���2�B*8CwB>-H)�W#�9m��h%����e�6�g��q���|V�N?�~��KaqJ賃�I�ː��;�$!��&Xg��gL>!>��s (���
؄��H9'�?��b�ɤ�X^���kXD��y�I	e��߀������s���$q�ָ�a^�\ی��EˉRW�DSnL��5����B��q~�ù���@_j�1f"�T*?��I���w>xv���Fi�[���/+�C���Pi1λ �-O@�7	O7B�3_K8�.6��`�E"�AZ��X�3�.��0�f�C�A�����N��\��'u��;��cA�o(h���`�{_�.�mm���un����]?9�L=�WLwٯ�DX��'�R7�G��@*N�]�.�njD��U�fA�(�]��%oC쭦��}j�~��w��q�3�^��z/��ۜ��ombZ�
xV�<�bs��f*]����� ����1����!F�����wbu�y�`��J�x=����$5��@�Y+���6kߡr�5����5dl������Ӧ�6��t�Lo̎�x�鸊c{��.P�)+��2�)J
��ܬ�gg,��?���9h���q���H��y�{�U����q|�z�[�W�c����Q6H��[3�?1Q�6�#q�<�iD��~;P5�H�;�C�Jq.i�y೯m��۸^A75�R7ԕea���/��|$�Γ7�S_�Ur�����Q�.�=����sK �×<j��+�2�_����E0d?�(�J���}zN�^�C܆E�ޅ�_8�+@H��p��+��k�q�?��aY�+�ox����گ�{5Nk�fLo2��>�(�)�1�;��0R����E����IED�J�F�l4a<a������G���v����:��:�T	=���R��$��\U�as��ؾx�M� �[���2씊����CG��^����"֎��*V`u��KZ���cs.�,A���3U�������ޘ���tc>�]`n������I��b�ٱZỉ����v��c��-:�D���&����-+tW5�PYyV���:��Z���.��I���'�&��?dS����M a�[�-P1mq�UȊ
��e��JF�{鏴�R r����Z��=C����X��f�.U�,2�6 ?��tJ��v��2�4e�&�ký����\%�L�
���y�&}-�5�`Δ#s71�^���Dq��1�a~~Ј��.�ͷ�����Տl��3�fH똻��L5^��=�>o�n����_g���K�^��S1�RZG�SY�BP.r�t�r�@���9׀�G�<K��t�	O댠�VHYJI�\��Α���s(��ԣ�|1�ʵ�pBÒB�Po�b-!�~��O�!�����vk�!�D����C(_J�wȑ��h� ?�#vB@�r��k�Q$p��+��
**ZB�����	2B|G�t;~>�_�b�]��ʏ�x��+��C,������s�6F&96��԰f_W������[:��R*�8x��U�;
`�e�e�	���4��M�9�M���z�ێE�=ג�8��y�6#n��Tn��{���h��4'�,%�����h;��H��W=�J���̠ܽ��W�tZ���
��s`���$�˼��>o�-�i҃#�b�	b�-)A�oP$#�v�.5<�y>��P���yC����]���Am}�d�g;�yO;F�� $���٢.H�x������\�^98�&�FQj�k=j�]�a5T3��r��3ڑ�`)�52Pȴ=#2�zB��gw�Uu�!P�]�W�U޲Je)�Ԫ�����x���,G^ �1Iৰ+����C�V]���U��߶�=;}��U�C )��HX̯�Ģ{�2��H�4τ�?nF1�_��X����g�?|r�ٛ)�nd��o#���(�!�ӹi�R]�9@M�6�=�O�NL����S���u��F���S4P�3����i���_����k_cwi�Æ���F��8)��G�=�6@����XJ���1����n	D�Tf���-(	Jp�͐$ù�2jj�7��|� � ��_*+l��SZ�ik���Ԟ��-��]�m��Tnoc��_��}Mx���_�~p4�E�~�W��O��t;�F{��en3�+������Hm�=�v��hyC��(��č��������P�D��6&0��^]Y���}�,F�$~����F��a�A ����Z�g�"�Uͪ�&�|,I:�
-�RT|�+lxM9�ִ�-�v]��-/��Ғ�mV6[���q���*�l�������� ��A�9��[\�=�7��� A.��a�)��`�;����V�����)�s}�j�X�B�j��T��m(�X��;oL���4	%���S�|�Z:�!L5=����7<�Q=��93�����(4ꛒ�~�y:| 'Aɵ��H��	�X>��t)�2DW-ˬ.�����۟R�7r4���*1<p8Jk�E"H���P%�0'�r97 ^S�c{Soc��'�:��2���|�ix����+�N2K��Н��r9owY���dS$����)h���3�^����MpK�[Zc_�ų�2�D̙Q���x0kj���3V$����o��S��s~���i���ہ�X������?,69D�Tu��|�0IWg�҅"�S����q��S,Ƚ`����ɾ5����՞�`@}�ą���ۭ�`�!wY�&P�U\�G_銭Q<	�t@N�/��o����g��|ۛbs��+��;f�j���}�;{��̞���G����,�+o�wS&:���I��d&�¡�l�� �8��E���g
��U�i�Hw�B��i�B����Ԋ
���A{wUc�ɳ��vo�\*=o�1J#�IE�Y���'8��F��N��0_�r;KeAR����(��^K?�ku�H�^ C�Q�l(��n��!gj9�9��P��/���Z��6���j>�eT�#8-��76�몍FK������@>�z���	V����"��3@>nߋe�^�A��"� ֝}����^�5�k�l8,��^d�)X�v�j�P'�1w�S��e/�����	��4��{TM��2�����%����Z�������!�t�u�+�g�r��Y)V�� �P�w$�(z��B����<+�g�K
lEB������ٍ\��t|�,�\����X�v�BLS���%(`���
P��l���.W��݄>ey�um+��k���(��^��7Qc�5i	T�t�?n�y����ᦦ�,t���Y!+���_����7݊�u�U��H$�Ì�j�q�d.^�`��5�|]���q&�KB�ں�Z�a�����D�q�Y��,��@Z���_�RF!�
��17��E����)�W��/�/�@�=�\ܭ��). ظǆn<�=��~�����%,��	�Ԋ�紹��2�54��IZ0������tvs$�DI�ۯ���i�����&�u�1����%~�>%D8a %��4J\� ��2�]���G0o;�J4����N �#�l���{����>B���=��EЄ/}/��K��y�������;�V�R����ԭ�gK�1�liY1�X�;D�f�����5��'"���*�?0�]�<�:����`6�%yf8��P�(j�Qv\j���\�����*����?;���­�����zI^QEf�$1`��I�{:׬o�g����ɍ��T�����kN7@��p���S��Ɋ�O�>�h�s�05
�dg�~:��B(;@B���H��'2��b[58X��k}uqW)�9��_�U<D�<)��|��Z���LB������5Lp܆��?���x�e����u-�"�Zv�e�I���0���ȓE\�����уul��
T.U�ʵ�B��L`8{:�_��wҹd�3<;0B�m����׀9��怼b�� ]%�e�p�_n/�]�+~���J8CO �?��z�+ء��B�4�|Nb�IāGE����&�A�����XBS�y��S�ws�m��m{L�L���MY�X3�̮lM��=����e����%(ƌ��
�@>�����<�7�S!Ϗ���뱵���;&ѣ6����T]����m�e\+nd/�7Bt�)
l!�̓�jX�g�ĉ���vs�QʺA��re>�F�*���Qnq�b� ]��p<��z\1�h��S�Q�������c��]�8��D�he6�T�������ǤH k�~H)��{@ɧJ�8<��8,ywKt���SD�p >���~4�zmB!�Xzak;zy
�N��Vsf"ݒ�&��G�t_[�5�3�47�4�a�+��ɻ�;��I�O7K�y/#�h��z�&1;�����"�h%�����tDu��.{i6�9�]vy�rǧ2�
�0�f`Ӗ"
\6��凝���y8�|�w��Aei�5v?F��v����ll��p�Lt?�"B��Њ,�'O������������3y(d946�ے>j\ذb@`4�>�/ �?b�pk�A�@L����It)�����svn�L��e$���,��+}�=�r�#��!��}U�@���`>��:��z�I$�0:p��g#�l�,�>��:���L�sY�(��>�Ǽ'��m�>�D����s����cN9�5^QUVȪ�d�pb+e�p��Ց�[l�9��˵��_����^��Fx�G�V#x|�lIY$5�A�n�W�����f�+�_b���KD����m�`�P�]CT�| � n���r�*�p�&�Ͻ��v��.�7,��4���U�^���ќ��K�;�lRz�?_8�F~�A��eږ-0R�����g�-���Ar�
��D��Ui5q����yMˮ	�3��I��4C������rȍd3\�DuI^,<J:,��3Ѽ���~U��O������\�5)S��*C�~~�w���)�op�@�-�K�� %�3�Y���Q��C�Z�#R�u]�6g/�L���$��=K���/��F��	�x�M3C��8�A���@� �"S���K�Ro����j����qw��BN�DXS�k+^?O.2I9&��!�)xD�s�Qx�x��P�'��z�Gk��v���/$7�\��.W�Z6�v���<�3� ��[���G7V���:���E��LB;	�4.�>�n���$���A؝$DyE��1�U_����?�ȭ,�,�O�0@Q��@���c�*f�qz1�W�}����㾩TP��h�ٙyd�>��I�p�my���0�vsB;�7�/o'������U�
M�$��Z��J��H�����xK����I�ۖ��w���z�qLD���}M`�Bͷ��%�@m��(_���˵�.�6E�IX�W�F�Nݭ٨=Z��\�EW*
���U��Q�q�S�r���f/\̆�\����}�g x���^T�������12��E�/|(<6m��f�&Ϋ�fv�  ZS�F"}x'�b559��@1�Uװo��UT��A��?Q����ߙ�]+ǫv>A)Y����^'���0����-���h%�V�~�O3$10Dlؙ����mz����A!�l.�H��)����Qj_l2�	�m�|�,閒��'��&�q;o�lr�t��\��\�"K���*ܒ��y��*⍩$ �s���xƶ��|���1�JxӸ���"�������ZbKL+�1H��끂�j7;��⭮YrV�d0?)쮲0}TShr�vcq
W �,�W���)l��jc'������#-��e�Ͼh���_ 
Fi�B���y�)�A_�ƭ �R�b�W��������5����w3�%��V���ҩME �É��/x`� F����L`�|L�P�<���RfM�|~���_�y����)I����?!����!���:�I�����ۻ��9���M7�F��P\;-�@`��IP�@���#�m%#�(��x�$�г
x��R=c@��8h���0�4U�ؕ]��si���IeTJ`I��֏P�Ր%���H�������p�]w<���T�of�6�.�a��;�I���m��쑰S�WF�/��D":1?u�^T	��-����V���Y3��y��t��4Ew4#�=9����`�j�N��`��eZ!�V�V6l,F�'�R:��INE_�b��5H:1Y��V�:&6NBY�>�h�
�c$���ʇ�#x���`
u���VA�]E��d��c��C��o���NN���e�?X�ȿm+"3��?K3�Fބ7�( �������5�R�hh�{��l�s�$5M�>99n,m`<J�%<n�}��V�GP[_�'���iP�Z9�ɱ�N?�L�
�U�a�,���]��:,
= �J��v���_3��>���sS��Z/>(���9��w�Ĭ�D/*@Eu)��L�qI^r�,(�7�$�6D���{�}�V�SXIh� �6����S�,�~?4,zx���`.�S�j����a�Kgr7<�y4+2
��ӎ��@�b�|��ex{:�ؑ���j���_�̎��l���7)BP��%�Á���f��ʟ,Q^@��P�A"y�嗊�-y�Ep>���	T�E��2���r.M������}_�V�9��A�̬d�-��*g���z&���K��h��~�>��>JwO�lފ������z���f�j{��vpA(<k�~���k���mv��C ψ�J�p��U/�i)8Έ���7+@��)o��"(��C�a�����9$c�ֆ/�5�V�1w3~9�n��7'����;�<�`�L���wq����.�q�T^��%@�}a��l��1mw��V�bv_�щ�/�]���~FQ�	��Je�X�S�&��T��:v*N�mml�~��雸�b6��[��ޛ��ᗮY����@�������ڔ��2	��e]���c+ ���z=j�Z�4��>��[I�B��D� �oP���i�L�״I-�@>.�3�g#Ua��Q72��JC<[�?�����p
���8krn��n��@�9F}����c��7�<я�PU?�[	VP�x��R�;�P� 9C�E�L�ǚ���F>��?���/E�0o�^�fbTg�溚�+C���Ԅ��ZM���;��Җ���Zj��{��b7���	 �a��Љ|�ɸt�|s����0�
����\o%K�09S���/�"\H��T���	��g`��#�� ����W�<��`�a�=,s�
kR��T�ם�s<�(v�}�����[x��c�8w�t���o�%
`� �U��p����)\�>�`�$+�v���:G��n��IӣQ*�hD5��:�~��*����X5s,�U����3���B(%�a� +��ɶB�
�"���/��h=s\~�5@��	�m+�+
D��ݎշ"ޢ���Rũav�q�`>�fT��W'�V�1�>�����D@�O)��y�mH�C9�ēS��f��^�>�5�]�혜-z���oy��|������+�5�������@<���0)�!BA�Eз$Fz���P{B\"	�Ղ���3�6<G��%��ՉK�Kd��ΡR��u��55I���KQ��K���ڕw���j�cm��ɱ��4�*R$ˋ��@׸CnGB����&��X�<��T�a\���; �"��{iW�<E�����*:V���0�RϿ4�����Q�n�LD�?{6,K1��܅��)�� #�%t�M���e���E9�l�Ԟn�_�3ݦ2�ɬ;�Y���� �bNwܦM��L8*Fª�Fc�u=~���&R`��5��L`׵	`�>{D�d��+l����2���n���X�^!��f}f��8��Ug��b�i�v���]+��� ��<�F�⡫[��Z��XG���(r��DPXt��,��oFz��BU�7���FO�3��1�wr ���w�����V��`Q�� ��X�TgL�pD���G=��P��s��T3�k��@�Q1�Pײ����0H��sT��fO �[C|��>(n'���cwS��J��"�5�Lň���	W=����C�o���yd4)3BM��O�[M����PTna��TTQ�$מ���k�n]���(u�{�;�Q���"�f���QQhLX$�9e�gfH��$��~F����_���x�ЬyOk��4�y�����;�����.|i�k�ݲh�@�d؇x�� q8;�8����V��F��nYwtzo���8�ڨ���������hY��J#5�E���i��;�{5�w��3r�l?�k�5����C�qr_�d`�����{ @�G���Y%��#��K��ߟ�^�'G+޲k짻ƫ�{O��Q�l`ћi�V��3Q`���?�;w iT4`�Ƶ�Ux=:�w#���sV�-��7T���j(ܹ���+Fh���E���m������՛#÷�ĞgG@�x;"�����o�NB��sNY�i-�Y�D2��݄y9<�V$�-X�W���$[,�FW��R��:������fD$?Ej����g�=�5,`Jg���֡Q���Y�{1N�e�M_š>��W�����q�te��,C/���-��=��l�'pTj���_��1
A�3_2�]�m��UX�@��`?���b������u�_Y�J<Z7�*T�S���[��)_�N�a��Tj��3*p-
3�����Pܥ�L��L���m���P=؟C�Ã5�)*UU�����M��I�/>�C/x�?���K`���n���/>��'��JU/����@�������@���f?D՟�j=�\r�|�9�C��fVi�1�,��"4�?��B�I����pr���qf�l�ő�rJ]�����	@J~���Y�:�<�M���"V��jk��i����]��h�����{���c�A"a��o�<+z�P��]��k֒�����^P_P�]�5�0<�ri�Y/��/A�Q�K����$��4��J��0�n��Գ�]R��v��}UƦ�8l��#_���}C�"��a�W�]�6Z���	��7� 8B��h��PXk%6Wv�K��r��g���I�I����5ډ:0F�f�U���c�2!�P��#�f1�SV�e��XQjn��D�����MG�[�4]�Q�9��քW��_K�)_N=��#��5���p�x�DkSy0gO�|��9_E^rw��XR!/�̒+
ߐ�Q�	I^��;~dͼ�� ���H���BnRPk�-�lڒ�fQԦ�B2}Ї�pYf�	wN�lD��o��n��
bQ(���f���yk�FfV��M�E��@��B��E~]ܨ�����v|��Y�b��45���(���Y�E�́<�w�����Xˉ.Zbp�����qچ͸PشS���(�,/�ۦ��Q�L����Q�j�E����C].;���M���`>���퓷���F�;��R��@���ǕPi:�2�8�g9�l�}��F��~U@<�AQ"���\��*.]ʘZT�.ۧ<�C�Kh>VN܁p]Y�c�+�(iw�1�d�N��������$�ͽ����]��8����p� &�O݋��4����ш�gn�b��Q���tp�!���%e����U�d�4����I�JE�>>9����@�[�#��{f��6O]�����Kx���ە���,����¿�H��	R����N�~�(=a��@��2�&����b*8�M����A�T�zn���H֖6�������f,�;�K�҆T)n�����pX����W��^}#9��t�.����h�Oèm��.jX/�֛<	y��������,]dt�/ᦟܞ|���ΰ�y,o���iT �|�RZ�ħ�Fx�
߉(�S��j�c[�����3�KfE!PRP���G�/���z_�ѹ+��]N5�|���(���*>�C�2�����l�I2�'M��ר*3�"��N+�V+z��ܭ���-�$���$��oAyT�Op� 3���(���_V�>�~��r�j�q>4���x�z]�G�,���*A�mu�S[����^I�6[�b������������L�W�i��i0����$X���c��^���9?�	�������T&u�}\"�$����{pX��	����o-��;eQ����̗������L�<�8�V���k�zM�J�)"h)iNi��E�9���vjˀE'Ё��U�:� ��ZK��3��Y$M�J���\b�ň4���p)3)>Sc\+&�n��<�zn]=�]���%����q�+kyP����HSd% $�\�Y�`��r<1��zǚ+����F��r�z��m���|(CJ�2(oZ�EhN�|�g.�m$�[�]��J��61]��1�
���i ��E54���5:&����2��P�i�F����gbKa�N��T��P��̎47c�����rQ�[�?p�7�l�&x#(Oe�L4��f�֒��мEb20��G�N�i�d]�˩����79���h.T�4�ܬ��Y��*mT��L}]���)]o������RB�(��������T�~0���A���"og�ҋV�������r�	Y��i�G�T5Vk���e�jM�B�I�~!�t�((w�,	���&Д��-x���_?��'�u=NLo�C�˽�5�xH\� �Y�.XWl&��M=O�o������1F�e::V� �6�#v���J����qy�*R�?�G����%%aA���W��Ag�\��H��h�xp�����}�\��d���-�e�_�+����yb��:*��.�C�Η�٫!A.��Ӡ�� �\/�������`��EKxf��hd�'��/�m��H���jj����ef��)�}�)()�ӷ좣P�uV%�D��+�=кJ۔j����GU�7�ls���(���q4��y��Ά�$�{�Y�4m?$�M�!�J��3�j%Nt.:1�o�}(�o@����͎݋��.�g/`1�[���8�� �,�}7�d�/�$gV ��KI��RhF��� �}f⼌ա?A_{	��d���[��n����gC��+7�`Oj���@�t�xW_*vY=|��m.�]���<��/�{yWq�|������U�688)1mȚI9gl���/#�H�H�C���e!�w$w�&��)M���Y�fĘ3�''����z���k�~�-V�R�%_�{���=5��5�DU��F���g�U�_��Mk9�v:g��&.Ҫ�n 3	��H�+��I�uft�!Hu��NM���ή�ԥ���?�z��L���'��θ��e�	��S�qѳ+k��Nȳ�Z_|8?�V1���O�7N	�W����ÿ�#1$G����@J�@I���zp��p?�L�m����E-��F	k��m�ΎgY���Mo���r3�d�m �>�
Ҷ�,d;�5)X,-�|H����0!�q�:���a����5\�ɕ/���մ�2i>3:DB�*���NJ2G���d�e�.b��m}�)?8׍�%��錬��J����F8�_�v���ۮI��C���*5BI�o���7q��g�il�חV�)�3��� a,Q��w��Ӆ�N�jęy�ڶ�Z���,�0OGT&�S�D�
$\'�0�@��}��Y.������
*��A3T�r�%#�]����b�����K<Faβ0F�
gA۷}�<�UCj��)%>H;�bw�,�]�$�l�Ր���#mE���z�既�o�˦�Miʧ4+M�'LT�Z��?Ϛ��N`��,+v�m����$�OVj��oR0	�'w�8?�$J����M	X=z8�2KD�I��y2����	.�uҲ�Ofp����)��6N�{8�*RrV�b���)S��{�����#�"(KL_A�id�|�$��tqr#�;�kP����W�� (�h0uQ-��FcK응	��8�)��ɢ�A`��\�r���W\}T0Ѽ� �~AT؈�9�u�uN��8���w&��:w����u�H�Y{� ����T�O���u6�A��[�2�>^�F���ݛ����Xq���j�I��/vݔn�W廸%	jw��!s @��5-xHNf��d����֓w����mT���v�*�ڈszS����y�*�}�����<����Y�k�Ʋ���oVYܾ󘙷�m�X���uY�7�U�p�T�:����	_�eʒ��y2#X(t�1&lgn�47���	Q���y�"K��{cͽ������!�9p�m�8=�:=���ě�����������TaJ��G�:�	�k8��7��,�f��C�X=�<�&���88�;��/~�'��(��x̣�%
 �
�r$Գ�_EV3�m�A��?o��4\Zֲ5��ώP�- �W�%�ߙ�x=kHC�g�YHA��˱
�uK��T��y�HN�jQ���0#�q�73��)�"���0�/Hy�g
����j�o� u�I���p��u}q=�89P�\b���&����(�	�|��õȎ�/��D1���2x�Oƕ2�)��U���5ս���MM���sWtB���&0��^�\��7ԫ��J%t�,7ז@�D3�:~WL&,���Q���lSg�wc�A�P1�U&��o���Q{�+&j6�.˻�K��L�����R���6�<(x5@E�}}�@�Mf�Sb�'4�H���W�4�Yɬau��.��`�̽���)\�I��Lځ�o͏E�l�B�X���7[ל�a!F{
7T�V7�U��.�Q���V�^W�l�i�����y��aP���紩Μ����!��}:'lzL��iY^�k�OGU6#�n�w�kJ\�X-���IH�
=r�_rĠ�**/��3���PP� =�]�}���'w�X#�� V�D���~���l��uaMY�
,ь����h��O'q]7����^a gcvE�ۇ�o�G�zⶒ��9�hC}�����T��o��B�M��;�I����
�k}��D�a�¨�`�R�zX�7S�֋V���.�k��)_����/x�uu���d�#,&����Z��̈́a�S��{[�!���g�`�1u�y���t
�������/y�Ū��0|0¹Z��Ai���^��~}���b�L�}�����G"�yq�^��E�o��U�`���t2}(�i���(�����)��:C{���.-`Y9$����|�m/�B$.i��K�b������j�;fT��Rm�P>������d������>����S�@`�~W�D�E�7��]X;o��� Z+�usO��6�v��W7Uv��X^ĝӀi/�'��E�Aܻ-�}zk5��_��&�9@C�$��������Z��W���.����vy�&NM��j�a���r_��I��Exb��;� V��}k�C�9��|��	�f�y�h���\DuQ�D�Ե��X����\fm�8q�1ڭb_�2�>�X�L΍�W��ۧ�X8� �bi&��D�h�֣�N_	�PP�BJ_�bQ�,(�7G���?���=@翇P�8\?����5��8�U���D��:[62�K�����	FrO<��!t,��m�2��kerQnB�`�Ff�0����;�:J�C��%t��C���ã���ӎX�����acoq�{�[��� ��(�LW�b������~��)��'`[G���ת���#vo�@[f�\Eu���i���G>�s����2c�O�W�Zl?a��2��Fv��;���#!z��q.%,���>:�bh���LU?�x^��T\N�]C@�b��8�r�b�>&D�MeJ�:�(���V�N=#���\Db�H=|/���MG`PV��7�?(n�Pe�܌�8=|�x�t�'\p����ʃ������s6��L�c�m�D�����x/�>�_��)�C�������WY܍X�I#Q�L�i �rxͫГV/U	��Y"�)�@9O	��?+���En����i8A���a�b�n�GZXn�.�$���л��	LC�$ �L�QX�t�����r�a.��	W�\���~�1 �@���"�`8I�"���2�#�������<W�pMҪ���¶�D� Y���c�zoj��ZyU����G�J!�������ʮZ S�k�`������+���Tݤ���|0SUte�(x��Vb�Z�{�Jes�o1�BQھ�N����]�|�՛���AP���ZQ���R��^�<	�k�7��������UK�@���>��n+�ND�hJ_�:G���M�o��n۩}~�c`7��?���Z�o��(;�%L��7��* �A�����]i���y�nܰ����c%;�GV6�y�n&���*E�q���<o~����2q�u���Zr�O��
��r�'�U��4�⋔r�E��/C? �}b׊m���.���/���9&�wl�!dv�ڊ=N�`~����4XhJe���S]�I?:'FH�e>Rt���+�z�Ө�5䮢����y�`?�G9�9�^r�\�9F������&r[ԡ9CU�߅@ջ�l ��u�r�_8 TEDg�qFκrN[x��9��~��n�>����t��ϺN �:�E�2#$���(�C�=��3.�Ֆ��B�%��Q?��	�7;�
/��}�ّ��%%�M��Rρ�za}��i�i�����G�,����5�Nʇ�ד��t��G�y�6_��*
0��N�`�^��^�?�)b��:�2��W����\�v��[;�Z	��-��`_�7���:<σ�q�j�1KA^���س��p%E�zp�.f"��R���ضj�ʦ W�m������s��^G�CB���n1��mõ�Yo��	m�R�cc��$,cwQ�@�{4}{��̖��� c="�_L�A	E��!�K�/f
�x�	��s�pqu�fѪ� ��-A��]��a��4��k�ym�>�WC��b�J�]�`3U�R*C�Ñ+�v�Py�ٓ�k��q�Mh'�((9OD��7�|��J��s�U���&ޞr(N2�ݸ���i��X�r�r��F�NT?�,���)V��d(z��0,ҫ5�!{k3b.�:l�z��� �"����5�v���C������\8���2�!,�����]yH����&�tfZ�P�r	Qfz䖵�o�6L%?=��������qV��@W�ӓ[�]K�Gp��k�X�L�?S$��R���D��(��n �)?ɵ°���U�]����aM�P%D欂1��l_#(���d}�r�ʤ�o��PO�T��a�&����!�!�$�Kd5J�=OK(:�M�:�?q�j�6�L!um^�G�с��X���}�R.nٍ�9||�b=SԴpR���qG�g�M�i
-/NU�tSQ���Á0�6�|�����Q���-0%��YyX���e�\1Z��mF/�4oh��l�s^Ռe���K�D�:����r%?:޸�"]d�}��5�?(�)x62��w���gS�1ʼ���,��.��b����	0Z�@$ş��?�h�,���|)���5APUU�����KgL��pnW����-��������Jh/ʗ�O!�%�$��ȭDyQxl�+eJ9{a�$��Y6�X�V�
�h�R�6iv
RrY��bnkS�$��z{��5��\����@����5��{RSR�]���U6s�p��Mr��J�`���_�i�����£��4N���0D�b=��P=����lVr��4�'�,ɜ�NXS�����)�3����.r-�q�K�ni�ll�t��]���Nnhb�@/՘�Z����� s[Q2���l�>�;sL�}��}��3e0>T����"�%Ȥ~`��z#։<���~M䷡o�m�n�h��A�G�$�[~.,�|�дg�d�̤�C�7�)�.����Oں�6'�FA}S��-g0X�Q"�B4>��&afݜ�R�:/{D഍����<p�����;�h��s�J^��!G�2�y\�.hT�>*S����6����l�n,��G!ŷ�������J�Nu����m����g2�'�g!f����8F�vC�� �BXy��j��q�q�E�5"*���!�NY|0�d&�o�������J��б������;���B��G��hL)�����3���;Fs��s�l�ڈ�FJ�%Ħ_\S�d��@��ǈ� ygo�b�D[���O�U����a�N(�$�Ù[�m��؀3�￝�z��ǡ,����'�n����gN�D抬R6���6b��g���[�'C|u���i�#��3���@��(��b%��4L/���]�	0f�^ű��#�0��������	?�K�k����4I�߶B߷���5�ˏ�RZ��P~�O��|��&�ٯ ���b`c&�~�PF������ �y�hsQ��23KyLP��v74q���o��ʀ��+�O�ӊ���wK����� 9��acƬ�z�@WU[ՠ:�g��4&K߱���S,�HTu�^ә�^���W�Ξ��r�yO�˺VQ7��(�h6<�T DN�d_�H�d]���)҆�1�Y�;�5�L��Ӣ�[�y+��Y���^6
�BZ{�G|0�S
X�I�
�8S�x_X�H���������+��x�-��5=��mgݿ �hf��	�������T`�~N��v�+�RWo?G�4��&J��0��C�X9�d�.ikbv���b�z�	iK��mz�Q��9����7�HG��X'=ҠA���[�v:U��߰��>���>��\�����8�N�s�
t�G��'Tk��%?#s��tK$�@��X�iQs�����NE�+e��������E�v�_1��E}��O��F���oX̭H��o���_���B'��S\��r?L�'{�6��~B��9_�ynj����W��Ѿ�g9�{{�Y��u.��hf�0�,�;:�ιLR4��RXU�������Xd�PD(R3����o����'�d���6���q,��Jcdi��=����aL��N���l՛};_�G�Ad�RGdק�Z��n8У�>���K�n���XC(��F��UR�-�Z9]xB�ƝǺXq6�̜�F��u:��Q��g��lW�f�wSYi/��h�v`�����j��Z�"��=a��P}���˼>B;{Ԕ@�_P8�,^-�jXu��TAܛ �P����y��1����t��$~9Y�A���f��!mBz��_w��%�4$�2k%�ǎ�7�qV�9��oB�x�b�d��I�̄��@�T��TJf���68�C
5~��^ ]n�&.# �����+e�Ş�lj7�\��'t2xM���Zx���{A�-q��Dx�zdI=�2�I��<!����)_T�o�X���h\�"�Y)�\��|�y�Jht��X�6�e76���b�67w(�Yyy>�G�HH��̋��dRak����#>I�j�x�;�,y���{;-��!xj�2�vd��w��g�vZ����BR��>m�G*�qю�O�#A1_��W��Y��񽉯��j �Z�3���&��f�����m�cv�ֺCF��	�m�����W1B���2�6D�x;��$a=����s��>��'��.Ú�)�RS��"�2��F�@��37��n��O�Xz=9+��^&MK4Zm�g)��_�TL(�t��8 yZ^c�-珙���
N�L<�c�WQH`m���>㤜���Ś�M =�<�"T�"?��-�4	f��)c��c��]{C�3+����Bh_�6r�[-�|}�^�z�׃;FnW��8�N�8��%�4��&��K�D�n�������}Kj��KN�k�����Qr���	�+y ~�_.�`� i�Oƣ��a���jR'�a�K�R#�1�X��~�׶���DK�����J��mXQ�߈�vet����fg�����ܸ��B������j1���*�J}��3-�f���Ua��ja�ҷ�<�D)6r ���r
�o�e
�A�we�p0�h��\� Uؙ'��8�j�.Z�5�G6\�^�>���&$J���6���}+i�+�CI2h��҃M�K��qg�H��X�X�����wa�	w��TF;q����ZX�F��/��FݹRq��0WO���1�p7������%X~�	���ːr6�%�-� �>fw�P����5}ş;&�O��������.K�T��ɀ$+6Ȗ	:��8��a�4ˋ�o�F�^Н�G ڢ�9\0FJ��w���>����J1u=c��)ݛ�އ��$ח�B%���棬z�'�K`�����Ѱ����=���plZ=K@������p�+֟� "'��8�1~�l�J�����!��x~�x�\���F����Ec͔��mt��G�(	��ǩ��5tD/{��HIsf�W�mЁR��lzf'sp�o�/Yk��vu�����{�} �����@�%vjMuU/���~�l�������d��X�n�d���u���,� [l�#3v�Kq���5�q|��_�����r�U�;{!���'�����i��ФK.�[�u0��lÕ���Z�ydb؋)�d˂�O����(h���P�@�B�8^|�հ4G^�kv2���0<�&�7ۮٸ��L@ۢ����A.��Dz�ɱ��	���Z-����Aa������� Nc2���(��ԯ���b�7�P9��m��z������>���9�ѣ��r5��%c��C��`�px'y#}nEa�'�m�I�l;1dS7"A�4�]:!�����G�Z�o�;��8��,�����'���x,$���A,=jI���j$[�
Diֻ1�;n>qRhh|�����Щ�ә��\��{D
�#<ś���=��W.%����%�e�dM'^��qLL�
;�ڀ2��_l5�ƛ[�V -i"p��T�n�v�"�MF�R�9?���(�+��|z]6��������WS�>��S�д��2��tm�S�ń!��T��nD���!PbS.�,��orFjO��?v���s85&֢/.�j�X�;�;���A�@4�����t���d��M؈\���)�ꎔK��E^<h�!W3� Iɦ��vܾ�;��"he�F�N�9�z/���b,=vK(���pJJӤ�/�n�9jI�X9Y�� �u`f�c��dyRz�zM���/8��+J��(�ų!}@�
���=���>�k�b�tb^��Q^�p�s���a�h��ECD��`$��y�2�� ��ځ�����h�3���0|C����<[N�I�b�J�Tn�;&�O�b��	�8��CW�S@@h��~������'�,���}�
��_D���W�ͩ�דkUV+�yش|>����~��O����k:����ݛ�����l�6��^$�T���FM8�w�D���&��C=�y���R�� �R�&lzY�?�7lc�JV#����H�~A��$f����}()3�kv)3R��c�u���=M?;Qf�
���@��Qc�l����[�J��� %*b��/-����a�s�g;�3q<Y�P�W���CaiFEr�e]�'�fh�^r�Ju,����^(�ް�,'_f�:��M<��x4���-��W�^����1)v�Z���!�G�H(b�����{�I#QK��?ɾ(G�"���ج��Yy��ĕ��d�܅r����z�a�V�\Y&�n��a_�7�TV$:�d���@����ҋ==oB���E�������K���-��$����kim`[�\}{<��n��,�ZRW���L�b��d�}.�B���m�u&��S��wX�h��TjT'�=n���2�՟m�G�V~���8��?�w���J���pp�"���Z#L���.���P$\�p���]9�(TF��CS�9��9a��-��7T������oM�X�+��"�r�x���1���!�x��H�}!ke6k!�rT���#��$q������|�	r��cv�C`����1���)P�d� �Te�925�f	oTD�H�&��3���������B�������j&Ǣ���hb�!4��t���U���*�6��T���R|�aA��?��� %vbc1���(8�Gn�*�k"��q�~h���_�@�:�I��ؐ�l��g��=I��e& �S�|�h�e����P��#�5�@��J
�F3a�H.���k���8i�T������D�ͼ�X��f���*��7G��� @��l�\�}��3�>���(qCv`�P$~�K�1R�����0;��n����PaNް�H���jBzJA�����Q���g�뗙k��C��<�#x"
����p�G�%�}��8�����]%^���sFI�)�$_��A�D������E�E�>�h��|��Ov�t��y��	i�����qο\��<������"����q�[N���o��ݙ]��ό]6$%�18��;\>�o����-��4 _c��v�l�n͎�gy��9��%��E�k.y�]����<��&O/�R���oF���^>�n$d�>��!(�L�;����ro��T)�^��ç%o�o�����gLLhLN���QD
L����,d�҇E��[��"��s�����i���tq�[�u%�����t��ꝑ�F"J����[������]H�����s'����$�\��[8�iJ=�"�P�9^)���v��<��i>3ޥ�=�{r·5 `���������A�j�F�:5FH9%���I��w���_(;��ྉ�<�{�a퓛|:@P��!�!�p3�K]�RN��c�z��F+eiaW�kK������_.4����x���� ��"HnU h���@d�m��U脨"42��k�B6QKY_����� iZ��՘ _�L/n1�m�+Uxε��x~�h�`m�#Y���j'��]�
���?-z�T���4��YpL#����f�����F��v �)2�R�.ȡ��3�mJ�U��!���of�5��+��l�aV8���=MS�BF�eG��	Q���_��klO��A?�;�T[Zh!�yd�b�1ͻY��9}E'y����u3e������I�F�n��:��(��z��Aܯd�+Q�����4� ��\w��7��̹��>���%D���3iy�P�ɥɻk����$	�;J�9r�&櫷��c�-�L��[��S�V���\���*PU?s6gW�^ۮ���a
��p �x��aO�",sh3�<�T#{��X󑻢߾;�I�!�;Υ,F���%b���֫��*�&ir�}�d���bSeo]��gq�k�`��?������Ru ����e�+v�i�ń!r#W$�Kw-���{~��/p�!ɥC�ڡ�k{��@ŝ	��K��Q�S����y��t���4�DiN��IH)� Y�U��t�.|s����9���
��ۊ��-��L9�)ŔL	A9!��K�(��)�x��0�1w1��'�K���:��4����"s����9@����%x
,Rȇ�Zy�\)=D�� zCBr*���8_߾
��G>���	3�A�x��%e �f�<�v�LDM�`��p���~��X�^AR+)]t�8&�'��E~%�u���"���"��S�����7�s�o'ѵ�@���L+;���y@�[���´�؎]�n��^�<\��,k�O?X���<ǣ��k�A�i��C�o7�aB��+n ����+�NIa�#�\�����e��i��T�eJ��h@n�U�XU�+̵�G�l�ؓ1�q�2C������8��y�ۣ�ޞ6Y{|=5���<�E�+* ��CV�`�(�dQV(��(ָ��D�l�_���l��us�R��VQkN+V��`W����Nɣ�>b������HoP�D8�|�7��	7WO�Η�L��ls�K"ZR5B�j�������OwO����i�Ү�ؘ��]']�P��J=���PE_�n6�G.��]�-Q� �y����ߊ��Je I	��`��i-�H.���УN+c��$��8��V��q��蟻s"y�Uv��/��&�?챮�w����Ü�~%.�gKw��K��^�Dz�a"���
��u$ԝHl�Jc
�)T���ȲF�
�
��FĽ#i��*�ȸ���_�{W��h��/I�\m<���b�s��`��8p��B?\d�W+���۲��`�Cjum^cF6h�6_L.��u��|��= �:����[g�q����{4EA!h�D=�ь�1�\x�k�A����H���
X&@H�=�����%j�z�(�޼b�<���|pV��v�%��^i�3���`sq��Rq(1.9P�V�	�#N�>�-27�OH��[��p���sI�0L|�<F�Թ��5=����:�L�B�7�	����.��,��i.t�Үw�?k<N�5D�6Ã(vz���n^��=D*|�r���-%� L�{��9���~B��3�4feԪu\v-cU��ŏG{����ZZQEZ��f&��О�A���2d�O�y©���L����<1�3ջ��*�:~9D�="��[�[l�]~vG��G��pI�3��ۇ<�`;&u-mj+�j���ӓ?MKI?�Di���^�S���U3f�-^��^��!޹��8҇�B�8L�~,��%�D��(-�S�m*я-��Q�W�z�=�0mՀ��10Zx�+�JP��I����)T�����`fo���Y>��Bhz�'\`�3����@�]����vx�R_;9������#���Ԓ�E�3�K�	�↸�cS��gi���Zda���5et��?`��_|늉,k�Cw��G�50�'j�>���%�ӭu�[�:�V+�����@��=L_����|�,(rg[;q�=����qɘ�+��Ƶ��ٽi��/[�	�X����f��Kv��i��N��
�E%xW&sE⳧v��+�E�[]��msA�,���k��;�zY\� �33�D�?��# ��6)[�Ě%m�
��u)e��Xi�;�:�p<���9��g�^�(��ޏ�h>��l�4@���e,�ƥL�;L�-r�",(���L�"u����ϲ�	^"AX,�3) ���Q���}W�ݹ	�4mxm���sp�?x��h�x!����`�ʁs��T�_wY�8"x�U�y�kG�1��X��|TDʏ�d�n�?��U>�5�Py��N�%j0.iK)��2S��
�X65�r��%?T�d,&�EP��꼗��s��D���b�#�L�V�mV7�c����ǁ��VH�5X�H�2�;�'s�Q�O�d�H�@	�d��#�n|��-K]q8���\�*�GMY�e[:fAC<�eJV@��ol�����4�q�%���̵���C �}W*^u���z�J��[��Nn�:x�u�J4��uRb���������:)ʎ2�G�nlb`�VhMDqg�D����}ߺlf���P-���)����x��*i�ej��+�6��٦�S:�5�(C�Dw�G�L5^i���"^��L�hQ76���W׋��DK��U/Nҕ��n��y���AO�O�6�De��M!�ߖ�`���~��Ċ�؂8�:k�]�'��(��
״�Qd�5&+n.B`���? m�p�Oaw�C8K���u�.�S�Ǟ��[¬�\��4K����&'���y�_(��N�{�9]�4��E\�k�"�$��6�����K�ƕ�V.�b�M��$��	Пq�5:�PJf|p����+���@�핕(m�:���� T��3ͼ���C�1:��o�NG	v���\N����r�j��T]"�n�jm@t�d�|��e(9p�}��A�4ƽ\�ЎFr���R�9���9��@d(O���R�H�*�K�M�4*-v/Sv��.cK���}�X����7Ty�,�q*gC,d��#ebd7� Վ��A8Þ�#+r��w�B?��k{�h�h��f�g�b�@�֘M��*;���)p
��V�y�4 �N!���î1��[�l=�7Oc��J��X������당�:F�8�})RPg&��K���ѣs�͛C�?}N�1�[\�ײ;���:%^$T%�/���a�"?��?sfɛ����A�b�D3A�A��ƻe���e�S@��#�`���(w���F���ȱ)�T^�� �'��d��d��f�]�ܬ*ǰ�}n׈��WN`�~��I�HixJ��I�H�HHd~��Lef�a��7�,���
,�.6�A�9T/��}D4�%k�7�8_.JS�����nm�q���Ƙ���uQ	x�eX4R<?�䜺��m���xӏ�1���\�s?a�9�TJ�,�]��QJ�٤��W�6��z'���l��wl�~���C؆)PZq�[Ÿ�W#�ξ�
đ,�b�8�ۮ A���B��71��Yt�ԕ�ݱ"G�{����
)�6�'F�u�w�,��:�sAe�>ꥹ]��<�v���U��df�h
���!z��c޳-ag���Z�D��P1��@�d�ޘ5��C���Zv��˼)Wxk���hdǊs.X����|�P�!��X/�B7i|:1m�O����%����@úl`�d^2e��rU�{��y��O8�CXKW�F��8��
���v�|�!I����.yC~N��� ����n���f!��t|�ۥu�P�/�.�3I�,u��Ó󓲵jw�,���P!�����q����+�����MQ�����%�]�j�,]銄�ʯN��M^b�.��%\�x=�s�Z�xrf�a&]�5�,�J���� ���i�Ki�_�"�x�M�=i=W�40�������PV����ث��i�FAՔ]w�� $a�,�Ah�\!\=p�o�O��	��_����N�6��Q �k&���٩��W�Q~��um����;X,��G<i��<Ss��.N����{km��B%?Όձ/qo��E�FOI�<��?ц.t����/�6�"��H`,���m���]4���;hU'u�p?_��&~9�[bop�/��Q�f�eo�D�M���r|S�Z�}�".��Yg�n2��-R-_����®����n!5A��Jx��-� >F��W�:���nr�PqB��*�� pi�ܜmj]���Ƹ:e
,��1I��0`�_F����a!M���e�
ƹe	������[�g��_�L��`�e���9+�y;絋�2�PY�����,�ڤ���-�`�	&��fq��-���
����:q�U5�.N��9Ц��Y O:�x&˲��`�=X�����-S(L�X�!�QdX�
����2�"�m�գ(���/(�v��{�"�η�n��K�����ô���\�ɥ3�X́B�dģ�`�/��ʩ]�2A��2gw�J��#�k�c�x����$�슭��b�1I���+�Eܬ�i!�wּṷ��'��Of�9I�W6M�����L������ ���{����&<AtUHa��vQ�<#w�)v	4JeO�G��Ƚ@?���(������Ab�	�	��'����6�}<D(a�<��d�ˆ�Q�mԥ6�7h���!��[����aю�pDF�9!�Ⱦ{`��ו�JDb5��"I��Y1^j��E$���CcNj�E��6�N����P�''����)�Bn�'+�8E:`Z���c��/�S�k�ڐ��w/$A��VO�h[�9�/�H���$��p>����	8V;.tSZR$_�j�R@�`y��7߲7��0G�%ב ��Cv�eH=��F���9�֚RvUÇvy�{3����,��S���IE��屢�1��A~>\�.��W`�uL��`��з��򠕨���p��ܤ�i��b��	��9���g��<�Xg)���a\'5_�����
�>&�G,�O���H���I�&�-d�}�g��ıY��c���R�Af�tjo�vNRֈx���wM��������TaOf1�G�
f{`1� @]�>b�����DY�0NL��t@A�E	]8����7a��K��N�d�ы���scu�i�ɦn����􌯇���ɫi	{F�p	��,z�����.�$D'��O��%KZO�I��$�KR���&�74����N�N˄W�b4�;���Pw��P������lq��.��7����G]L����U��V�\�,��&��pVM�ޓU}Ҋ&mK�3_$w�2�a���H6�и�}�M8�� �R:5��ENt+:���'w��������{�;�5�_=q�=zo�����l\gGn)�"�j}�|*y�j�b���s�@G���3Xz�6iRG�x#w�&�o2��Sp�lF����M\.���� ��^�6�)t�22&������Cl��cRaZ�sM8���2t_��DL�k�*�]��oFA6�o(qq�
;�D���}��bG�Ft���P�U A`%�t�h��;��=�EN5np,�%�\V���%�K�*���v(�����3���e-���l�Y�-㥋G�`���܃�Ȅ]���8?�gh�����������m���rM`@~"�h��ţi������kk����̬�U3'��SE��Uj����!uRh)���>?b�t_P�A㢲o�T�Xc���}
}U.c�;1�
��;vSI��qB L�����;�1�_�e��2��TOl���y' 꾫%k�@5�C�L�K�y�,�S�<_.���&[E�U^�Y�(�w�c�p\�e��@�=��[Dep�Ԛ��|�K��(M�f+c�ש�x�����RCN����-m�9���Y�06τ��i��������Oh����>��Oe%7':��������OA�=�6�� ]:�P'�M�G��t�i0Ǧ�}$u�	�7�+zx�і�B�7ז���)��L)��N�0�"�dtLjص��"�A�"�[��w�'�N#�eO�������\-R٪��N?\���1Z�L��Ƥ���u�vCO��`v'�V�L��}��?�1���Hf����J���y<fh.��Ū��p	�U�݊<0��G��/����V�FI��h=�/�?Ȟ��f��,�Io"1ɰ�}Q�թ��$�`�t�
�'������E�>�nZ�5����ZB)��
�S%W=���5,�����8�K�"5�;�(a�_�g�;)x�}���xN���\M������X_��B�nX�BN�$l3.E[����y�L� �Q(�s�@ʁ1h����X���Jyo��ռ�Hr�z[���r`�M*�tx��c�Bj��޴c^:�wO�ËͲr�R
�7���nSk�a��J���6�E_fPE��T\�5����Ϳ%��| ���R*j�9Fg�$�n�Q����`��b)E	%	`�K�Ȍ�CQ��tO�ߙh�]!���$�uVǾ�P}����u�l7��d�2y�q��
N+���K��l�|LM�Ic�K!��!�����f�	b	���y��.@���o0q�8�m
eC�nN�b���,�T��8��xp�����6l�M>�4k�N�
�:V��vrU��G�ND�������D���-$dH�BDᮔ�w5����I��ڮe]WX�֎9�ej�tF�8��.Wk���l���7T��ə]�-�:�?��Ě��հ^���.-��@�)��/�&u��2��r�<����J�'���{�w4�pYz.J�c��Li"�b�8�|:�-2G�h�mi�7o5ϯb���r�_�k���+�`j̜��ït��Tio�U3���`���R�'���z^�Y/�9tLugz�؊��wF7�^��E���g���/(L�~�� ���I_���U[O�OӍ:�9���[�����+9��N���W��� �ȥ�tצ�u7���6g�������V;�^��V��C'����њ@M��:���lCHu#��>.%d'hf����C�%�5*[D&i��}[R��~��Xʹ���F��]��HE��Wl��J�Doh���O��)�O������ C'�o�I�Z%�ȡ_o�^N"9X�"�+���udHe3�ӱ��K �&>�wFZ��y��>4��m�#�Xo���P�����Ʊ������U#�s�Q_E&Mɦ���c���xW\�<���مG#R��E�QN<Q8���T=�AR�ck����)!«�������S�+}�-#:���3ƌh����ZL�<�_3D��/�̿*��7��:��dt.B~_Ԉ��YU����;Mm�v��<yw%i���<3k���o�g�ө��!_���[S�x���8S̍�1qn	`x/�Is9u)�����@�Kl��5_�P�`0��7j{�XXx�_���O�,e��4|
��+��g�Κ�����X�y!�4��,��UB�Q[�ј
�͂n���;��ɗk�h&1��\e�hӈ,s"����"��ҡ�Oҙ�;s
���c�������v��_à*��fS�εh�ۖ��ڑC���V���\CXf��VW5�B��V������_�T�:k!;�Q�}f��}��tN-l��g'��w�tt���4�$'TI��5βv��ajz<��9�4~��4]��N�	�mk�Ï�!�j��1	��,����a����]L���6�5�2݋��d��b��ch؃_�|�pE_0)rQ�Z�E`�pW�_��$�.@E�+��~=N���~���B�̩R'/Sf���*L�C|����J�=�'��z�K����4��ߪ���6J�zh�rxP�{nv&�p#�D�p�.�(�)�������Vd�����nҼ8x�ڄ�ˏ���P��,7�n�虤�q� ��]��5r.�����`�k�B�Ew =v[���;��]��i���u�>h�dn�J���J��Q��܍�C�x�mw`�?�Á��3x%̘��3:;pX���W�Pg����0�~�
�1֞BhS7*d?P� �h���af�h�j��_`������f�Igb|�!l"����p�K{��X#wK�	1��������-��Y�W��/��$		�r�7r��3D�E�!�\���Ȟ��0�Q��S3.a��1�_VZэ�v�"@��~�������0�+��p�8��2���H��P̝.���M��Vf/_�eO���嶀��ГH��)X�`Ŵ�av:eƤ?�O����<e�hΜ.�hҽ)�>SRȩ�c(»�x)��`��o����nݬ�D��(ʰW�3'�}O[K��+1�L��Г��禖[&Q��Z��=�A9�����k���Ө�Q0�Ll���(��36gJs���ּ�q�:V�'\�bJ^{�?��Ȏ�~֨Rc/R(#��_��4V��P!��v���V!���?� �8K�����w���;�AF����[�#��|�VLg��q�hC��!�g�m�?$;�Q�(a-W���Cc��>��Tե�_�aGIԳ��A������A�����-a�1Ј�5��$־�\A�e��'Bu��>7}�(����0m�d�*V����>�����z���p�a���� 䒆Җ��������I��;�e۝Cc�)����bF��#eaL_�iu�`�X��?��۫ʗf�;'�?���g`��NyoHn��A�S����.qC�&E���#���dX���(�AZ�f��p$�ab͝�	6�2������'`nL���C�Y��L��:=�q����֗�v�׳ {O�Ap��Tn����0T�l�%)�� ^�
@a�7���]�A4���c�q$&�܇I5���c�Bʻr_aw?پ�����f��\�;�iYc���C��-�6���w�D�ȱ�!,Kc���'cI_��)�4����a����՜,
������~�T�[5�C�qy��r�WF4-h<�F;�]�e=0���^)�����K6���f#l�>7�.�f�����8$o��K�n8s�[N+填��q�{o�6�~O!cF��|��bP/M-��t1땊
�,���N�?����.���ˌ�;��jN8�{a1�
��Ƽ�7,�Ih>g�$����`�3sY��5f��y���z��D���Pi:��^�Z��#Mc�(�D�[�"Ui�k�P÷��U?t���w��$4�~hF4 .mﰜš�e����5oŮ��{m�Ё)28�HnL�a;�>L�ؒ0SO������T�Q�xsk�0G�`_�A�����X%�l��dD! ��?��I��
eP����5����9�����	�3�q䟥L��쁥P3��|��a��;��}AJA����Q�ٴ����I��?�y�����NQ�o�7�I�h�õ���Ŧ���ﱟN��*ՠ�c{���N�Ss�>�Ŗ�! ���M��Ո�i��,2�.X���e���_��' �_��2lT�ۥ�3+b�r�� ��Nd�F����7
y�F����6�5���9O�-Z�#��OJ�EMz�Cc�?"	�,;�h̎�Ѫ4�)�k��A���� G�O����I������ld��	/��0S�c���G]L�� �B�o�l}'0Z�w�a��=�N��c찡�c1ZS˙�@�	�`�ނe�y��BC��<����f��QFj�1�\��N�j�jyZ�A ��q�p8��-��$̺��c"Y1 �J�vtsc����%�'�+�e�Ӻ�k���v<H�[��[W��aܥH�拃v;f^��`�A//S���L�=c�Eq�J����M���� �!��.��b�h߯�_ZH���AA�7ڿC�Z����֪��KK�˯���(�b�o f�r1 ��)S����
p�1j��!Z�v����8���J�B�j JTUH�7��A-�.�W�E���楝µޛ���&�k\J�|����<j(�KV�Mz�N��"�Tf�l��YTv9ɾؾcH�	���/#[KY�Q�n:���n�	~��M��V�ٕ]ք�j|ɵ���b#��ѵ��/��Q�jOQ���)]�g/cW�������6�.(�v]h�g����^����������LV���z ��|����Qn�f���Sţ�n����{ƢC�f`�����H<�]O��!�b��!��}��|ī[*�O�)u7q��B�|�[[� F�
��6�	�p�&�j�y�-�\�/��$nW">z��g�5P�)�.�s�L��[עZ/�A�RZl{�܋�Š�f��g��9Yb�lk�F��9��D4F>�Cן��.n��i�dNF�i%�c��0C(¥�Iwp�Y�0����ą�\��E����n����`��&9�\sx��;`v�OT%���B����Ϛ�jy������c���"���1�~�cT��4�f�xNKx1Qǅ8<b���X+�Z]�-��|�,����d����o�hu��)��8�pP�5k��#��k%�����jH9.��vr"��3�F�Ļ�hU?A��]B{�4DPSJS��GV�-�Y���cx�L5^�'�+�l2G4��&U�Ą��g��A��mu��4?It��&�q����|�ɴ�I��&����M&���hyh���B��.�*��B4��ʶ�Q�|ϰD��澗g �Wߧ����י8�p3(i	�&_r��"n�����^�6�	� b̐9�nϏ��\\$�Ч����~��y�8¬TJ��EN�ATr?+@Dy����u;$5�q����53y��I�Z��l��lZ�(�1j�u%�$T?�ܙ9���L�d����>kPau�K�ᙷ�$a3�OV�;ú��C����C��ʾ���EN4)#?㿧���)*:r�����ǂ����O���Pt��y	G��x.F��Ijŀ*S�&~I�u���lKpc�v�����U��[,ý�?��j��ߥ�/��L���� \��Ң���d�W����b	���O��O� ��޼�L�͝��I�,�b�!��"�2{u�'��	G7��S��h���߽�Z#��{FĊuf�W'�$��e���Y������e��X�	VY��vH�cݏ�-CB!�W��Bϴ;�\~��8ҮG�U�����֨��_�{��nu�[]��61()/���H����O�0j���B�^`.JO�Y]B$Ђ���9�_ރ��i��`ƕƌ�'���.�!�lAaiz</+����-y���,�_����rZ+�H2�����}L�ʄ��v��
��M�0Ҏ�\�:l\�	�;��j�FT�`�/�ϩ���-	ib��ɮ��b�=h���B��4�(����E���*�{h.=k�V�m��8�9:�/&���R��.=�5�d5�����쒱���&��*x�PjЦ�`�v[߇�>�`��BVJ�e¨�z�6יb�=���1�s~�]0����Y���8��2���I��,a�)d�X��6M�u��u,]x9ؑ�����Q���D@�� �`ϊD���C�;i�L�m��?���������a�/����@�A�Ƞn޵D5�:k���xhXw�@�2�#�fBL�=D�����<���8���6�i����o���ǧOݺc��sQ�����]2]�i�qK�b�-٠��@���G��^K��zM��y���C��[J��K5Mu�a��Vq��l�)�X�`�����-�}'�H�a\������X>O9�>yW�tT��XS����ă��UƗKܘy[�%0����y��	C��7�@J>^E�o�ݷX<��w��,�`ܧ��y�5V�HZ�  w�Z��fT"���&|�y�;�/h<덁|0Y�4b������B���h�ײ։ew���mQ{��a`j���]/r]��v]^!�O4����TpP�H8����K�TpDq|C����A+�#e��}1�����/�>_����~�3��Fz���[O��O�֔��^�h�sƯ�	FX}3�_p�U���%�2��"/���e��;ot�$��u�|]8�91ZQo]O��45\(�5T�yP I���㢽�!���E�Э0Q�O;,����P0�@!PU�).���=`����@�.y�S�
3�K�?�5uJ4Bð�L5	�z���VOb-NqK��B�!���RZ�kp��Ӧ���+)�%0��x�~ο�خ�����Z-�ʅ�w�1�?�u�������\��
����9�@�O������a��v��D�`�C�o<�.r9�ю:v�Zy��y>��)��#k`�
D	��kY��&�D����ի�?�,P>�t�=*Z�_�	��/2-BC=�X��<QgQ`�o���1M���Fi��eX��7o�%$�ғ�jYU[S���1&�B"R��4B�A\������-�:��t�6TE�P���w�
�D�ؚD𾚚���`�/����q>;�+Lw��-OW2��I'D����^m�Ȯ�Z���Po�dKZX�>��Wpr�3.ۿZ�)�`L2�ad�1L�oC��k����@�%���6��S�z~p�Ð�0�vJ��wk�4(t+;"�9/�^%h��ϲ���:	��*�g`)A����[�1�F��j�O�ǘ�_��P�YX��P];�S^�
a�6�2����d�������;N߮X��XMq[�ģY�����B�m4��SԐq� ]7}�q'�N�f�J����E����b����R-8y���6]#�l�s{T�EN�0����)�(R5�㍖O���uZ�d_�t&�N�*3vE	q�ҩ���f����v�������z�&ɔx<�?��,H��w=�J3}���ɠ1D�(]"(V�����r�}-i Ï7E+a�
dF��-:����DI)��0�\��+�q%�DH��(ٱt|��f����{VDK�h/
��~q?7�b��	��ߟ�K67-S�Z�,�O�K��+�v�����3�Gkу��(��h*��"����YY�q����<��|?�yZ�&@G��Hh�����0��<��;[	�Ѵ}u�y�WqTpk�:�g����*�k_���Z<1K.��/�;�JenبnT�������Xt(XW�ȥ���VN�l�G�5���{�n,,@�KݨCuuI����[{�g�64�g~�E���F�%����Y�hr�ǘ6��j_�#J�]��z,�'%���~�R���RaK��&�c����C:#�>+rIO�SfuV��-�ΠMEu/s<�>�k�遰f�-����L��R4����K��'B�p=ExZ6E�����(���F
{��4�hT�Qf23{���}9S~�ѵ$]x�#��)g	e��+��n���s��N�?�����w��a =������GL�}�b�/Nr���1�a�oy�J�*3�<r�G�զE�K�Xy(S��ʱ�4�O�iB/�Ɛ�r�Ј�d�s�0���f�Fߤ��)+w�ȿS�LYk�o[<����C<��4ayw��M����Z�<u;��e���8�@*�}]��}�Ay��d|�r�h�B v�ѯˬC1%<~E8�%����z8α����d\����ZK�ZQ��
c\��.��5�|�k������?����A��4�bR�8�[h�^�:�����: ������х��zW��.��$�~��`�ET��I����v���F!�$@A`h G���S�J3�'�-���62�2�E�R��m�v��߮���9�s&E]-ת����t�?55}�p6Q&���O_�ꕩSo�n��%䘒���^�;����:]��7*EE��u�X����3Tu���?��n���:��Θ���΄��ա����n��""��'���9X����� b� ZX��e�tlɊ�V	��ݚ��p�h�~�9j��$��C��<����&�0�N'd��M��QE�g���!��nr�b��5���K�,~��9�Jxt�zcď�Si�O���_lL��7P��KXK#	��iE �>�E�΅�:���c��xVY��_>��s.�VS���=�od���,�'�,��5���6@�o-ъ�3�9���O�}���̳���I�Q��h��jvs�Z��p[�D���F��;� q����	Z��X�T��c����wSj.�K�����<��5J�M]��� |������.�]4S�&Y#�?˼�5�AL4�.�T\{w����XFH����>J�j�� ���8�#4�=է�����e���I	h(�Zeu���G�L��`9�&��������5����`����t
��	n 43N���㜨�G���0$��xW��yl�*�#�C�1�}��)������|\=0�f�6�L��#D+��-�!0�����Y�I�"�aN��,�_���ܖ$8!F����g�Z(sT�-�|���;�)��.�Q�<�p�&'�X|ݩ�'�N�B�}��vI#����ŀ�3A�0V7��t�)�@�P�ӧJ�=H��`ӣ��큃��d[�}5x��#_(���x5�_b��`K��'&L�Q#l!U�L��m�ǯ��A�U\�v+��+�u6�F���7���
]��Tu�@d��#��
<���}z����[U0@��ߥ��_���+*��\�Zr+J��5�C�ԀP��^��(ǔp�\Q��A�
`���/�V��)���`���Ը��)��DO|������_����yR&Y?��T�a'>8̮�롯�g�X���sJ6�ˑř�.;�^��E�쫵�3P+1�ArY�O�yO+i2�����2�g���'�{ZS�䄓c��|e��}H�=M�W��Y����A��um��z5&"�D_ͣ����'��OЫ�Y���<`W�Vf�0��A���W�ܾqj������񣱺#�ٔnW8���lCD��4��EK��λZ�|_Z�"�%�vc7�1����S{%K'*
�W?l���Ls ʳ&�v�{��;��Kdɧ�����LS���5�k���9j�������|��usz%[#�����_���D�6n-��{"w<����O�Js�
P�9�=n�~8�����
+)�Ճ�cB���q�9urf�5ah04P��FfA�O�O5�-=uE������au�4L9�����Q�tυڴ�#Db��ױΓS��〱��z���n�@Y��@��+���J-vg��+-����������~8&gA�f�=#@tm�%�	��U��}a�̍)�lKKH����A���2���m����ֻ��b�G�]�Д�6��A=k��yf��|������3�n�x����'
˱
��0{�*\�u��U�K= ���ؾ<���RS�N����F�垳rB�3�ፇ������-x� ����nx�~>�� tǩ6f��g��/�97"�d�pj:+N���]UP�S�p���P2�l����A�uHvHfXq��މ����<�l�"*?��A�A���ގ�9>L~E�8������Z~���%�������۞�Cro��x��;�~aw�k���x���������Kk���kJz9U?|��	uOh%Xc�0�λ��#�|#  (~��/�Gg�|-bɨj�X��Ao��! �mρٙ����@�|�*��IYJj��2���l����J�%k��Y���]��\6>��[��U�-*�t�kw�ܩ�5��/�#d�D<��*S�1�ꮘ���R�ǴtV3�xm՝���) ��yÀ���V���5#�'����i����s� ��g���c� �Fne<��R��)D5��W��u4�]�����<f�Io��{�l4Вsq,k>��m��Ϯ�a��}.��w`������G0kH�)��k+�_v��J�:n��{q��>?��)1�W��ւ0��`]>3��P$�?֪:�Ĺ{4$������<f��0|%��-�Q�J�M�~�F�D�/�7�[��Gбi�u$E�/���Tz�f9��vM� _y�{���#�mx!�{�Fo��J��e4�-���ϒ�m?�e� [���W�9f�+K��ТZB���Ӽ�_ͿC�r�m��xȯ~ԁ}_�E��Wb���R]�8!lN�3hg;���Ƞ��L��v�5>wڄ!i�E�a.q��Ez�������@�f����W���ɋ8�
r^����I&H�~a��	����}���lcϞݟ>��_��}ߔ��C{�Be�6�S�,��Ș�t#�˔�&�i��b��z,��Tې3%f~*(2�Qh<5�ŲKݘ�+s�J!��Fլ�� O]slOX[�nm�s��=R2���An�8��t�
tBGM6�u��F 
q`[��eR~M��A��wĒ%�����n�?;g�B��b�EP��}HF�U�b�D��O�I�d��a�>N�o�i�˪3���j�«�Pzw�^ I���r�����'-�"�˛��d�}�I	�t�ZL]�h�m$��<O�d�i�|�ƯAa�*������;��ڬI ��+RZ���N��pP����H��R��*��NLV-ZUF��I�>ȑ"��zQ��r	5�+��0�ɿ��j#.𸟻oA.>4pa1��C��l!y���ʻ�;�.��A��d��w������k�!�%r��w6Ꝫ�d\Z�x��s}�
[�S�ٺp��:�Gb[�̢k���ke~��N�|����wZB@q�'��Y��\�tDj`�~f���hy��>����yk��4.�^�QͶ��4s�g� �ZU��A�1N��|��0�!�P�K��f��2�^�������1�����6�"c�N��@�z6���ލ��1�F�I�#�q����{ӕ)�.�.+9��OAl�|�?)��<9u�JN����GPm�i�������X�H��e�qU�R��ѕߗ��;��S���a�I��_���gkM�������$~I��}e�cX�؊0�����"aQ�&������y�� _}��Ek��*��`���'J�
RXdd�#��Mo�`�L���`�m<����9p�'�)�fMM;��Qω�>~N�CF9h��� �K�>�N�a���s<��hhq��%s�DlD��o���)�==��6�QX��ö��o�B���|�s\7���e6��V;��9�S��B́e��`nM�Sv3^Ef9�Y�>{w�,�* 1�Ɍ��+Γ�v���NZ�0FmT��񑾔�T�X��=m�����#yD���ޝ;QNp�0b]�F>h�r����g�-/P����c��3��=֖�
Vrl�hӖI3Yk�i�|�Zx|8���[9�&�\����Lg]u�cΊ���O��5Q;�>�����µ��@��Wo��@�F�d�ۡnB��?4�/{��<Z����S�2�q�뙾h9n�aDl]���ޭ��n-�,#	4����a�$��f�ᣲ��aײ�aڒ8��4��ȴ���4����SyA1Z���1�d�O6��ǖ轕 �z/K ����[�C�?�X�B���4� y+�'��X��6���l�����5\_LDj(�Pp=���[�]�&%W	��\�Nʄ��TS5$���Kzp�[+���9�}�[,�F�K���y��5���v��� 6�e�	J��Z�a�N�@�h,?�@&z��@8�w� |��]�*�[��x0_91���bz��o�Sa1���y���W֠� ���S��8��=\��pZv�S��[T�^x�ME'�Ւ?��8nJe����TD�����(�jVj4�j���h���U��=�/��$���^����-@�E� ~+�r3�Q$ �&D�C�ZS��1���	4=��4b��	�CRΘ{��+5穰\�R�%��O�s+�.�0}K�3��%��~!���WGE��e�+=;	3��Y���S6*��6�?�^<]U�?	�&��a�J�"~�Az&`�����|��w����D
��'�������/��s�u��>�䭱6�"x|~�H���a��G�섿��<;�:�s��r��b�-q�v��6�F4�t�n�5��S� [�M��c�sy�0�1�Chy(9�6�hX�s�)��H��cڳ}Hu;_���#��[F�ʝ�n\oiӓF�|��&iH �R��K<��#�
�}���K����h�%@���kY�v���Z���H�ӵ��B$�q$fr>GѨ%�=�Ĳ��i2_YqE�AXRjU�2ǁ�5@��P+qd����
�A�޻����(�tm�'(�S��V�
��&� |�-����`4�v�����f	4�XIL%}/���KF�;Y��i�E]ԫe�ۄr�O�O�4���vk��d /�f�8�����i��4���Ǚ�4�T��\��>x|&-����8�ϟL)�9�q�n�y`�,V.�0V5^� bu����7�I��->S��y?��l���
��1~M��'S�3�N��43�\��S84�$ۻM7hiW�֌*#I����u�Y�r���tM����ţ?���J�w���x��Z����t�,�W��Yj X=��Kd��ȯ]�>Єg�N'�$��J��0-Qʕ���Q���ޕ"E���c,*҄�56��iuN���q��ή�[q��b��}�	yu�@���S��<��|�vrŨ��q1o_�w�s�+��������{e� Ҳ��$�ԝ�n���	;":�(2Z�\��kO����}�!�!D�C��S·EKm�P�d��#��O�X�@eZy� ���#O��_L7dK�g�֟���wD��<a�{���:�_�NA�[��7V\pY
�� qi�,ٷ73:�]��������e�8z���������T5�����p{5y��'��l4��k��WK�l�nWmY4{-����B���=.8I�h�����Bڻx?�96�C�Z�.��T�}�7��� E����rpIxՉ��v������j���vz�(y*��G��yܲ�R/��%�}�>������oʚ|�w��J�5�T_x��nY�(1�c2�b��M4/�+��i�^Ɗ8���%u	�3��ͼ&�%)�@A ��b̬��P�����MjI�����k�)9Qf������OdK�0�~���r�݇lU���uP��K��u׏���F�udS�.&���(E��+e�:P�#*�՟����&!9��i	�����H	�p�ӷ���݄��b�rT�;��sBӦ΅G�m2T�Kq&�ܙ�p�1umв�����Y��A*�7Х�X��l���ت|hC	�y�Y�-�\��N�yr��5��ǻ�yP�d�S����*�;gl����I��'���9l�0\��k��=5ʂ����3U�$�sba�W!��j��7��N��u���g��i�t�
x"ɞ/�UGˁi�9�ON���$
�Bl��R1];�4�^��Rx��m=ƻz���ӷ8�챷n���qo���V1�N�A�gK�(8��f-XS�â�G��Û�jk��Sk�>1� u�֋�3�L2�jæ�N���������M�
�CA�.�5 R7И ��O����K���tF�ޅ��X�,,/?� h.�E)�:fOu�^!�R*Ұ���WƏW��%ee�'������h�:�1{Qh�?��P
S$�,��$P`����N��޹I�*�~�s%m{����+Rp^M�Y�&Y�����0ñ�K9����]�b��xF3X��R�/�|�J����� �!��[��&>l��)�.��5kTJ���tE�����sQ�y�(�J�Vxk�A<ʺnQ[f�~0���t�C��u,ؘ�J�9ȧ��V�N�����̜n������]Mj�/��h�&��$R�~Q�$�1}LEVF�*�))u
���|�U��!�OQ�WC�p��;���H'y���/����$��j������y���>��f�C�H`8�d6eHq�|�����r"��lEʈM</7^[����	��G��3wy�p��͞�Y#%9lQv�vĩ�e=������ LW�D���Y�����έ�	!τ�'�^ ��AA����k^>��kɢ�m��3���ɳl�m�%&�Q���(��� /N�uw�m�̳��O��*�����Y\]Zk+�:Z��2���<���R�E���kqt�7�7M���Q�G׮�.�]��6b�֢g�ۏ�W�)�Kq8�Ki��`��x��I�X�L�f��%�v&w�췪�c=�R �"��;0�x��O�,�ͪ�� �O� r��u5�n����3�Z�&�*j��g��2�/�Wh.Z����,��X�S� �P�0_����h��?CfJ��N���{9�����C���'���fg�m�_�������R��
xH�����.# �0�R��i	�V�1b��=,���ɱ�����wb��.���3�'T9�"o��¡���`Ԃ���iI�Ҷ�ǅH�3HQʨ�}�&6�I��O���Z�qL�Qv�W�g.��A��n���4v�-�v��?�ъ�p�U~w<x�m��&��gZ��绲z"��~�grl���7G�I2S�!Ғ�3*qp�F`2=gɦk]22=��j�b�]��؟C��3��~��W�:�Q2|��OoC2=$8`� ��1��j�n���W0��̈ҹ��G�:0h����}��A�γ�bƂ3�0��0יX�Ez��x�6_.8?Re�f*�M�c�Gh2D��7 �`��m�+�/�܆X:��QɅߦ��<щ��K���<d�(GHb*�ƚ���|�<T��h'H������4�G�!�|�@f�ƖCh2���a�->#�M�RI�Ҕ�g7n�q��eû������$]$\�H�7k��M�t�$�.Dن��v�V�7���h9p�>"A9�5s����Z7�b��}��Z>�&�g!j�얊𻔿��G��r���*��g)��p�
������0���}2Bx~��t%^�Z��m&�{Ɨ�ካd~L����Sx�����sg�6iVThEG���}�M�1~�G*�	R������5w
�ƪ�&��g^���Ww�*k��UOT���B���4��',
��Z$�km(s��WW��ȿA����"���e���#�����N,E/��9wȳ���c�W�7*"[|ȹ�$���}=!)ʔ���[�X��$	�)-�暸�uA$�l�Q�lʹt�%�h��j� �F��R��R��ƥwv����_�lu'N+@p�{p_N���F�3V���xp5�&���ǌ�e�X��)�0T�ď4��{ ����S��>q���+7��+KfQ��bv���9�;.�?����V\G�[/��#(^�D�J�"%�(O�!��zd��_f� � �oWx"�o��L���eEj����mG=�Knu�R(Ms?0ؾ�I���! �h/_5��p�ͻ|��,j�v�Y��?*"~cq�?fzR���(	��M#�1�0��H�jU����i�'���5U7�\�{sO�j1[[Ho�)�9s�/�V�I1�r�ߥ��E:�;�_���������%�DO44�ܓ��hi�Ky� i���6�]a%�Ҟ���=���ڄ���:�iF�iE�)?H?N�s�3���5�ѵ����Y����q���V7���D	�:���Ź��9T��m�]�W�R�d��6BK���B>D�b�+�<���=����`c1�3o���m��V[�b��d�)�\5��l�B�~Vє��К� �ȑvk�3��vk-W�2��y>��*�����L���Ǧ%�y����b�FI)l�Y�!i�_����9�i2fa���7��xEuD��u4��<�����u���Z��G ��4����2u��M,�{�T�D
�u�g�	Tz�덕�Ѓ�~���R�_VX6#���f��3B�T��E��el�wL�:��������.1�ͱ��S��
�f�XF0��	��Q�,�|ٺi�uOT��ڮP:'�v�������A�����;�P��$��~������X�<&��?5��j�������w%�a��zF��9��{�[4� �7�NO�7a��#�։KBY����h��x_��sF(�?�4��+	�;*�T1
����<�6%�ɿ�e�'�t;cǠn]�S�NK��?�Z��j~.,g�����8��d�. �H��%K�zM����{R:�tCZx=��F�-^� �{�k�wK��
=do\y�J��j`I�J�1#��t�@�6���H	z@=��O�W��/[M�v��0���z�q��5혖(<��^�]w#:�NgZ�a���J(�帐����G�AZiR����8�*�@ AЭ�CP�3B�sc#w�S�L�kvKC�TQ�{%��b�~+��d=����8�v&���A��'��xh���,;���-��?���@!Nk5_r#���U����{�,��he���S|=<��@��A�b��};.-d�3f��}e���Q8?�����<��G㊴@��UaB�Ii�5)쭖�HU���$��G�G-���3Y���\�t���B�" �Bp�g�1�j5s�?�(� ��pt��	�"�W�A�����x̆�^s9�Ъܭ�P�v:ޜ��|So��T�l�����Ej<t��ܒ��g�TV?�0z����?�d'�1�f�44���Xנ,t��x�0���k���� ��V掞��o�Ná?l�D�J���$��D�;F��{�6���Gv���O���ʱ���!t֧�8$b�(P�nNs6��P��}��Q$���K���V� )E����M�f��f�*�\�-�pAⓔ9�	J��y���, 2}oz}q?2a�9{i���/f�Fb���W���j�>�1�.!��r��lW��ٲ_X4�����Ž\���=\\Hq��
��'3u��ه��OV�~�Gßg�-�ֹ�S�dF��$M6"'��G� �dw�i��[�ϳ���>���D����>,���s�[��3���s� ��W}:���'���]��K�yJz։tG	����8���	��2$�����0?�4�4���P/�R��dY5ݽEC�X��i;k���y`�W�A�P��bHf�[����,��t<Oͳ��}׀��h��^n�߆�z$ck��E!S��Mn���!��?���p����������ţm=�'05F��j�$Ⱥ�(I�6ʳ�糠s�j�`�Q<3�
H��-�4ry9�m����X*��P���c^����ڡ�*�������0�$g����qퟷ0����e׊2Rd. ,&݋_u���6�~&�#�ڳp�P=|������`.G��Ц�|��f5���s��?�$�K����MH2��!x��^c ��j�����Uy�G����f����L��9�;�S��I��JO�Q)�J�o ^ڴ
���j-^Gkڶ1Ect)]�W�~y��???m�uM|g2'`��	]�M�(��X炕>� Hm��!lI��g���h|�nÿ�k���	����>��f�>����w��fX���4��4�|+���ș�麒˕��"����z���t�?����6�u����CV}(�րg=ί�q�B�C�ߺSe�i���CcF��j}N�����ܾw����]�  v�M��A��A(��5OЀ��L)R�
z�n5ڰ���ԇ��:�
%��^X��C[��X0G�r�P%���V��oS��呰 7#�#V��Τ�Nj@���-[PvH�@X-�i�L	�3^}�0�Y�2p"mC�B�4�Z�x!$����$F!�'��&�v]f�_��^���N4��S��7F)�$K�0��A<g���sDύf�aß��U:P��|���Y6�h|��J���&8e5�Foҿ]�u���+l1{p����-�c�&�p�e��e�v���{�:_<��d�}W�6}��L��Z�I�F�Z�F0�s�L��{�i�_��m��~'�Ow�vf���9D4��w�w�*v��<A�-��c��
��"���>�7��>��-I��ϴ�Q�+�Ԡ@�6��_�8��s*qh�[rB�RJ`x���� �(0�y.ë���yb����\r=�V�+K�L� �y���K���px��?*�U�ͩ
�+2-��b�k�� jPxH Ѫ$ϳv��֘�	e�Y�<���E@g��b,
r����p!FQ��{��������D�`]��:�=vK�����4��]_��	�f*]�&;{{��9�;h�K�Mm7)�k�1�o��T���w�WV��nǳ���O���b��,� v�(��%��t�;9�ї�6{�l1�CI���6 �W�<\�e����ҳ!���?.��A�,�DX����pQS:��րg�:h�#�e�K����N��?�,���nS�9/aի� �D��@yxBJ��G����+���BS�0����Ĭ����ۙ�㜰̪��$����=9�%?:��y��.Ds#� da|�I���0Fz
��]�J���R��J3u�&ϱߗ)o�	S�T��\�F�c���te�����M�C�ځ�4���v��Ұ�ג
�?����N�P\[U�|@�@=���we �Zn�v�ZZ�ct�<=��>��+8�rX<�؉���j~�e�	��L��������a*�)wQCt-�X-�/2��w`)e����� q�Ɖէ���ԣ�����wZd3��~@I�a�f�R���Q1غ�$��tT��yқ(����>���E7�}�wbf;�6\��6��
�'�i.�����#�	;��k�tK/���������b]���4��Q+4
!д����0���	:���q�|8un�{O��V~z�����1�AEp�f�%Q_ծ�q�ܖf�x�련�U���W���ې��),ɔ�H1aKW(���	���r��Z0����+I�%g��a9e�����x�X2n�m�4��1t5	��]a�C�د����:��:�"��Iel����h?�R�V�͞���e]�7Q��������t�Lꗧ���PJ:����Në��Et�H����Gz,wO@�`I0�y�)��Q��Zo �)���h�$�ݯ���I�О�sĝUȋ�,�X�{��|������zN�@�y��5TE�}�����u�� ��!ϼ����_���*�X#9��Y�
�w���t������M������8����iK�D� �:�1,Ϩ�����v��2�B��~`���� �Up�w��Q���y�Q��[���Ϯ�E+���d2�J����A�bePi���_��s�r�i�.c��'7K	�w��$j;��ew�%
��8`W�g:/��;�g+\�G#	*J�[W@�$"�ϳ��1��f�t�)�M��l:��N��0ß2��I-U�7���Q��D>2��!�, ���\�hW�쑾��U�7� {��uY/"��%��Gг���_Zr�ұ�EM7����T��B[~`����1j�_�n3��1�������yb!�o��qV�rNr0���O�}����M�<o�|�)��Z��pKiP鯺j�a^�f����~��
�7R�

�4TP2qN�aԢ����c0T�eK�A�)C�G�J)���7%�����  A����=}�x�\̡����Ф�P�E�_���z��~_��`��1����g�
�s6z��F����|�'�rp��-y
������kRY��m�'U�j��	��+������f>��x���C��g�:)�������މpʲ�����녹c��r8������@�.ePx]B��ei���\�a�EN�%�E竜W��?Z�a_�6hb�X��-��%C{V>����Q�$$V���z0��`��y3`J/E�	x�K���-�9�+�H��D��*5����<!i#�o3��f k�ͪ�K����]����,����	�q�jnz��[���<�Nύ�0�5L�e2������Of/ ���h�_'x�Q�ƀ��W̈́�W|t�'�
��y�Y�*���A;��d�C�r�Jտ*�����-�A^��{��
�kh�C�iEY�V�]����1�"�E�D�;8�p!�.aU�y��C#UE8x�L�0�H�}�ɶ	ٓk��5�����SA����a	x��	p�L	)G��*Q�B���;q�m#͝�y�!�:m# enل�jH�h��w'8�.�aM1��g�q��F���,P6fS!�$�O�G/P�y�_����nIx�S�昘gh_����Ʃ�0��[Q�cv�S�;�F���s�}xf�F�رͨ^8�[��}gd�#�W푧It��S\��U���o�:!d,�i|Ms��|I�Ꙑej���D-�{NOS���W��:F �Z`����l�vF_%��27��ʁ���U�h2ф���󑋔��Ɍ1*�!M"�����+���H�������D�/�*,B�__����2��ٲЭrɋ�G���yk���<����2�3b�4ED-Gड] ��e*Ze+E������xvڟ6,V�]b���m��0�"l��P	V��x}G�"Em�"ₛ�厹�� U$& T�g���V���W��V�>��0���R�1���f�߬ǒ1��wl@V����3�m0�n��g����&@LUNC�X���0�y�-K����r���Ѷ(����*���ּ�6Y�V�#z�D`����S�;M��8����\D���m%3d��*M�p��w֓�gVgSH�Lyh]*���U��R9�:���_&�
�tH�B�$�/�R�@��D��Cbb��f�>�Vf�!Y*t��Y�a�Ϩ��tEC�=��Ų9�!�T�!�b���uO�eF��:��u�+<"��c/DjC�=�U,��Fn{E஽�[vwex��p���Y�!��N�n�t�0�.v	Oӌ��膛�NGm�m�A�_��� I��Ԋ��0Yi0B7z�*���o�
Y;�݉���4=j������!ts�(�rW�?p(vñn�1�I��xAq���(�^&��ݼ���̀�^���~=�n�R�.�a��If�r��=0 ;���!nB�śt=}᎓g�ߐ�eQ-�]��J�5ЍlҨ�2i8����5L�!��MSYF��rB3lB'�;"���x�أ�8ֵ�kMr�Sy������y|.Z_�G@��o+�2�ǅ�񜴃@o�)�p�=���ԣ��#����U�(���;�z�;��
/^Lg3�Fg3�6��LO�9�V!QL�Eet(���]��;�Ն�4���7ПDQ�;h�lT|���t���kmY�<QõQ� �(�e]�Edq��39TM�W3ҫ�>O����,�<s��8�[J("��g+I�]� ����N��Q���.���&�+��2
�qu:�np�Q��ʡ�g��9R�Ug7��������c��p��
,�5��g�ԛ"�<�O׺� ��j/
�lQ�?%5za�w���G�d>0㛺��N��<�R��&��K�u�,��%�8�B˾�v.N�5j�]33��?b�$1�_����LJ��5j9�S5Ц�r}���	=��wO�H)Ď=�ħb�2mmt̼\�:vt����n6+���b�A�9�EL�l���޷=څ���A�`z�X8�!.�������n�nRxy�/Q�n���2���3?�4�T<,�>��L&Z�/.�*ްB̅�)
,�7"2nHW'���;�&߰��L�ߖB��ʦ�>BN�B�b���*c����cDߺ�#�>�.1�@U=�L$�1�h��� s�A�Zђ�a< 횄���O:+�T�B`g�z�K�sp�,)]���/��G��� �9�!q���Z��@� n���$���4�hE��������r�{���&�c��`/:Λ�D�b ����[��8��p^�SoG<��A���e& W��PT爓Z�)m�n>�+���h�d:�Oc9^�p�;)�N�&Qg?��d��Q�gХґ���k�\�C�俻n0?ҹ���ATbO����D!E�� Υ��3��R{��߁��0t
؎��K�A�QG�&=H�5*;��2(?�H˝��ײh=
hs>Wk����|x-D�����R$;S��2>B��i�����ӌ,��A*�CKv��A�Z��q������@�:x4��X���Ҳ�4�/�Tu���ƚ{}�-~�!7���ɼ��L�Hb��!ͣV[��ثGş.82މϠn�q]� �K���[�d���0�ģ����Wh���2��q�_��q�N�v��Ppn㉵Š.2��_(K�.�jM�G�/�߳�`|��03ǿ��M��(�UTrz���։M�]�K�SS]��Vl��R��,�o*`�=E �x��a�A/�����D���bۖYS��t�w��	�{��!{�T/�OWӭ�� ��
����\>��n�L�f�R�d���t��QI���"}T����{�ڧ�0�-]�?�@	��S_����P� S��u��ϓ��w}S�1��{AWB��0b���/F��p(��P�r���pN�A�P
��4��[�{����q���Hf�Pb2�J�e:����\,���M^�:�î�<�xj��O��N�op 8�q#������\����P�tQw����^��J|��\�
���]a���
s/�ۻ�2��]Tgq+v 淫_��ZDdk-DSz�r�kV�b�S0���uheC	��=d@d=v����QؿR�F��b�DN#����eQ�fN�g�������w���[���������؊��� �5`�_41nH�˿�&�-*�����	�da��mT �-����m[0;�[_B�h����J�L��Ra &��k:r:$/\[�'��P�wy�Ý���� ���5h x���҉"�,����zix�!�D/�F�4o�c%c�͟�_:�a���~�%-ƄǊ]�3zM�5���:*`��0z��FQ;��׊������x��0���#b���\���$߻����b'�z������:N�|�����e��u��n$�N��\*�2T��p�X�rM���7��A`��w������@8�\0�=�Ʒ�5J�0���:v0���s0c
������d;�flYx�CRR3��_�Z�A����0\7��ћ�M>]L17��ߝ,�3L4	��[�D� ��z׈5�nϿ_�D��U@�:��mb�@��1�N�[`� �u����;>�(0����Y�|�BJ9��}0��d$���-4��Y^�`�z������ggb#/r�߻�h�fzK>C�`��D��Ae\P�\����I��U��d= sr�����+��װ6?����%BC2HB�)�ԺB���=^�κ�����7���h����)�(�z�>��.��X����B`���[*��$1A���)�|4�/������RY�X�W9��I5S.��<�0�I�i���0`�)�w#���X�LK<f_�a�9�^3mm�^������L�LؼuN�xπP���6��x�g�j{��՚��tѬ'R�;��څ��D�{K�=���>�����w�[�]�g����_�X��U��Qʫ�?�v�`n��К�'+�G�X�Y^�����0>t]A��42����R71�傗���3�aP��`ay1��.b\�Ty���!���oo1�\r�/T�DIs6d���l!���6�@�D��� 7au2"m�2�J��
������.�?���z�����Z|m�ʱ�!}�{���:\�����"���*�[�ͪm"ό[��d���-Ц��]Ŷ���yf4*g]<��HU�,5_�>7m�G!��+p��PA����2V��r�W���W.��A� 8@;JEUiZ1R�R�f���� �_�9���g�a�:���1��r8 ��:�~�[N�P� b�� �����[�έæ���F��I�lyg������/��v��'�?_X!�&[����@�À����#��;�B��"a����Gx �n��62E��12��g���;�vJ�MC���)��{�{��e�oo �Ls���{�$�˃�Kgb��4�vRf;���j:�#ʍ�F�:�	�e���s�����R�9%�.�mYD���@�%�Ǿ�������O�eC&قs�WN�s�!�_�w}S"�A�&��B% *ܗA�(��8�8l}����{�q�cC>x)��Eɹ�I�� _N������s�҅^í,����O�'u?w{��/��*Bz�r�}���&��d��u˥s�������]��O��+v�b���W/@TB��А��3Pe��G>,�r9�@z�휐o��s,A¨�s�(@FX�g����X����b����E/������+u8����CK&�T$ើM�(>�9%�kh���������D]��q@N6#7s��I���x�W������)A���m�J$��/q�{�S��4��Ҭ".@ l��2oPe�E-~p�8d�IJ���FZ� ��crD�5��Qd!Z���l6w\��2�BX�z��T:����4��,`�s�FGFj��q�q�Y/�q�<؇7K|Y������_΂�`�W��x�}��۲S��h��;Ɯ�O*uj��]meR�cZM	�S�����
"Vܧ�@��z�R�~�uI��SŻ(���+�
�٣䛁�i�֡�Vv̪�K�`�_�aKY��߱��&R�5K�8k��p%�y�֤���3�
�F*�ǫ�wj��A2[�/qF��R�E��󳼑�^�Q3�%8Z���mB�EY:zjk<г���۟g����/2�m�P���c3��Ø?um-d1{&�E��d�ax��x��Ŏ�������1U<R�b�]�q����쿍��Q�˦�w���E��y���T�)��d�A?Q��$3���X������˺+�+�>�(�x^-�z�G���v'4_}�ru[gD�B��znI,P��zV8.֑H,���Gύ;��r�~t�z�xzٖW��j}�6���r��0`�T=���f�:�PxSd5m��9��ԍ;@��Ү�#Z�c^��o��pi$\yf̍�w�t� ��易�Zx�A��
�rp��J��&�5 �S}��D|�BJ�!��o�e� 4���g?�+����4��$Բ������0� �8�є�l�&yo��S����ڠ'51,���a��t�=�02�S�j5_ل�+c���X��o��S��!.+����M�˶���7�q���K���j�"���j馤�&\Pd����U���pda��i�*@��g!�u"��XyC�2�/��q�l��Pef�GhX���/�kd���6`�7�͢Œ��Y�Nz��?�@�
D��\9�Ⱦ �9z�%�i���c<��wI~d�#��<�?6�% N�X�7W53�����p�����B9��ĳ㋞�X�fC��#�[��WWW���A��"i,��H}G�̮8a��Ϲ<�H��n�Q�t4RK��{2�*�_�I!�KGO�;h�vD}�"��Gf2t���|FZ7`C�4����`�i�(��������Oy/z�:-�E1z�����EK�x<�ݤL����P
!�-�˦�%��\��d?����%��.���8�^��~����I��� �yFTT����t<K�����4ևh���h��Z���b��(�������9-\[|D�k����Ⱥ���^�$��F)ZS�s�����w810.��R���<~h4�����u4=C51	`}TңV��T�Q_�{��z[�X|�D�wv3Ln5��浾��a�{�^_ys�P����(���J���u����.�hV1�jt6�eJ\і+l�h.�5ZG�E�v��2v�����>Q|�~�u�	�״I��kӵ+C ��3�	�'M���f9� p8�mA������{cW���帨��+�E���o�6�Lo�p�a�sҾ �<7�'W��A�B�XdXr�G����W6��8��n��G�(@�`Bj
y5�}�ҽkuS�ir�?�鴉� �u�����S3D7�,�k�� �>��C�Fk��Kv)5��h��'�˺E�l�v�?!�4y�`�d�D��A���`�!�#�i�ۘQ��?�v��BI�-H�B�M�ہ]�*n�n���e�KD���t���[O���`��c��!��DU�G(��G;]��r�q&$�?�n'+��Hŧ��(w�oH.`���I\7pé�[��k��w^�=�TZ1�?s���M�Q�����`���Ϝ�tK��j��f�aG��5������2�)?o"uB��Ԟ2���.�����y�����pJ�s�m�3�G�^�`^s�{�X�5�� 
��b���u S��X�]p�ָ˜�tN�J	�#�ٻ�[��X�c�Ih�E��8֛u�Y���c��
~�C�aO��M95)���m�(��[bRA���1Rf@X��9=�Z�X��$]y���-�S�zj{"���M6�O8ʂB��'����zWx;JȌD�S\�%WV~��sZ��z�\���"-�>!��f�����eBI��I����Ev��o-���B��� 3�I$ݓ�Pо܏h���M���\0]
m���]-S��Z��Ds�S�{��Qze:��{Dp��#Dn+���W���ṙe�str�Z-���/or�����LL)��u"P����aqf�E��h�������f"L`�	.���e�9zL�Iε�e~�g�=}�߹�Pyw%��FӜj
������G	�w�
6��<�p]�5m�����u��Lo�he��d.Ѵ���%X��(/��#����N��V$�y�|��_mm��s��rf{׈�_1\u#C2�y	!�tdre�S�J��)�^M&b6'|�|>�f�M[yA��J�;[ԮۡI.��NР	m���v�p�ƱHHw��Tt+4d>U,-M%�/��ZI�4lԱ�	~&���6�x����"�m.���̕��|��7\Ŵ���7b��q�4*1�����~"�^�A���q.k#}�: ���N��cB���kmyZ$tu���&�F�z"�����9�)w������+���u#\h2�o!�-�{��E�{c�֐��C��Y$"B�^�LJ鈒�{�]#�#��/���*샞�ΰ=�ǡ�DU�!�S���*&�4�l�oϹ�&�x��`���xʄ;$ˠ���5����:��?��'�;�����b8�Zܪ	�����5P�x���>D���*5�4�ò��������l­ZԜ���d�VW�P� !����Ӑ[Cg;��$�b`ר�j�ޠK�*[-�Qa���Q�I��өU� J|�x��D��'�z���U{��}���q�(�60�R�@�	�b����H��a{���]��Ym�)[~��8#����Z7�{yHV})��YK�8�M���Hַ����� ��a���i=Ŕk�aݙ�_-�3j��-���A�Ѹ�~xćN�F����XeƂ�,]�sh~��$���]N�M��Pڙ���/�i����CNL�(b���5���^)�Qap?v����ab�������ء��'ǭ�&��v����kv��&
aY�0d�6)Y|�Xٕ�m˺�{u��ܒUƦ��*i
�XGz�d��x�&jݳ�+�� �Q�vr�:(~+�����.����K��2��vqU��Y����3�B�}�čk��K)�48����Y\.��	�AE�(01��Pҿ��_�),暴X[��{����:4���;m&���8���n
5%¤��C/6��6�0O�f���@��L%Zl����}]������>��(��N���!�6�AÎ�0��7�
Ns:��9�!�蛵�sـ��3B�O�t5i�_����m?B��Pv��8ά�����h��H��@q�(I����I�2ټ��e�G�h.˺8��2z���,U�Զ��wR�Bf,�;U��^7!��h�@��?}9��`��h�G��!ع0?p��o�t!o�[������Glb�j�}]�[�3:9)z~����!g� �;�m�S� �a�z͒9�I�=Lim�s(���􂕀��t}�v�N'�I./>��fXC��lO�z�N��4	�>&hVrLĘ+��y��$l��݇b�!�rf�5<��!�?B}Іg�����.A�,pI�%q��㖲%� /���}�^���@Ͷ�{s����?���)?����uX)x��F*\�n+8RTY#�M�Mv _9.�1���j�蒨�r�����A���}�3��B}j��y���"NΊ�E���52ʪ��u�����U��b�d-��6i Ȗf[������}LM��g�'E�f�x��č����N�o���L74dB���q����n���4��E�����z��ċe���=[���2S�����E.��6���N�l|��c��ȠQ_������f���t53g#�����
0��J	J�� pذ�Á����=?*��C����h+К��$�^���-<:�gm�W&�\��LCԿ���H�yd�ۚ]#�a�x܄�uv@��o��3��B@�ok8�wT���!�E��Ce2��b���#Tr���@�$�C]��-xM'L�H]*�~jIC�Y���F��^T0u��]ھ���_�A���p��o=᨟dɹt!�/�z�2�`�b�8�9��,��em�"�Ӊ�?o6%`����e1j�	��]��}%cϤ�/]e��٣� +�H�ȶ�?�(���q�ZO��͚h{�Y��öx�ikɸ[ �p�P�9�7g��B����y����6�B{���O.H��E�����r*�tp�;^*�Z���ሿu2�ɇ
���c�Zs߃��t䆆�k�]h9�QZ�����ΐz��I��@�
Y�
Ya�Ɛ�T��3hb>�����x_ئ{��',�5��A�th_~3X�i`T������O�'���W�:o�0�S�ȶB.pR��o*2�a��<����Wk/]�L��d��1#�K�܀���U�Z*~G�Fr��<A��qq<���{yo���5����n����[�X�w- �C�&���_s�'UTǂa��_�0�
�͚��L��~�@��2� � #S�ʜ���T�A��ʱ�k{�oL�pUuԙA ��b�$����}b�P��5n����@�JJ�L��X"�f�R���_Le�d�D�0cF"W�d��G�������x������o� N���Z�6C?���C��/tYl,{h�O��=��w?C�8��=Ӳ���["H���y|�N]�O�k�2��zʧ	�̾���{�������6�F����p!�Sh�O�3(hܲb4Y����I¿�TN�u[��al�M�Qø ���*��u���z�x'>Y�%V���� i�F;��a��Wu�n����L�m�zzV��AO��sm��r���y
& �P�*���YNoЍ�9�%4�t��b�r��Nap8��b�٧�^ԗ���z��F�=>�!�ƅ��HP�9_Q�B��;� ���&f�����m+�"Q��Y.�z�A��Q���L��QX�[���n�P6 ��z����j�2V�&��L�׺�lC.��1����6���l4�wd,���xwF�y+�j^x��d�9{�ǆ�\t��nw��P��$X�@M�{�������Kl�Ag�P���RG��\=�d��U�%�+V�^b?W%���(�4>�E򃉶ha�%��Ys�U�/R-�x-�*�r���#�{���rC�w����e�,�5��C��S�G�7ٺ��h�+H���.��0�6-CC5��9F�bD�����+f���6�[$�[�~���od�,�4�*��64��:3�����G1�E�����Ef�0d�U��9l��H��)`
S������b���(Y�֩%XF��>�=��<�K�����Jq��L팈w�=��c)Sd9}O,X��ӝ��j�73�`�*���u(�:;<����<��w2�q)���J0��|E$9�o�K�4Ve�}Ʒ�*|w,���9v���|'�e2�X��H+���$/�:�툑`8�5�n���4��	�$�����+`e�7�ԩ���Il�1�:\���&O,���d���+A]� 4�zaF��?�d��v����zڴ��j`���!���%b���b63�(��k�Kҧ��oL0��E�%@�ݶ��"���Z�HQ#�[YlήD�����}CL�8~��d$�«ʓ�3,��	iﮇ��!V��DXf��(:���0C��S�p���	٘d�I�UWξ�����L�}�λ���ر����L�+�/ZM�#Bq¡S�'��2������2,P�a�e&_8�Y�0�^�V���:v�e~���WK'��R��nÈ��ο���6�lH�[�++�a�O~  ��V��F�KRц���	���W���sk�T�m�4'�}�3e��7�&��ͬm�-�T�Z�[�x8Kh�3����=u�jh�P�h*��$�c��4m�Ƶ_Ҟɺ@e�5#�e�2M��Q�e�'h�pr�, 0q���~���v�(��"'�X�����롿���k� ���o�`�P�%F���RK�����Lڐ����]���@Dk��<��c��;9�p��ūTC���b��X�*+�gR
�O`I�l$��E����VD����29A��>����[�sA�|�5��v��d����}�#2�mζ�[���k����+�ZW_��0L8�kDJ���1_S�0
Zp�X����qY��mq�(�X߾��.�W~=�x�K� \\و<�tkC�N!��$0Do����t��_3��>�U^М���"YuTC��#ʥd���QW�0��^4ǿ�>����ۊl?�Zi$��pC��|�h4�f�������J񠶈 a��}��+(|���U�~L��.�f�ʀ=���Š�\J�(/�=`� �2"�sXI��Z�o&#���9��[ɴϥ�7�b�u�ź�l{�=�g$���lS��9'�p*R���5� ��i<"G�ˋ�a��@���_1�F|4$��^W%�vX*f��1MD"�$��q�Ͽ�J~��I/M���E�7p.}E\���.42]Mh�vK� ���ċ�&�` ������3k�u�p�J�g\�mH_%}	��G�S`u��׿򧢋�R�SKk��(o�7�K`��WH�MI-ޘ�O-PȰCb��)]$�"������uܥCӴi�*�l�cvA�Rox*0������';h�E>?{m|Uu��|(H}K9��~A6w�����z��;���c12�W�tB&r$~���w9[�Ҿ�������|Y��t $�[�n�s�UO
˸��7�gy��<�U��z6v�)��ŵ�<���������+3�.��q�����	���|��KdE_5��j�t�w�T����m��_nں�,�+���� 8d��hH��#�I+h:�K,���
Kƒ�tj�����փe^x"4�i#��P^��4	�JQ�iJ� �'��=n������儺N�y[�EK��IL�)�����ј����$��S���Do�И��o��|G)���;�,��?	��\3��'j,mdS�(�Y�c�����)���eNj�u4�h(h_��:yrJs�4AC�j1E��0chq�J��F�Uo"�[8G����Ck9��vPO��gL��kAN7�Dj-(���J��v/7ST��W��0;�(�o�/
��_�ޏ����%��E�d�\[-�!`�B�f����# ���~
[E�:��C�rUm��2d��*�23� �^1���V�k�a����򊾆t���%�dts���[��Edx>�E�wr~��w0�fr�1� O5��~�L�z��7��䴃v F��F4��3��a�
M�����;��֬�Dζl�e<6���v�'Z:�x'��aJ�H� J�7�߶K���Ft=A�si�&�+5�=o�t�3�ٶk��_뗴L� �BfNN9�)-ℏ�T��C��{j�Mԇ�V�|12��h�@��<�&�n�i�,�Qi~'9Љ�7
���=,aO]�?%f�&���h,����^�i�P���>v��Ґ�º�f�y�ߤ1Ft4{}B}�?W���]P���K�C�T��뇢Ӷ��{�zS�Mt�����dH�b�qw��n������"~�3��AY�5��S�W��,#�ۮ��j��B��o)�s��%�}��I�.;�����gDl�e�OP�O0����N�����m�� ��~.��vih
Oq
;��d ����2����)_�Td~e?��^YTJ�\B�?:^+l}�v�+��e=�t9�\�d�HV�z�c��2�'ۛ��˭f���C��뉜�;ͻ%��FJ���L�.�X�#Ԧ0��Q+��\o��'�@�@�eT�������paJ:/,�7��P���I�ٛ��S�V�r��oTΚ9J�� ��V��k�0O*��/o۶��#��	}e �&�b���/�)?w��_jՙ�]A���ÃW�����D~��ώFy�m/K���Sf�qǃp
߁�#~ ��lË7��s��%~Wzft=G��U�[ZQR�#�����BTR���9�ߦ�X=k�H_x=���`9O4@��	�<���>�݃	�5)��=V����k���\�d��y�>�~���F�+�Հ+�Ò�g��I[�r��*4Ņ��&.U�}�3b�����B�&])�9K��<�������T��v��:�8��7#f����Ո��8�Ǐb�$�MTDW�fb��w�J�w�I�u�8���L�kI(16Ԩ�LIo�Ii�}1>�Cԉ±|�T���ۭh���5��a�u����1��rgMY@��S\"8�ؖ�ȇq��J��)%�F�����rJ�a���k�#��A��9"(�p�.oD ��8�\$�?�Y�s�f��:1����(�Ѣ�B*�r�Ɲ�V���x>_�T�����o�`{w�ԫ���󎨍x�G�c\9k��3R������gf Շ����\��u��Ne�=7z��U?��Wf�~�*��QG�C��%������/� f,�]�p�'x�D'y��e���0�����x�ikLvHP�`j���h�`��!�2uQEx�}zi@���0j�KG���?G�P�m�ꎤ&p)%����1�&�[wuB�z;�@�8F���g:w��¶�$KH�����O\p.��r��@��,�j41��%B�|�\ɡ� ��Y�c8t=��;�_2�y�8T�2�X��ڭ����q��l�Y����o�0�y|���v��M��i�
�M����2Z|�5�l(`+<���q��׈jHV����~��(�]T�us��^WCX����6�p�܌�B�o6H��kc��!B4�p�mT�U��g\咜���@�aE:�OI_�p�#�!*�K�š�[1L�l>'|]$��N���-�f�Oh�R5�B�͘jA�#?�L�H���~��W��g-��$�#���$��>J3�闈��^{���E�a逓�C_�
@]Btpw]̆"5�ʤc%��3(،c�:J�T����m0�{���[��R�x���N���|d ���k�lǫ�a��J�髸��� �>��ss ����Ty��=0���k�؏���}J�e�z?�hv�H\1�e"Fe_'�9f�6,������6��$�o�	&�q��<T��#1UQ�v�]o�,`�n���D�����k)v�g7��c}�%�w�o��/��gǓ^.~�$��ף�2��f~]�$�o):o�Pܦ-})�eٍ��Iǟ#��G�t�������MF�b���]	
GT��T-����
ݜzx�(RH��s�*��^l��_lc#qr �u4�u�O��YOSe�`�N*��ǲ�d7����a�kH@?U�'�٫q���D�����.�\w�#������ᳯ[���G��?�����3#��#>��u+RҺB���$��v�:K��Xa�T�_�ymS(\�F��8A�sF�@�,��IP�� �he��s���O,o�#�4=����,��7�ǫR�I@��q�ґ�&�D�|jjRYs���N$������r֩�P`a*�1�q���ށ�^<"��9v�ZC�
�BHJ���tC+x�@J �%�2sa���H��GS��(�P��ĳ�b*+��C ��r���K��\�L��a�Tz%��O�%NE0����mJb{ ���;���'�A=��p�D�&pU�*H��KH;�B���Y���ݮ����8Y7�V�����߼`z1ԇ�W�h���{~�Lx��zI]��@
���k�.�vWN9�a�w��__���v̡Ma�0���h�6c��a�<�`Մ���Y4I�I�ˬ�c]��Y�e���`k[UZ�Ұ�-7�|�-N�|�iA�<Oe����i�����2/g� ! �@�x5rq=He�G��T���Q���;[0���7�77A?�a�:L]"� O�G4�p1��1KIs4!��������y&̋pV���ҥ��:���D������������|9�(���{�N��s���C"�z$T���5S�f�(�^��c)�I5�4���>����_�u��C��l�2\9�����P!�q� H�W����1k��hu�t��BW/�˒M������z�A����D ɓ>n�Վ^��1����4t �(�9��W|�wl�_���b����\,8���'�>:kjB�iq��=�n'<S�Y3O՝9�e���F�����ij��b�����gm�\�MwJ�<�y2zVB����C�����V9`:@�an����#���ǡ�%�u����z�ݹ)�Û��h�Ò���sK'���g�� ���M���y�yI�]�WkB�g�%���z�6{16��[
�������%�^ȝ5x�:)�SO��q��)��h�2M&Uץ��q��v��L�tu$��x��T�+j��������άA&fVw��u;��$Q2#T&���}�G<p++=>��g*K�ȯ�$6��򣖞��# (a�v���W��pné׀��~$I�>����=SE�vȾ���`FЯ*n���p��3�@�e�L��7���q� 5��`%�EE	����$�~�{9G�y$���\`��_��CT�?�ʖ�p�'����Jj>_ Q�`�Y�Y}�ϋ�8)s7�)ݯ�a:]?�^C?��wD�~��%E:����y*��ˣ~�.�;�B��-��&�Q�� ��!���v�4�pT�!ń��6X�p��ђ=�<�d�����,Ρ�B
h��?���ITbK�T3d� Z�Xl�d��s��5���O�DBv���P��LZ�H�<�Ft�N�K^��=ˡj̦�7K�	՗sx���<�xC��CH���o� G�\X�����ҡ��ܫ��"ZG�n�7F�rfj��?��1�� i�<�yB!�q�#[Zm�[��� �R#i��	��{U[.gbO@M�Z�OZjn��Mі���-���6Kں�L4�po�o��U�`��@��Аh1�+�N�4/��c�'Q�8T$���Kf:�lB��uҨ)G-��$v��ף�!�+�Z�_��8��T�і3IftST*�2F�{���[2 \]�
��~����?.'`�KԘ����{�_T\����(IG���T @��Z [��53�.{�����j3[1t$/�i;p�%�S�S
��D�M��=n�*�c�(�����1sg�|.�H߯X���cy��[=��ص��)C
}�`!��e�F�j��v�]S�?0PR���y�V,�0�X+����՞�yu��)�6���W���|n?��힧�y���!�g������F�Cp��|;>d�"3�j���o��K'��yE����g�\����UU���w�{��� ��^�@�up�g���hϹx�R���jGG4|0�@�
iv�F׼�!��AS�F�K��������W����ۂ`�	�4�o��@�O�Lr
��V�?G��Ղ���WBw� Ј�l
}����8J�I�b�!)icqq'��L�q$2�5�N��8RX�bm�����;s���f�be�R׎��wY���`� i`L;W��?�e���J6߰����J���q�w�Y�$��'�-�����E�z㪓����7��� .bYV�f��?�g�y+�y�B�=�P��������΅��n
��3��<��'!I��X��_Ө��g��+�H�rp.��s�3�r2r�U4�9.>�(���R
�z;��>����%A�����!��j��,�ͫ��1�6̧�	c��jSA�;	��y�:������|J�x��Tf�#(gY� ���ȿ���A�L������w_�*��d�]�4 _�(J����~[<wq�Ao�ٌ�P��N^������G�QYr�TM�W(B�w_����Sl�OQ�DJ�Ӳ*�48����B}�-�zs:��Md��_��u�|�jY&���g׼�̼��؅1Uj��Vc��@L� j[�G�8��XǯLz�s��E���������䱈,&�P����.��&�R�vu�=��bD�0�-���ɖ�ކ��Y1��'�%*n��������5�dČ|�����^���̙���eLG��c�NW>����
L���C?=H��2L�Mt�,�Pde�3�˲���M��� ����eoP��5B�-��j|(����(�]F���{x���|�$��na���c�w4�C&��3�qd�<&��h�įM�$�M�9�ĩ ����E7m�^��-�Ŋy+_C��߶�W�8I�������D���;-f���
�[��;zF{�cN�_�Y�&�07��ry�K�,>��� �le���O	O3:/����K��yor���s@���<0���iG���ؒ\�G�ʡ�?�_��jԷT9�gySM�ԍ�TԖP'�sA���Qwh���j�\E������KpM�ֻ��ے�~L�׫
��Nh��U`˕�$ûIҮ��x���)��oI���,�����ھ��%ZK���dFf�MYՄ�2�$=0�ݼ��V������q�vZSð�Yq̸�O��M����YhM����DF���r�CC�P�eo� U���z8��ڇh\��$	~��h���.<��S2F/��\��h+K�gL����2O�n��&�'IC���R'��S�cM W����bz�(_��.��~�A�S;OV�Tcw�7���!�GpqO4�X֕�$k���"�e�,Ҳ��R+��
�ik+�� �_�FW:Z[�7������xO ��t�Fh-�s��5�ݏm��S�ۚ�^�.|�;0���Ўh?�?�g�=�I5P��#�~bN8r	�!�Z�_="v���6K��xM���J���e�Ő�k�v�� �2�zg��cq����2�Z�p{6	�/V�Πi '�g 2i� ���e�C����Dw�u����.���T�_+��1pE��Ik{K��_0��$��!/��x�y���?��A��$^�-@Q��3(e�4[��i���?�M���U�x�q��( 7J�S����x�/	�تB��7��\/�K蔏�8�u��R�T�R#�3DD�8_�o
\C�
���\�/�~]A�����s��	�������-fPQH��X�q�R����eU�,�=�H��9�Sg�vfT[J�|#J�`|��
F�OCh�
���Ԯ�Ȟ��-�--�SW/���|@h�l5��A�'�3�FI��K J���˵hF�����j��L�� �h�l��#E�h�i����3/Nb��{(����v@]a�F+2χ+3�z�������9k�:�������B"��)���w]6�w�{���Z�����CzH�e7��0��E���B�tˠ�TTT��\Rm�~+b5���2H�F ,����\�X��^z�9������2MA轣��d=�`a�v�Y��ۈt(8ɋ9�'�7��~H�Qp�w����Fh���HF���7��΋^& �ey�2��;�8��8Vu6�vb��K5eu�6e����N�|�=&�R�o�ϭ�%�h�����G��o**o_@�t�i���`�5$��U�`�X>.T�?h�2X��8��^��<X�Sj �9�/����$x��S;Q&�(nmg��O�mǲќ��C�C�UQ�BI��!�f؉�M��>�*3y�/���9������Ԥ$���l�wE�K�~\��Y���&F$&�~X�w��N�b�Ƚg���W�L��9�:T��<�P4�d;PH��W=�7z��I�� C��+��~T{]���^���ٸ�"�ES��A�O��K'����;gzu��� �׸��#9"����C�)AC.oMJ��/H�҃��)o�n15�����}�~�!8��KZ���3FL�ص����;?�_�|�qowXV7r�j��ʲ#����,�~� ����DDW����g�芝�-/j�xg2�ͼ�FQ���Ex���L��"(/��F�k.%��p cA�9�����yb�2�c�H�%i	���`,�Z����]�O����w�G�5�|X�xz(�b#�؍ⵑ�ZWzL����	)�~�7E+�ʝ?�䌴�F޷���,�Sd�27�����9��'�vВ�b}4Hdu��x����R<7w?��t���&,si,����v�����2�\�w�sO�bT�s����B�]�!�UX=���YE2l�Ņsi����!��8��M�3����@mAM�NT}��G@;�I|����}��$!Tc�?5�Y�?*Ey4��{cr	8<��З� ��xF�=����t�xx��C�É��aͶM20(%��n�������j�ǿA����F�k8~?�#������GJ���P�@�M���k7��'�/jq�eϗ9*�av��t�q����P��{�h���}	�8�ij�����$��rL>�	l�3uO�W]7~���+�aJ��^fc�/�
 	�n2۲��ɿ�ƾ�@�f�c��KgY#��W����ȼ�B.j�Hy��,�C����B�� _�$Y$��{�0���q�K},�&]T��F Sg��҃����]��'޸a2^�0vͬ�\��a��q�#��#���e.ߵ���&dlƼ`$��"��\m淟����G_�:��1!�V��P��2(\�Ν|���xDG����_�u��ɋ��#B	B��6;�.2�v�v�OY�{I�\1{_Y6
uI����B9�hO�Kz����;~?��B�P�23��5Z���%���������/����)�f����E=̩���F���	�Z���P���: �^��J��T�r���w��K�W�H�_���m�߼�NU��-;P�=h?O����0D�E%��N{�~�S�h�I����y��Y`����U?6uUt|h~��@�ؽ���||�F([��VW.�@,��T�Y�kx�]����\+�3�2,�0��C�-��9��B�����\�|���zU�Za:�nܚ��(��MT5��d��✠��AY���6�v"����k��:t�Y�-�O�����?��j��>��СÈݮ�h��� �W�u:�vs[-{�;��[�R)h�j������S9���`��Q����{�����U�m�	�����&7��}�q޸q��.���4]WqI��O�:J�;�!A���V��EM�l�{�����$�Oe�-�Uщ��@ߡlW���[$�H�R�����ZvS�x��ʺ_a]�����ӱ�+�$��솨O)�ť�M�����F���%q
2w�v�[&��kx�l����%B����0�8�YȢ��w3{I*�[ac�������qfB:kaCL[�QJՂi�}��=�:%%�ІH�d�$�:�����6��,��֋���[�p���#����ws�_�!oc�L�$�~.J���Di�+���z�(�ou�������7;G�?vˎ��XD��������D�GpLP��Kg{Dt�6���b���.r��^��V�;Z�#&F��eP�z����<$_Y� Ud2��'��F��$"6u�/9`�[��K��⎣p[�u?�r�ӭ|�	��7X��y�(���~= #L���d�J��jwT��hFje�n��Mk��''W�M[�{̄��`������ݞ�0J�0a�<�g�Z�S����V��_U����,"���/r����=y���a�x�UHJuwo:RW�+K8����%��� pѰ�Lx�X�	�7�%T��{]�6�	jq�]��1�[�(���Kk4m+�_
�ɖ��d��7;O�y}��Ur�]����z����O�/��d뻹2'�=?�����ߕy����ֶ+������6�2�]u�1��.y������x� zJƃ'��#��%��c�Z;��s��g��O8��M�=2	�&X�z�d��v[b�E��n��3}e� +��ވ`�3�޵x���kY�F�y'b�X��"�� ��m*�/r@B?�����bm+n�d��df��4���!Ą]D�O���� ��X�侄e�L�y�g������9J�
d��۬l�j!��X�z�#"h�,�̥�&����ծ\5�{��i�Q=*�;�Ѩ�5����$t�H΋�x�����1i�_��N���"���HFH|�V�ssmkŭI'#� ��}�+6�b��2k��疜��8g�3�*L��^��WR�_1so>h6�����5�Á�ߟW�)��{>���]��H�lݮ"��}Љd���~���E�Q�V��F�l�vW�&w��.Wdz�>���:�q�=�����W+�1�M:���r1]ᒢ*��3G�f�z�0+��ʞRj���(��oD��	+��l�(R&�'n����G�x�ln:p��Wi��1'lϕr@��s٢U��\hOA�ki�'4j�ʬ%VS����P!h�ʸ�3���l�%)�h��V�\���RA�gBQ�����R� P�$�Zt%Ц������ݩvIl��}�L/�)�?�1�>���QaP��;(�̽�6��u*�
"d`"P�yf������^6Ɍ~Au؏M%�73f{��f�vvq9���p\��侷��Jox���'��y��	�ښxy&gہ�IN�	z밇�ƛL o,�
�k��$q4�BC�:�l�����Z�O��.q�a����c�*z�`=�����tZ:�P�W�g�9BY-���z۔4)��bl*�O&����2�S?�쀹i�S�\M�Aqc�H'��P�īWb� ��龜R�4�/�i��hBZ�d��@�$��{��p���O ��K+���tJ8w�5Uw�?a�����v*<vbi�W�a��^�hDN���}/1�,��ק��Ͼ�\zK�Z�B��(R���y,f��\2㍐SoXC�7O|�"��-�q�a2
�0C;6�������`S�{n@���y�P� �A5�d�����Ͱ�)�eE_��5��	49#�;� c�d��=�6�ՕG����p��gS���}�ͦ���%3�7��V��=IL���(oC
���nW6�c	9��Pr�l�p����8c�9��U%+p��'e~��T��ɽ���4�a���2���C�U[���h,�eb�&���0T\���2{Y�ul?�ƅ��=�ڝ��K�x�Jͧ�FÐG�p�YD�ul�qd(��o\��H-��ؿb��Tܪ��Y��iQ~�VC�k�^�ϛ� �?����0T��e�|���@�j�	�YI �Q����]�<��?�$��"�*uI�Ql�dU��Ly]'�?�Q�nW�ȄjW#��S4��X������Q�̯���-b�v�� ��b�l;N����M4M݆i��5�K�O0 ̮ �Ùɡς*�8�o�!BT�x+�J�Mf�a&��
8����,��E�GZ�y[o��O�T�v���w@�՗�����,s ��4�����'8cxBK+���tPh�"�U��4$f���ʹ2���X�;D��>1+��@]Jg�0ɾ?l[1����!T<�|�Ɂ�3Y�����^��=Cr�9��Rm�� ��kP��p]���5+����A���Y[0�9e��������6%kO�/�2l�mD_O�m�r��Fj6NVy5�����'�$�����^�٤-��V���݊��ݩ�J'g�=X5����j��X���4�"�]zV&j)'Z4��6V�`��>ѵ����.X�\D��a���Yo�$����^�Ǒ�z�]�v����f���W"EU�uKa��%:)���쐤RS��D���}�r@�	M�@"ʩ��S��I�CԞ�~GB&�j�~u�X���~l�~^�NO��wj��o�^RJk1'���:��i�rk×B<\�z���n�Hx��Kn��k\*�ųDe���<����Īu�.��UOD���CP*^}��=�Y�R`:+Tb'��,���(b�+���mJ��?.1�`�b=ۍj�V&6�Wȏw\�n럺��JFĠ��^#o�!���]�x��y\� m��-����)q��\���X��#�"�H���?���$#~:�I�s���@�����Mfj
�r�������;4�#ۜ��m��@4�۶��H�x��@�@ubɠ�sm�g^>�D����5Vm� ����3������θ��~��)���*�`����g��x��T���ה�7N!��	�о0��͊�D���5�C+RE?�|P��}��&2�4�������0��A��(')#�M�T�}����t�i/�b�,�z����B{6+N��e�"���Q'�'j��Uj��ٟ4�fÈ�j�;�bD���wP��⦗�D(@�м�#��x���v��{
v� Ü(3N$C\��R7�J��Ӯ�}��6�G��Q��@�
�겨�;x�dF����qL���J�;d����N��Wq0`r[�c3v����Zq���@�m͚�V�w����>���90�\�.'���A��Â�΄jP��;\c����+�����&u�ɬ��/�ia-�� �g���r��`������Ձ�O���㥿~g�x�
8��u(7�ڠ�H��Te�F:v��[l�YQ�K啛�:K�̂��*hBld�`-c�YW�{�7.:�Tk}ڏ���!F�r����`�O�<�z2��(5�����5:ЋB]o�ј	����18�S����B�������OL�[�hMp��?���ѡ`�H2]�ڝ'OZ�&V�$J�����={�hJO�j,B�o��.JMU�̦!�k"&�����ɋ�V��ؾ�Z��wG�_�E�/x�y��Yl��p)5����ƫB�Ì+UiE��*�t��`�nl��F����n��z�oA���~�qb�B��pZ��)&|y��!cKM��~9Ϳ�ہg/}J+Nq�|���o2c��%[��|���z�T%q�{���A��ʁ�oZ���F���#���z��θҳZ���A�Z��n���p^����hV���đ�L�3iG�Y�0A�_�*hN�P^:�'bb���ILcw��%=�[�cߡ��iJ&����Oɡ]@\H�ϯ��_3G�O�H�4�7a&*��P9�@%n}D�Ip`-8�(���Q�4hj�������4���2s�'��#�b��^����!�P��cC��<��m�g�dۘ��ie��
�$'�So��!3V��?�H�.�R0#�i��U
�)I7��a~���zq�R<�E��È���}�`�= ޝR*��N��6l7eI�%C��	�z0b�������_�	b��
wخBZj	\b�9����rt��ͣ��m��<��|*��)6$�HGr)� ���Pr �scи�;j�b���OջPSn+;�=k�F,�~p1ړT�2�&�ףL�b^�*�G#�J���돐SO~if$��� ��>%�z�q4���&)uA�6ǉ;D������dD�i+a���$�kng=�I1wdtW���xn!��.8��l\-��=V:|0�u�����f�WBB=�d4{ѝ���"]\�)̬����.����_�B�$�&��S�,,?����:Z��[�@h��{nz.��8�cv�s�����/Ƭك��#��  �%$���M �U�I��J�Ҁ׌�2���+���٪�w���8����-��`�X���`'l �L���5!�3Q;An���ީ��"���F���bC�X��V����U�D`��?Z�NL��������U�}�<����j�WcV��ֲ�DO����K��9���Ry�F��k
��B%O8p�qp��V!x�+]�l���81���Ig���w�F�U�ʆZ+��S]��3漨�UM�2X A��;ZcK�����e��������r�3޿ʆ���Yl���v{�D\uS~�M��g���� St>AF�!����SS� ��z_�.X���1�`x�2��;%M��$)O&l��G ZA{R~3
�2&�8r��wYߍ�����-��Oh��