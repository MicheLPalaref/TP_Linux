��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z���$Gp̱`��@n}�D����\��D�]����x����@R�� D|�ط�8���V�����`kj��̢N3b��C~������L��A�T��c�l���~D�����ӘFy��P�1�ɂa̓��;R�30��T�B� �H�чk��ێ����ʧ[��S˛���|�fK�`�J �G9�]"�\���*Omm ykM�篨��'2pxmK�E@�W� JD�h����{ħ@�W���*Ck&��Y�/�*�CԔ�ۍ�U�jz���4͎� p�s���V7��קk�.���E��&d����%s�!�O�+��%m�����+���v֐x���n��?�x����f�Ɣi5]��kfE�K�v
N>���}��Q��=o��5�?�V%�~�%��3mA4�s�_��ށtl.�����D_�M���9�� �@ �`ؕ5YM�U��L�Ď��l�_NKˋ�$����j���q��~��h|���i�2�X_;���ʡ�!=f�׶~ֆX�)א3�Q4qp�/lfݠLHGMp0X�V�Ω�P1}X̖�j��S�Mq\Cd�BT�rk�F��N,��h�v����V�M�±�)��t��F90��ti�+����&k�Â��@��ڕ�h4��D�}��吿?���V��Sh�վ �x\��u�;�?BZ|N�Iwx5�s\4�E�^����$�+���o޿D� H9�_�+���G��/O�n�01�*��ߕ%Y�����Km|YzQ�K�v;����~���̷?�<X�~%�(��hGڂ��cd"?	����HÐ�7Hn��F�]�c��d���|�-E��d�e��:�
 tv#�#Q�'�o��v`�E{�}�V�b�V�7LOF?Z�;��x���"����ϣ�SM�G`L�N�����iԎϲ-|���B��c
�d�䰤��\��6b��#���A�K�O|䔮�Jnn������?]���0��ʷ�}�W�D�!�M�іc�!cR1�l�94\��W��W�|?�[ǵ��X�}F�����߂cU���F[ƍ��E�^\vZ�o6�Ew��WkȿuE}����:���`�!�dLTK��(�TۡzEoZ�X���ҰIN�܋�dꩥ��Q�3���]cd�
ē�,l�P~B$\�/�[I��h��)����i�gV�Qo��2���ķ�ƃV�8m����j�ݏ���޶��A5�f_88� ��A��H���%�tP� ��vϑ�C���6c�s�5��Qah�3 �rsR�k��x:Z�*�\z�����V@�i�Ce��l���<nM��pq��[�����-��*�+m�Me�H}*	�V�t����uɿ	Y��[��<��ꦛƤG����-g��#�F�d�ӝU� ���'�CT�ּ�u x�����/fa����>�!����ce`'�yF�Kyoe��f� J�4�a�O� �)؋�!�gB��
�����^3�ϼ�:yp��������1У�RM)� u�1׼�`�L�&�<�!}�1���4��܃�\hͭ�B���e��4�?�m*�������^���2o�Ӝ�ho)�8|���������V�y	�%�2\tRS�7�|r�'��P^vb��Q>�Y!�h�����@��*�[�ND����ƥH`�I����F�;w{��9q�ݮ�P��;�A�����3���v��M�wMZ�YC�ųK���������z�� -�@�)���l�y.	��O��B������G��0T����_�����?j��1|D�v����N�Z]�w:5�q�x�޼��1�9�	�[�p�q�4�Ѻ�U,\�`y��xK�M�x��,�'�l�����M�2��+�0�n{���C~��Uv=`�d"��2�Ȼ��'}p���éf���HwE��U�V����bm� :����\�_d/Eu�,��T^ړW�fcwj�r����욮���i�����uR���j�nK�ad�1b��=9�d�Z�1�u��6W�~�ZS�����1�������b>�
j������Q�w�khW[��-;#���c���6'�ӗu�x�L:�0:�+�;;�4�tH�"�߲�w�0�t�T(����7��%V	q���+���������B�ę̱�3��	F�l#��AZ����s)���h-��b�J�Kq�=�M��#�W���l�3�tS;�5��������j{�P�<�ָo���3$�z��[���չ�h����䧓DI��&uM��h	۰3s��NW�Г��r|�v6�t좪��T{M�l�O������)��2��l��ҹ�����a�Ȁ�����~C\� >Լ�?{T$��6�\=G����;�r'�Qj�^-�,Jl��w�i�7gc4�>9�f۲�"�L<�@=_���J���Ű.���A��2a�
��}�w�S�/�"�4��d� �*H��Z�@&\'��u��B����?w��Wь�=.6�=�ϼ�K�j_�Y&��ˡz$a�3�g�!9���n~�
�S��;NY��䃥6��x�ۜۮ��{�U���xPqYB�+�?投1����5��Hgi�0�o!�����T��<�R��Ϡ@ԯ��^�Y�M�;".�(����}��}�t�a ���i�dc��T��у��(~�r����K�eV�u|'5>��,يF�$�s�	�];Ic�'J�[~sCl�N#��<r���������\�Qx:���<3��6�W ch����c���
��I���K��S����
��].�!������&�;��/c���Gj�&j�$7����b�پ5^�p\N-��q$�m�VX�!ӈ�K��p�t�k+A_Ss�ա,Z�1���]��˭�f�	Pl��:QnSQ�V��⦡�^u����=2�]kC���^�2�&��	vC��+MM���s�Yy��"h�y5V��ά#�(1�jnN��X�n�!(}�_���Z��7f�[B%�:�5\w?4�L#Ĉ������ҥy�cr���P����T����*��ڛ�XN��`�@�P$m��ڹfca�k�����+i�A�%��n�5�q��<to�� &]���*|s�6�f}zh[�?\�Ƕ���N��Y����
ڎ4�1����M;p��Ԍܽ�Έ֩��Pn��G������D[��Yx�aT�/�����}'e���9u���xp��ѝ8��Ͳ�a�;v��;���Ҝ
�D'��|�C��m�8�z/0��a��N��>��A�68�e��=�]z�0保_Ѵ莠i�/�QG9�yQZ������^���������"���w܄��"+��lA���)����.�XB2��`i��Lɒ�,9��	nq�:�5���]:X�P�xݶ	bpJ��(ُ��4�Pd$��]k��]q��5Qli���I�+y$�5b#���>�`b�e����3A��O�>M�O1�Yߜ�q��ꦶx��+s\ŧ�L���l�U�CK$aB�ni��}��%��P{|�љN^��p�G�*ܳ�=ve�?h /�T�S(�U�3�MV4s�C�q30&H���)b�G����=`�|Y�ν4��k<��7�و`��~�3zkA��8q2�k��ⴖi+�9_��o&�tp#��8}���C�;�-�N� �1�P�\����}���D��x=u��ټ���AT��$㏲e�Q$���d"�/D�:��c�9%��W�3ǀ"i0
��)x�U����P��UA�S;�q���$������tk��s�^[�$i
��i	�K첽S���<��6[�����9���R�%�3������*�~}��CG)U�^YD�e���!��*�gO�t:��'�N�@�>��z�C@�vʭ~�V��0�{u����A:ô�����֦�A�]����������3�6��	��<�hY���mclҦ��icؐ���jG0��_��:���"t�Q��r����jo��P �@f��H|�m��"1
Fu�CkDvT�S-"����n���]7�v��Lc3�mx�m���«ݳE���
ʙ�~6�`�Ou~��s�gz��OŖ�������e���Ml9ik��gs��Q�]�̅(�~t�m�Ǭ���/�=�Od��Ķ�;�q[�ĜG�2����]��Pb|��
�<�v���(C����K���ME�B��O�W_K���)hRx�vG���q�~��%ٿ�nӍ���b��K�����2�-�Q��#bXgѡ}Mxo���ˌX�9��k�P��!��j�1�j<�@!��c���X��Ӝ�����zU6�����"C��Xf�RJ���a��|�:
����J��e<��ڜ_�R}-��}E�?�̋�^%�ѩT�@�7"���<h;�P[����-�����;.ı������l�t��3�O��%;p L�]ý�p&n47B�kt,$�VU�C�l����a%j��n|�Q%�G��M�|����;F�o�j
a	@AP��oU�∂`�S�[��Y�y�B�ji%|����)�.nLZ���3�G��۹`m�<x.�_�TWa-��.���D�����:@�,!'o�	�����f�|\54	-ehA�w��"t����f��k�0۫�����Qi%u�yV7��R�G��r:�����G��<����+:�,�M`Ko��)h�@�[�)͐�>��Yoݾ��S�5ߜ���W��M%�zn��-�^���z�.��#-N.���l�G˜fJ��V̉��B�hl�Y].��~,��x��4X�ɴ�d 6;����g�'�FrxTYr"�<Q���q�ĩa�K�z�ndT��KRx��BcS�_o����:���ER��n� ��n�46l��)ؼ�땿k=��s�:�����Q�{�-L��G����$QL�I�'_�8�ȷ��G6G���F>�w��4;�wc���j�dcD�B���,{k5�?.�9o��͋�_�1<4H�I�[�!g��S���U�c���." �P�ÂK�������=�4��Q�Ys��s������.F�-B*v��:�Tm����IZt#��C�����G$�������m<�%����@*��i�F�@�8/ز�Ӌ�9�A��P0M����Ke �c+��*��h�V�.�	vs&�6�H��K����m����wQ��.��q_����It�fKm�W�S���9iԾ���/q��7A�᤬	5��Is���b�
���<9mN�gŌ6^�'V�S7�U��_K�"�#�@��\��a�H�ޠ蜻QC2@��+����0��p�l��t
ા�p-�lXXW���%���n@���Q�ȃ�M�=E���J@C��Z��ɳO;ڤ9fݫ�TC�� An,��p���**�Z�n�7�9y���s&�1(��"��G��@���H D���c.�~G ��m&��8\����, d����IQ5H�"|����\m���q�&��*G���F���3�ߊ[`Ń��p36U�s�Aa.�I�hߝN�*�Gn��5?�x��X-y�Ƶz[k�f�C�R#�ȝg�X�b��/�\��x�f�*$τ�T���Z�z�4w�W.I�Y�r�ʊU��(�t[����O&��Z�Pho|���@)0�N0Y���4�0�=W(���⵲r��dB�˱����-��J! ��1_�I1wܷ�������VeC�mT�(�D�j���B"��O���Q���1�'#e4����P7EX���ԃ"�6.�)
n!H>�t4-|���b���e*Iؚ٢ѯ�7禜�~Q��}��}��P�'[t�S�c^�c'��i�I?�퇵��%Mw���DЪ�ԯ��3�Lo��ë�#^�<�g����x N����Oǥ����fS���\]�q�bڰh\��!ll��so����9Tە��q.�1	h���Ku��|�xi$�b����&�'��(��Q�z���'lv9�b�LO��32��7q⭴�y[tq�O6�{Y�%��2�P�N�Z+�L��
���"��MB���|�����|�'�.�*�����X����k���`-+	;1�,Vo��kV�X��b(�r���gKNt��$unb� �Y�@�YS
�b�*��Ғ[ʈk�Y���3�;��B�Ϟx�L��ᄂ)��\~��劢�;h�uC����B2��+���H,�2�8��=�:�L�לS��'J����\��^P=%uf�9���c\�d��QJJu{�д��\~�,_�L�f8�̈��~�u���	,��Bl%c��s#���K:u;�iP���>gp�#�Ȥ����?��6QY�C�B�O܏�H�U6���]Ņ�M�n�A�����M����j���נFޜ��-��cK�!�Z1Ė���B�{�%I���[r�26�D/��i���aP�q�u��+�TC��%^���u�MH�*�]��[�$O�f��^�E����]H>E�p�,,f'����;�|/,I�w�A5j�/����2T��o�8Y�Q`��EexM^^�����_PR�o[({�Y��.�k
:��UZKP�S>�|�.�"���r��U{�V�e��I9���C��?+X`���~�U�֞�_-6;�)��j,wt�p����@�FP�޻�M�z�����k��r�^Fn�aQC�f�O��!H�@a5 ���ʊS��������!B`���r��3!�
�9�:]OgT�aYnĀ݄�ttp;x�
��<W|?H������Ver���WINQ5$aP����C�2�Cq�M��sz�D
z�gGսp�4�|i���7��3QuG2�T�XS�}=��T|V%EX��k�8 ���L8j^3@U�;m����`/;���>�Wlm�g��F{�Iȅ�v�<������R"� 
���>��?I-ȶF9�R����!1���4�#�ܨikv�(I�s����B8��)�g\��T�Uv����:�/�k��m���s%�5��:V�����u݆�Յ0�DA�_��!�[�����F� ��EU��~�-���,j����ы����Цn����y6����O2(Xh�l1`���5/��Th�{��̕uB�ѯ$��U�u��#=N�+2Q̩-/ƣ�=>���ӳ�?��gL�8��+�B�"����wf�ϱ!"��D77��xk��8ǎ�"��Q�����xf�C�(��EHy�,5ر����ӻ��Ɇ�qu��l�;'~e/Z>�1���E�&rzE%<s�1�	HȻ)%bN��s��~�J�rJ�N�$p����*��B�pr���ͫ� H)?Tn�[t��b�3�9�X5wJ���T���qJ���q��9��y2�3�R�J��:N����z����\e�����0ng�������N�OԿ�#����i��Vs>���T+�mʏL��=���~�3�s~[�;v�Ay�%�o�ԝc��)�J�n�pVa�x^"�o�H�hӳ�>����"�Ż?�WۼFX:�(��K�oq�����Y!;�Ȟ��,�HS�_�)�j.��Y���A�a��r�-��Oc�h3a��b-�M�{�P֐�֧�~�hB�7ߣ�T�z��M@9�*ؐﺔ��gR�Ч%q'�A�c�5YQP4�D��і���Sv�q(,���F5Whq@���\�?�'�h+�N��ŏI��� ~8nz��)wU!���0��Յ�~iQ���NU}�r�@"Φ���B��Y(��0ǥ|u��m��FZ\����$��@K{��wE^@Y6/��J
@��4���P�a��Q�7]�B��I�6�K9�[�Q�z�%��H�KU-��8����u2��3=B]*��D7���3I�FO���W��8��������X��Y8�$���Y1�}��ݙ4N@�آV�Z-��Fnҿ�4��?�-Im��|����
+��.n{���q� n��&I3�;LE�e�(�a��0A¡(Sɩ/*�pC��8k�
����W'@h׸�!Ҳ����i��y���NWE�I��l-�A4<�E��'Q5녺@�i����;7�֌N���HLJ*.O����W�DV6q�0tY�s������n.%N����U���P�E���X)����#�������=�pu.�d�w%b���p����CCGJNs6^���+�b������GL���M���3���ڊ.F�}`���)'��T�<��L*!R8K��+h{e���A$&��)��W<���">ί��:�,ڥ;B����]g\�9�F+�4�Z�{E^z����Vn��[�9ߑ�V8L6�ֹ��|]:4�+���v&�W5is��eN�����<�����҈Y�Lcl4�^�jp���9����W.AQ0�*2���A��I��K��s�B澂읆��:�����}5���v�U�$�%	����I��s�� �b0p\-3�,�
G����/��U��Y� =�*�vȾ�qȦ=>i����zG��*n�y�iQ���kT��`։/��_h�IK7�D΢hmq�wYQ��r/����J9���|�8
XӅ��tN\�ߑ9�����`�H�����Ac�T{��t�����6�-��OB�P����\8м�R��2	�w2~Vi�W���h��fZ����T�q�8~��y�k
cR��lw�ӻS��Bm�o�����u�$�T�~L�����g��Ǚ�DG�Q�;1Q��@Tz���V�1�uK����!������W>����� @o'��q�Rk��oI�vN�8��2�M�7��F�� <�f U�#�qJ�o�<��8n��H�!�$�䎦#�V��%���GQ�h�A�-��jnܗ�n�,%��T��` �Μ|�̪�J[M�-2E�5c�w�3ݪ�0P�N���� Ϛ�L�V%�y�?�+�V�8�枤܇H�[y���k�T�eVaa%Ф<gHr��"�d�iL�Ck���4c�A�JQӮF5�h�o��q���o�/(����^T{	��m�X��eX��4��I�6�9Z+I�>���?e��/�O(@7�aw�Zק��)��6�7���{��O�5�2�d_ec�$���F�qK�C:��$<ˮR_�sahtVLR����L��nF�'D��.�7^RΤ�DvT�'��x��=rp@��W��������r��.րv��p��29�_���
/N���%�^�Uk�f>���^�{?Ć��$�Wg;AC�:JU��TB;jaxm^��E�v���2�L+�[lX?,U�'�v�b�+ϯ��w<i���F��+��GM��eI���lDbٳ1���%;":�r�:�^���aZ����_&�\gcy����V�U!�d��\���x���♤0 ��=:�B5���X�������0�w���a�!�0�p���$؏�[	���ӫg�윕x�'BN����]I��N��<A��!s����T�vD��^�w�k=�U�����
�Թ��a�FN�cKU�Ѡ���������
ł���|�n�>�b���s<!���F<7�Llt/p��=�/B�[ʭE�_D� �#�xI)`��$�ov�$H����rI��9ܱ��Hh%:�u9����u�-#�7�����+k�_�v��QpC�aՍ��nE���֎r�#L���ِ����74s�FRa����`p#FE��P� �������a��Y�VI�3~���P���yy�����){L��Gu�1w��E�b�>$�\��tE,���`��~uIn ��2���4&��k-ބ�|��̚�`�3Dh���(D����U���O�O��}�z������bʍ��bH�Y�U-&��:#�jmB[Z�`���e�3bSW�R���$���B&U����]�aa��%H��}k�+�*=>��V���l�	�蔞�����x�r��0�Y�p����p�?�¬��u��p���4wA;>�ԶD�����S9�O0yK*GRypr �>z6��\O�$�i�n��gj.���%��*-��Y&���i7T�n�4�8�$���I�D﹵=��i�|Gh�K�pQ���zS<�Wu����b�ā�Su�N0OVV�w͢�inh/,������øJ�^�)�zo�?��+�꫼L��/�g���������i}:��		���]�ˤ9���4�-�34�S�0 �稒��n�20k�} 8bcw��M��$��$q����D��%�z�-��!HWvJi����/�d�ߤ�-�M�>�F�����S� ��u3�-���5�Q���^�Ic��;�+�(���T�r������3uq��Κ"���M}�%t�Z�O�z������a���wj���J�$+��2��"��q���{8-R���_7�(��h���ry�\����+��+��/����M�Ĝ�Z���0yŠ�O�	�ݲ"�����n����+z�$�?�8��{W9�S:EE[Y6��.x�8�����#�Р�%�����ŧW*W���ģ�Y�
3�E�l�; ��er*A���+4� �l��R}�Sh9�&��-�(y�4���6��CV�|� �1z��ٟ��^^@ͯ�tN�ޏ��[����S�܀��@��';���	����X�����B�>0����N�D�	ъ�gnE��x�Ň��F[ecq$��7��zxP3,ꏬ)�K���!�-:�dC)<�Q�J��a�H7�V ���ȳ>��`����N��!a=���������䝋ޜީ�l�F�����q��{���߿M�tM��e9o΁�U�dB��n6̟�=���mO:N4�j�7���j�� �|EIձ��̛s>ɤeW>����R��s\{�{WO�٥q���?�~���	a7�q���zݸc�k����H9n�U����vA�Eo��d&����[�Pf̇!J���Rÿ��S�\l\�Y�d��~7�'f��z���|xڸ�;��f=�v3~�jiq�r*��H܄����'l�PQ���ةk,���`ہJ�MT��z�BMoA���%�NU & %��1�|���E,��������%������zd	����) 6h��D��GT��m�"���c����Y2���g�Wk���-q�H�w?U�ǐ1����@4��eq�8o��*���aёb��.r��=����ӯw�kf�ܗ^p���b�-�G�ᑢ���,v$�hb����,��1W1�hw��5�1Ӄ��j��϶N�4�%���5����_����V���-�F^��x^r��x�G��X����m���|�c�jt��}Dkay)��[n��QAȀ�Ǎ-����1�.��K짯�ڛ���;��	/�Y��e{�����H�F�I.�������@�}|׸
6R�>� LԬp)��_NJt��x9��m^��w�v-44T�g����ܮ�ҍ�5s�����B�Q7�f�)�?߀L��U-�n5�9X�1�Q���e�Y��U!b������9R�N�ﲘ(rw��>�(WG߾����g�dԀ8{��~��X�1��{'D�F~���仄b�kJ�8������䑪=�9͞�ZA���Ny*��)΋�z��t��`��!��߱�J���Y�Z��(�PHZŸ�r	R.ӡ^���v��]_B\J�${��δ�h�zWQ}�~#� y�Q}G�6��ZK�$rJW�N�'�X�ľNqw��Ic[_��.�BV������a���M�2���x���a �c��"��j0nPW#���&<��x%~�ČbAP�u#����T E�)�M%��������;�0�cH���k�e~o@�!���WLi�F�j=�iv޲_ ����D�4?�hc ����t�{���)?]7������.�Z��1�0��M4	$��gZ��t�w�ڻb�2s&�b@�/A�5�à;[��)z"n
���5 ��n�'��DG��|��ls$^>�����oA_^Dq&h�����3��o� �6�!/��NEBi�]=m�>4��I�~r��5O�r�4���;����ll��G~Z�y#��)&Z�S���H�$֊$�MS��>}_�޽��r<��Le��˝�~�Ӯ�Q
O9��扴]��M���h��`�6���n}-=����O�Nm���&��ٿY>�l��H�p"���ő��e��B6����O�S`O7i��a�Wݏ b"RA|D��Ҫ����Fu�qKbdv��E�p�w�>�-�`��ҿ�K���t!�z�~�\l5{��5X<^*�鐜`�-�ߗ�����蜟�,�XVS���1�c�B5��8r�+���s��X�a�xZ\�8�2�m� ���<���c��������)����`�t&�ȟN+(���o{I�{G׳�ړ�V��x�F0[	{��� f����q1��|��/\��s���A��(��&�?K��䫺E��O��6���B���fq�̀�l&�9r�Eif'��̓3|+T%r�֏)����f�E٠%<���qʧ~GF\~1l>(��6��8(C>*�x�p�����Kే��a��Qi��߿v Rp?-|ere��.C������81��e�e�q��y孼��9�_I�cX�<(�����ɭ��1���A+i�^�h{I��+�s�h�}��6����S/#Ͼ[z�+D&����r����w���[�i,�w�����ݚU�[<O�r ��`����"�\��R\���ʌ��� �qȬ�A�Ӿ��k�;
f�ږP/�k��/'��Y,�����s�Z*	J��	�ppd�x�{1y^��?9�O8�����>c�Hg��Ntƻ�k��z��d�P�\
	�n���`��P�L������ó�- ���أu%��/+�ܼh�ը�.�jɞ����.��R��R�7n���h�h�3��-(ZHc�/�l����eII�S4�#,�`���9�+Ѥ�q��`��y�5g��oO��X���������i���\�eK��mvv�pz�;��ބ�(G��eK��m34�[A����)�����w�{�eGCB�%����r!��Ԥ�/#�1�*�A����A��z���ʃĔ�WL1���b&�������ħ��'H���$���.u�R����.�#�Vs��p\�׻�J���ˡ��9�z,�R��R�����ˠX���2dWw��6�����^4A �5��e��a;�^�o<�R2:	OZ�@�<�^�p|�E����a$�]�����j5�W��#h�:�H��k��>W$1`�*7ڏc���n�����HS	�U��Q>Z'�Ci�e��%W�l1cw(`r�gsIM�]��Yn���:슍w�~n�G��~��V~�
��_�UC[Sќ�qކ���ف����Fb�r1r@;��wC�t�.��!��-Uڟ|i����v�'��6�g�Q\��3)?�o@%
�S�Py�Y�A��n�p6��d��謌��)��Ѳh�-���o�-js�\������)$�	GQ*��1ե���h7_Yx&�AB���.�p)��h��}
����5e+Š�G��qr����gC�p�o��x�1@�����B!kn�cAB�Z&֟���qҦ��]f���#&���c�|P�_�O����,���p���;�y�s.�(�~ۖ�k��4I��v��qh.���銪������pWP����1f���7i+�sw�D����6q�O񨺰�IgV���m+lC��E�
�D�����.�׉<�)�y���'N0�椮��R�w�
hw�ݫ��ھu�Q�
��Ʀ�"_��� M�2���~�6�AF��R
z1����rr�u,�.;�ԧAz���������/1O@g��Lz����º��O�)4�T�żΫ�j,n�9�${ ~gr?�U.�6%�B�'����� Lp�]Ϙh���`��<h� ����9��|���@�
j�_�+}R�N�v�u�rt�QJ�R)�C+��Ӿj��7��=����ه�ƛ�ĸ�.�K��#�Q�vl�nIT������V�}�M5�T��z�8-;����A�ҷ�2��~p�KA��������$q�;:YC?bj�O
�a�B��c$b�Ff���bî�'!`Z{�E]?�p\�ݽ�����>
#r��b����!=�Lt�Бނ���U�A�� 넡�-�w�o�?_:��u��������/�,���m���?��LX��Q��S�O���yc������Q�y]��ݢ��x��"Rgν�˚E�A{BS~��03mƿs�X���t5 �Z��
8���jé`��E�G�;�	�CE�n�����#LD�ygDC�d(��
m�@K��us=c:;d怃�W�����ќ:�jp�7����~ă��_anw�}W�I%lm&�#�6�1��^8}�༅�^���"�*K?� "N�a[C�?��9�xQ��0\}H�J�����������
����ҝ���M�e�e'�U����=��Dj^R\��v�=ؕ�-�G���~Wiw��==�ֻ~�q{7Q�	i��H���u�ި�)�-MO�2P��L=��l�����ң�z|�P��������I�gL�ΰ�Ќ�i1���Q��XQ����h�o9�v>f�;�6����xrGr�L%�`��dEaN�k$bj2�՞�U�ӧ��h��"�� �����p�ı(��<dIPY��a�}���m����J'�w���#�DO�z9M/tVl��K��N囝��T<5MSigq �����r�D9��8K��d@q����W�D3w�4d`��/z&sTqs(��#�"��r��E��Aޑ(a�a���rő���_ey!��9�}^�Q-���S0��2��F��@�L#�+7L
���9h��T;�t�� ^�
HlE��I��}յvuxDB@�m`�Rn\���~J�W�YN��m61����b�o��<܆*Vx~�Ȁ���g�l�R%�B���ٳ��Z�dh��I�F��b��J�-�����i@8�ы��%Ԧ�[�i�=��^�����LyN����Q�
��nt��M%/7���z��>������F{�G���N�(-p4<�-�DH��Q�eu��kA���h0����+ �&�����v,�z���(�[�A���AS��Tm��/�$�n����s�4��{t{��b� � �*&m�H��2F�r�Li--#5�h!���P!�E�Y����F�7dDU��e�	9i���5D���s2aKSE�_=��=��֭�C���"k��P��������G>c>�X���C�Gi����a7i�v�g#(3��fߊ�/5���k@s�˖~���g�,NO���WY~0�ԙRU������(��"��:+���u��=f���� �l�lV��p9b ��~����Nz���5^0��".��3@g��9�t���n�8�bD�z u��I�)~0=��H:&���A��X��]��E3Sۈ���D3�U�[�������&C���6��4�$�O4r�sG��w@��I�����10j��F�"����Ko�k\�_�� ������5�Ћ�a�Î%�Lc���@a�v]�$���Wj�1N;��c�f�����o4M� �@�V �[�ɱ|I���;4� �O��}-�h[l9 $��b�)����TI���Ği��U3?i��í�c�g�)CLi�mxx:�U�X�[j龚�;���xc	>C~��u�$>����_:�+Z�cPŃ���^��2�� �;��HA���H�L%�PE�Ɖ:H	�w_�+�����qĴa(�Z���D4�H���ҍ^'�>�K[�|�\E��55 7� ��V�7�^33���M)�qn��I���> 4H����PI2��ټ^��Gq��u�à����9#i��2F���n�]�	\��5ǃ�|FU�n�X-���n��;�vS�t��V8�v��'�[J������eo'G���sE�e^Q� ng�:�A@�����I�=n!��ȞJ�~��vJ]��0�y�>�)��q��}��kfc�����ں��Aq��P�Jk��o���w1�8k;���1L0�A��.�N��ۭVk�G�K@ÿ7KE�uF&�~1��T�tH��㊔�z��0�֥���w��s��V�&"�jM��oT�-2T�G����,D�~Ԧ(n����O(���d"G����7d"�)7'MU���w]i��QOS�7��5��(��	�#otaN{�.����z��;J^�������w��+��'���E��A���� �Ia��Sː�Ƃef����%u����;υm�f�CeڮE�yQq| X����1 5��n���w�%$!t�9r�xh�b�G܌:I`��X��F�>�e��L�Z~ ���l��y� QS���SF�-h��:�=�"����:��[��|q�8_�ȓ٭%w�a�nǗ<w�x��S2���ք���l2��T�HT:�ׇ/5�[#�x$XGZR/�H�QDV�۸�������0�vMk� ���Tr�3�D��9n�3ǁ�w_�[x߅܈��Z�<���BD�(3V��ޘ���w.y����4=�=B�9�Emi�\��g�$�7ڷ�K���1[��˹H�#a=�2�|�ܮ
�~���:-,`3�aG��{iΉ@	�Oޜt�+���,X�IU0�GEd�d�"����O�!�<G��2a����dT��;���͸�����!��
�Z���N3��2Տ��`�f��v�B��m��?A������3	��줳�r�q�Q�T/C�^myS2?�в��ی��7gF"�(����[�p O����:����LI>dD$������m7��l(��p+%�߿;��07�%ǄY7�^-��פ0At͝{��<��	��R�T�r�z�Bk�V���K�����E�ޕ�s��7�ѡѸ�m�ɪ%��f	�9��|�f��|��O%��W��,���.}����Zq� �`���y�쟟��!Z�{m_*�}X�|0ų �?~�T.���r�1��r��8��K�ܦ�W���.�P�y'�p-��k�����;�I�$��(�@�*"�����&_I��WI@U�g�f|�I�!���,^�(А� ��2�p���pn؟e�b�m���� ���l7%P�q53���4;�t�y)�-�:������m��:�kVV����vJ?��9���	S�N��z���e?N�$F�A���r�t��5W�h�"� ��ထU~�� h�p�����9$Ky����1�.�i#ښJZ�߀�άc�.��cƣ$慑�_�ʶI�O7�ˬ�GFb!�*v���הn�{A���6�2��W���%�VU�b¸�1%ѭzC�Ħؖ�GCx �e`c?����w�nXʦ�o<O���5�dEԬ�E.�%Y�%����#�v�񞷟N�ّd
�G���tr���Բ�_˻�w6)�����n%Xm��0�GcA�/d8��id-�ƿɋ{�`���zP1�Fڴ{���ܘ��.)ԏ��g��ԓ���L���M���xN�%QR�ܟAR�o��72l��⁽�:p�n�Rs��{�#b�����u0��繲@o�b#l*�V+����D�ӭ�%\�`��J���DR��"MTX�3�����t�JOt��q���t�QZ�,9�u�T��A����
#�e�[D���7'<�fT��7�y���r�B�F�h�U�X��`�˴9���6�w�Tc��$��$.��[�m�>ܩ��>[���NH���o�Ǹʟ�ƝQ/�����h��fz0�6{܎���.�}�eJ��Lg�Z�K�� �uӫ�(��z��G@n\���@p�Tc�;��_F�n��󑴤�N�X|�nh��XZo'9�z�7@w2��Er� ���.p8%�4B�I���PZ��x��V*y5y<��~~o�m��l�A��[�;>Dڏ:�O�C)������,�/��\jr͗X�ҳ�c�Iޛ�������ḭj.�ä�bB%�5|�(
/����8��	�y�sVؕ
&�7Pv5�R%i�鮀��\D��1go}�2xc�Jq�RÝ<X�J;�Z��b�p�V��Y�&g�H��`�u�3�k��MXVM�0�#j|�'�S�ܛ�r��G9^	�׾¬q��� �P��gO� �� ���o �\��G:�>1��y��噳�ؚ�iW��R�j�l=<�~�����դ*BN0����|��`�7�2�}��6�+@�-v�!��W���ά���+-�|	������|��P��+Q�z�pSYզ,��E��X�W����řB��-%��<��3��.�_o�m<�����dBs�慄� �Z�͙D����h<w�3��OL�{��,�}���^Y���Ҡ�t��f&hi�|滓5c��>��z�����t��`�,.�x��8�+X!�*�=iH�4��P(
�)�u�\��|'�a�m�͆:��܌���Ӈ���+�*�Y����K���R��	�G�>���.*i��w��y7�~�ƞ�iZF�;ŧw�ժ.�ڦ�sM����œc�E�������;��+|���\'����.��,��g.��I���3�k��n�T�J��̔���j3��Q���7���3�Xw���@|{���)���*�t�~���;��Մ}�0i^簗�,�9��Ry\çh�������1�f4��uf��s��pq��dE3Z��� �興}�Ks�z�n�����	�D&ݸ�( ~��7?��8|f����,5�w}F#�Aj7�4���
�K�p�f��'��:����9��ѹ:z��P�g��ӏ�_ [���J��$��A}�/�A��i�=��N�����^bUt!�ӻ���=^d�C����qQ�>D7��]���dI����G2�YI
�~��l��_�AW?D,f�����VR���#�_�������D�/�s���1hO���:���gX�rw_�Ӭ3���J�k\n��S�(1��1�%���&�B/�օ���:](��^�9�G4J#rd��p���D���n��M������{ ��¹�����0l�ҩV5��Zr������94�;ό�L�>�	V���o�k^c�[���:�����u'#]��

��o��xO������NY��x��nn�}6��G��D��?(v.����z��ow�����L�!᛭ՉM�Ǒ��Vcg��ꌁ��F�ǁ�ͩ���S�jޏ�o��nd�Q|��B���2�	�O�Dʁ�!/oN��G<��.8|��WVjn��$/��	 9)�;d�h|�N�� �Ȭ�a����p�NThA�_�T�Mㄫ3bќn��*�g2@��	���H#�����L(T�����Eg��i��`�S���E�>?W�,U�r����Ԡ�3��o���\[i��:���b�B��g���ɗM:�!d���m��nb/�Ɣަ� q��MF4���eA��%��~�/��$�k�(|s�;b}��80p�BfL%��g�+���+�j����D�o�k�܀��ʴp':��dc�}G����n��"8�V�8��bݎہ���Q�;���*F��=�s%ܲ�!�[���Q���9݆�2�T��������n�vV�4�5�	W�;�,����{�L��>C��C�M�I�vW飺>���ziqtMf�XF��n���*���*"kmO�1��g��c��4��0���?׺��H^o�I1�lf�zUη��?ho�FM;2Z�G_c����5+�|�`{Z#��~@M��z�xL�!��.N~@���Lj�T�]�6�׫@d��%G�)�bN�`���Ӧ��բ��),=L�Go}N"��u����u"�ئ���K�kEѭ�jǃ��Hڤ�� 1�)�k��^c������L3�p� Vѝ	!k���6���tQ�4;4�W�����,����W��W�
?
c)���b2 4�/��w;┺j������M�">��R�aM����e�V̆q){�����R%mko�L����v�.�vr�H�'��2���&�)��Jvspf��|��MU��L��wj%GQ_�\�%#����rʆ����s�
fs)�\�B�_<?�a���$��^�9b�l�&cb����E��vcq���Rc�Kl�B9��k(W��İՁ�U�t�����vpЂ�O���@����oX] �͵1@�Fp��-ֻ�w�v�������$-ӡ����S'K�aj-�+�ˌ#����G�?u�8-f���z�D����g!h?�P�kD	��%�(NR��n	ɱ6R�B�J���8�{i�g߃�pM6'e?�3H�\hu�!� $��I1�ʠ^��9M���S� k���p(*Jv�Cʻ�L%x��}��u����w<��&Z���|�q��!��+���B�J�.�� ��Y�Jf6O��L͇l�����ckS[y����)n��x<B�]���4��1o���c�b�+�������_P�b�)��a<�����#Drd��j&��K���pQ����IQ�i���B��e[��_nˊѺ�`��Ct^�ή��y�h�D���3� "L�s�?+����'���j�B�t5<ĭM8e[���-�8"ܣ�Az�R6���#�|`�F�5C(�?ΆUrd�g���M�u�`.�g�u1�F�?,�g�� �`a<�jݿQ9�4����ֻt�����`mY	H0��n.�h�Ն��J�Q��fRef,���{.���5q'<1�����8�m�f�m1-�JA8,�ʏ�BM�@tB�
�wϊN/�$�>�(��r,��*ď���B]�m&\��0�\%Cn��*r�7pWVKۭNU� ��s✬��H_s�ux��{5g���S{h���}AK���M��}!�Ğ�Br�>5E�d�E,	�WIT�A�_,�H8�����ۣ�D��$u���)U�V�c�lW
��l���Z�&Z%�Á"�Ay`���s�C&�{�Ϡ��joR¨�&�������}[i�M��؄�A'O���(xJ�_W��#����<6�
��E�F�Ԍ�b���+i�z��#��q�E�� �2�4�^�i�-h�;.d�5���ͭ=�Zj����Lr�컅j�[��;���P���^Q�q
^0&_���Ėz��'?�I�:mj��&�/�b蓕y/�F�����Fi�pU����O;�N�*�J��F��Cᶪ3ʁ��� �M�3��B���5�V&�@�a�	�?"�{�_2�0N�Q�R�B�QCA�'�}��S���Z�~��q0�rd({O�{}�Ȗ�<\ƅ6�?M��+����2�}O�~�io/Ba;^���'�wa'�(�:9;�v�����/��O��_�<h�)�����O�&�i�f����ǳ��bQ��/w���S�u)�(�e���=Ԑ-.К�d��3k�A1���ѻ��1�d��Q=��a��TeW�x�aWq:�FP��	��%=�]D�(^�a9+i��7�8�}3�����w��\��Um�h���~��-����C��n���<�Z03���Z��ͼ<���$<Yd����kE`B�o������R/8q�
�'���wɖ�)d���RY:MQ����@�!�#j[dm@���j~k�w=X~��oA{NB���]Ѻ:�h�V������W���N������#���EÉ���q!ik����IO��Î.��e���%�$&˛"��9��S�yF�ϝ=Q�ܦ�T��N�p��5}/�IH��ګ�6+�`�@�:��V92�Si3���Z�k��mt,\!_,΢�>����<E��z�E����D�ѡc"�����x��'��P�E�.ȩ�������X7ϯ��_�8�1�h[�Jv�'��S[�I�A�Ӻ���N&E�ߓٗ�Q��n�:�/:�]��P*�	�r���myN!N�vN��Wn��j�+���K��/����T>����FS4����9o��瘽ϛ{�D�Q'�^Z�I�Tb�z��N��p�������6L�Y�hr�m	��2�(��h�V�j���K���°�l�aj�$9�s+z��QR��Ԓ�X����� C͎���~�����3bW��g0��
�;����<5�1�뇾�|���H�st܌���wI�4B�s�f+���C/�p����E��i�v�������b��j�Zٕ�Z[&�S���P���Jqx���$����^O� {`�o��:��B�D�ބM��$�tx��Hh܉<ʽӋ��A3H���v[_���v��MA�sK�2߆���;讯��fa�&� �ɡ �Sx[[�El�Z�/@^1�W0	rΈ�U�����>T�+���Ӛ|���5(9A��W�Y!�]�@�A����3O�����ۀ�H�s��i��[����$�3Üvz����µ��ܜ�)" yFy�ՍȮ9<��v?ζGă�+�g�Վ��m�L��U���K;Ӱ4�o����㸶�\������x��gn!���UC��J�~keʯ�Wr�6�rG��]�Yj"dB�$T�����X#����j���xa��	Xm1~�c��۟�D�TOLu_8<ɾ|��O��K��Ne ɵ5߻����C�%��}/y�,���Q4@x�C���S���  B�����[��<-ǰȆGYߓc��&�v�#ο 4+'@;��af�����w��4p��-}�և�WI#qL��UR.�4B ��%U� i�7I�sj� �5�Ȝ�l�P;7�4�%�Iy5���AV=}\I'e�A"m�ҡK�#��s�ڰ��C6bȁ�%x{���KfX;��z:� $^�g���ƈ�4�].;hQJ���E��mbO ����?����(?ۈ����b8�n*l)��߭�E��g�wD;�i��H��8;2�9K�[IA<w��g,F�	�����a�1��ܞ��N\Wwq4<�c����ʸ�q �3�G�<��,K�
��]}���.�KN�&��s��	/���@q�%! ���$s��-!߅�%Z��Pߞ�Z��$2����(G$:�M�V���]�s7�D��|�s��a=�5N�<�,t3Qa�o��#���t���脱%!��h<���3KB.�R�5��<�,o$\Э�9��:�J�.3�3?��-�F�m0D�����WU%Ĉ�
P5�>��4{�F����l���%t��2�y��~N-�]�R��kr�Pހ�C$�*W.;���my���A*4�d��ʨ�)��*�[a��ܖ��Y�����jM�܌� ��Ϊ;�,:���X�m�L���ԍ'$�D�&>b��"��ԟ}",��gHy�'5WA�j囼|UF�|�I^����XF�|á�f5��{�:���󢃥��8�!'�5D��"6��=�BX&��+M�w��/��tg|��խR&�'�!�7�Ū��?Tn���Ҷ 4����[
���"%{d�B��.K������?M�'T
��ч��7���X�'4��X,ܗ\���)�wm��	�Ԫ��v�X�}J�?��� �{�~�J�]K�Ҷr0��1�R`h�{�!�#���'9����X�R��$wC�os�a���k��{�YU J�����u:���謖yRG�5.�b�r>�a	rs�\�/
y�V�6+��ƃ�ba0|/v� ��������]�<��c�`+�^��"Y=��O�)܀FM��_��>��*�h���֐�ھc����̸ګ�!�W�߳�����\
�{o�!��ꊤ-��Xf���x�	���[
�O�ْ�p��ii2�
Eh(©��y����k2�#<�/�p����v*�4&� p9�,�g���Y��Lվy���s�J�H���XOH�E8��L��c��Q�> }�ǜL�lr�y��dL�ҏ��s^�!����������9�#iu��0C,f���j�(�e� �.ې����^b��{<��'>6��'h��RP���uWn��{XY9�:����K�7�;��	{�3�,�ɴ̃OGn?�������̎�GCE�Ĕ%�e2�-m˟P"�v��k�H�6�VC3�1��Y�(�c���~�~��Ύo��Қʝ���.Bp?���(s弜����u�3��`nE	-Ѫ�B�7�g/<��$�ub�2ZxaK���%߅���6v�2k��+����-����]oc�<!�3�a���{j�A�� ��Z7O��q b�Fnk}��k�u��3I���U�vc �D��ՠ{H~��-�3�?�Ar�t;7ﲏ�yr4E��󫏫2�	�������IM-q��Z$�u-�gu��#�ٶX����+/��?����Ԇ�J3nYmn��R���ο�S��Qʶ�N�]l������̿`P�����A�Ȟ��}y���j��ص���晡a����+�Y�,�b��)�<�^�c���m�W�*��]�OU� ��m�3(�YV�����$.��P�w��Bf^n��%�[@�Y����4Y��щJN�@�'pq�l�`�"�[J�Q<���`�������üh&�,nF_6<yWcʸ@#�4���J_�j�.�il��O��5���� �5��"L��^��_N?_l�.�jm�&f�[�����V�,&�h2l�HZ��:��#�>����t��ʑO���1'����.:HF�å0|YpȞ=�y�MguG��~wFc��n�p� VF:��K���(���f�ԜQ�/��QD~�A�֨e��Nl�&�vg4SI�ܖ#{P�Y�@�iY���YO۴X�w9�ZbJdn�YU�����4��ȶ|�9k���Òͣ�[�pʧ�Kt8qp�6�2ʍ���ϕ�a�e�ă��j���4z��@�^�ٵo#��T
��ܓ"ʮ,V1�-�LyPBx�܆�mD��I��"�c�0L�Q������rʶ��%�V�	�G�����ո!N*
pT�]��5�#1GD(��_�A��k����L]��Vy0*���/��l�1�1���7d9�h��q�ϣy�?\���ݰ �]�Ԗ�΀Q���	��z�����SM�I1�(wL���ho�ߪH,O���u�Z� ����>^-���}%�g?)������k����xpCFp���$��[�<����={�J���̚�����K�C(��lXT�{I0�jO[^�,�fݪ�� �y�|��	K�>Aq��k�^Bz	c�ˡ�#\z���Y���E�8c�cpg5](֠-\Z�^&�,j��P��M��lye(�lC��Y]�[��T� ��m�X��Q��z9��r���O1��"���Nj?���S�\�F��㎖�����j��P�3)/��_1�D����C��er��A!{�-���(�@�*���L	DNh'=����R��=C����y�r�CG��`	��p�=�"��?ǉ /�X�j� ��u�p{��W\��������u5d
�b��q�'o?���Y�s;@��uE�E"�:%�De"����6�]
�c�j�kY�a�=a�U�	��,����=t��j����݆Z�-��y v<�������י�tTG�G#���[�&�jR�B��0�X���	�
��(g�9�M���W�=qyX�q��z����b񳟇?��`s�۸z� ������M{ˮӄ�L<�D~7UM��J�}��͞ZUf�}g�h�5Dg�K��^5�)Q��l��xg]�Z�p�=��pR��Nt�B��hgK�U�q���|�8�󷜆�Y��[���9�띷�Yf�����O��Q���~S���<2���Pn �f fNtx�GS��˕30�uϏ`}���5�?,IcW�q�~�K䈅��3��dЂ�ME=��
_�m������{rN�6R��!�b�YC�� ﱥ����c�H2b_
is³A>�eL����_�|?��{>��F-�V�>t(hr� �&J�q���0II�q�0�[C�L)�����V:�e���4Q�tpA�!\��|��ӱ��Kp�Vv,:Z�x�x@�R�e9�A�<��MF\�<ivD�x��h��|R��̖���-N��E�"Z������^�@�o��3�;k�ȟ%m��ε�x�7V�1*��\���N���F��#k��c�C��ӛ�L@ �>wfT�?0A��m����c��NNf�jio_��]T�b�����{tJ����=����1�7[L�Y�%��>c��5�(������#)~Ybe
v󩳓%�g��H���@?�v?n�0r�ī�v�C�.X��ƿ�3�d�ɿ蜛�+��i	��k҄��'f�����¯#�1�,���t.�����Z��c�G�$^L�b��V���Ma���R����28�llD �8W��`�7ʋE���w��~�������L����l�9����u啳�.Wwb��K��������o&��R}���#��xO�=e̪ȼ���Lp�z��/���ȿ�Rci-E%�^�(s$,�M�'��)M_�^9!o2��ü9q|���PA˲�[�K���i_�20����������G����W�">�^S���c�6e�$c�m���i�(�ERy�(NcvJ-�I��	b����d��L��{n�zi��%t#[ܐ���T��๫޼b$��E.Gj=��~{Z����J��ӧ�ڗ=�]4����ʬ�������-s$X�vk���aj�b������;�I^� ���ڋ�0�/�g?L�G��Ȝ:���#�g/�uDx霒A����^��ځy����d�?8������@�i�Uϔ��
��Q�nHk��m.0��F��.���w�Ѯm;:*l�ٷM�/Ou��L+'w���;���P����+�Z��^LaRum6Y:�ڀ�)�� 	�nΞ�Ry����z�h����d]Y�4�!i�\�9(���OҴ�7ǹ��\���E�����1r��&\2ʰ��}G�3]�Zt��0ŷ����� <q����:!8�=��b�V���ʎdE�2���8^
�e��������\����4J��R�MNP�3.�(�g�:���vn!|/�$7aD��I�-��=��El�4`��Jfj`�#�^��/qUL����z"���gA�x�o`���q�v<}��,������ �o`�!vm�����-��#` �hͯ憓���k�[u뙚��H�3���"A�U�Е[�����p��7	L����y;Y0TpEf|������o�͐�;�%���ta�=Ru���sÇ�2�Y��|Q�i����w³Q"���A����3J��?t��\e�.wU����k��T�PyPѻ��W�I�cO<ҝw&gX$��)�A����n���tEM4����v-8��~�v��*G9���l����G�Z�bȩ�(	q��@�Pjhn�QZ���C����K�_�u.��� :�F�n�]�Jg��Mqr��$�j#;�P~R���ߪ��ZI���O��g�Q$�WR֯w�%���0�9}�!"ޖ���Vf\���e0�gm��M�U���D�%a�a9���ت���˨,��UL�>ܦ,��~��y3PX���O@�S�C"��Z-36�!1����\20h*=?Y��>�RBa�@+��P�W+�p�wi���l�r�c{��6���<�Y�7�!�HBM��X|��brZ�Pχ���yH5�2�Q{,3\(�LO�&[�ogq!���|:��DDb~V��ƽ[���Tg�x��dD�+����(���ϡ2�|S�%�_b�\�b�������ؙA�?S��<0�TQ����sL7��
�6R��|фz(�sd;�pS}�q&���U�c	��!�!�M �ƥ��R;w�=�h^���I�}-� �Z�IN4�p ���>8�3u)��N��wG�8@�"e,+�͠��ndiɾ꺏S"����K�K�"��b�����Cb)�&ʆ*����\���.�&dx���F�#���1��вA5\7�����8'.hw�%@��樢���!޹p����7�>�C�b���G����y�}}������GRRo�K�
p�g5��q���-��nޮ8�7k?��kˉ���'ݾ��!�g������޵�P�/�-����<�o��ڭ���TeM��be�����MK�%A�������Q�54�vi��d��V͉���G6o�n�p����0̮(v|E���c���G�%_��� �x��stWh3(��58��2�g��hl�+��B3,@j�E�V�Dz:���/<UE���y\W�gIS�b5��އ`���|��=&ۙ�Џ��v��$0�ӑ,'�E��`'����O\A����kܸT�z�O�F��	Ti�t��e�e@�-�Q����6�?�o(TW�|�M-	^ȉ���������~\ts�y��"�b��������-Ԇ��Ƨ4����+��Hf��{-?�/���h�����Ǎ㏲���fP+�%0�w�2c�Y �Za>((�і�;@��ycGś��y��mÚ�s!��}��h��j�kXh�����#1-��[��r��x������6BL���i��v�hWK�8p.�����R�WA�A\�d(r\��)F�N�ZU�X]6�$*����K��0 �48���f&�F��b@�/�bA��'�&�JHȭ�;�qZ�<���FyE���������x^��ZPqI��^E��Å��9w޾���Z���������م�e�s�jd�O���0������VN�U_x7#�d�r�#"���A��m2%0@�Ly�L��j�1ZD������h�d<��O86���ѕ��2��cz�߽���=F4���
6�&��J�6��p�'���g�Js*�m6���9�P�X�d�te�s8;WB������[��W!o3� �=*����,�k#��Osd+;��(��i�L�Z\���k@�Ҿ���dRKJ��$������6�?}oG���g��	=>ĥ���|t������ץ�`�A�3l�h}E��^�{��6��R��-C���Z�P��?�hv�C���Z0#%�+�wB��d*��&տ
��J�z%�������f��%4z���{[/��ǎ'z�d��ƿ�Պpg�F�{��V~۞^jzJ]�����Id���Vy�^r�?K4X�GJ	��n8��)��?g�A�=�gz��|��OK��~%/�x������i���J�h����+�'"�v�T	~�����4����V�����[ ���e�SE����!@���Ml�n�+���"�o���*�~�첐�a����>k�h�>�3�EKC��c�������'u����K
������b���~�Q��b.j=��n4#x�"P�}M|ƸA��h����EP�1C�@4(@��o��8���x�ꙣd羶�w�f��r*����s� �e��Ըi8�)������O7 ��ž]6�+�_��A����2��6�=�໺�5�F��}{D��ݤC�.[:.m�����5[��.��C�n;C藵��S�����{���U�9i#7�0ci��q-SC�"��^�%��~��)������ep:�+<��b��~{�vڢ�2��Z�F��C��1YA� ���E�;��`2��_��fJ:�2��e�Q�s��ӹ��`Vy"v>�_��#�p���M��	�j7x�U^�"�9�PW>�cy� �1 k5����X����b#��y�q5�{Y��W�n��-Y�;��:��H-�~�.���I�OG��	*�E�c`�B��K8i������i(��tt��6���`]�I`X�NM3z���?8�%Ϟ����>�ou����پ�J�����Xe$�]b�5����/&��ă���^F����!�^a�G�dU*�^7���	l���/'!��˞��D�H� x.��{s�"�tln�+���f��_�:m�gx�B7:=ІQ$�o�8v*��\0����zl�:��p�ͳ�����ٚC���T9 �=Zu;��1� OG����k��%'?�
���ŉ�x�W���@�S�ID�3���Պ���a3NP)�v��N����q�,�1��e�������8�0��Z8�̈́�X���5MX�Xzm��A�*D�I���Z{U�@�F#0�y��bʹ�.��k�8�j�����So�*Ω4-D��x�b*%0���?�4������|�3��M��!]�����m��R� e�����*<�nM�T	q�e�c�.2����:�̑�E�6P$o ^&9ٗ24)�����An��-��7�a��A̗ӿ�Rҿ�y9�pW�ב�Ք�	m�D1P�`vLV�1VM-��?ӹ�O������BC�<�ARC�w�����<�����l��tH
�7`�F��daN��1Y8v�C�S$vw8����6!)O��$��<;���ƀ��ۅ��S��o`O�n!p�yE���$~�%�,j�x��^�u��3���SQ&H{Ci�e����-��n����E�q�������ia��F�l7�wHi��%�=	˦�_k.^&�:v��;=$��$�+��
��i��� �6	�eB�v��)�J�^t�B����������j�Kdd��Z,���ޛ͎�r��nٗ$��n�*W�F�,��Z� ���l ��X���ãxX�H9e�jM(��/|�H��b��^c)A�w��c���Z���[��k�֙֬���q�e��[���glY���r,�f�����w���fKH�'I�7�����6n �
ڵ�4�Vb�� �,������NI�(�V7lxT���b�dl�f�Ee�c��&��q\� Z=AwS�6���x��a�⽾��FO���
�׃|ЕC�^�jҰR72_޸	�jU��0�I���Y����oz�J�E�U�����([�C�f�E�tp�'$��U6�=O%$WV�ņ�n/֋=���j
�ce����x������A���Z$�a���V����0����*��9-l�5r�a�j�� @�M��9_$N�x w �����ոr�ƹ	���?W���I?�m;]���U���.%}�������N?�B��������c���m��A���|Xj�k�c�'��Or��PW6,��"ǀ���x�d��۶]k���aI6�t8����7Jc��3��n;�U���OUc�����%�l�" ��T���n��i�v�ߴw��(v�ø@I=��������tC�wQƐ,�s�X"=�s��I�^��9Xv�x�Nzӷ���D��-��FR���ڕM��s���`��ݝCm�.�5�s����4o�'\)x���S(*)�,�y
Gf���Jw�\�u��Ů���d��_�֛�m!P�$F2������x7*u��DXtT�LP��x��*$��[�<B�(���Y�n]��n%|�-������q��W*H��#ݮ���SU�\X+3���I8�A�K��ND�!��OX<a)�~?��E���!���&0jp��^*b
�&�*�Q��I������O�oO�xV��l���%��N��@;ů�݀��S�;i*h'z��:�7�˧�����7h�ϹKT����������L��������5<�����dHA������ܬ�^,���
����2�������9'Y%���(;����ۭ�+x?P�&KVC�zGH2P��A �A�9u�+l���HP	��neӣ��bɕ�K>Q��(�πU"���.���и =,�^f���Ž��9.�΄<k�)������Xz��K1�y��eV�-k|��I����ZPJ��J(����8�w��r�m�:V#r�)D�CC���Mc���kus�j���nL�Q���[���5����?��Ҫ~NC.�`�k;�`��Nهl��Rg�L�3vY�PðƎZ%wX��ҧUO'���g����2����C�o��[0�����A�U��C��j�VBY�&r��Tԏ��,o'��@M5�8�D����"�}t�.�Kvl@�յ�
�Q[�����1����}.�/֡�����{l:�u#R�P��
�F�u�<�D�N�uI�}��a[1<7u�E����#�4�(m� T�G%�;�8��;S�!Q�i8�ZlN~��/}3S/hc�Xז�c��s�����J�h��˯s�&�_�]�����Z�B�t�7�'����G���G�5�>X�e�p�Ȉ.s��U���ʘ��W����R�́G�|v]�8k��˴@�gm.M
k�xU��b�e�H�6W������)W�F�o{0�8�� ���6cgS�G)蠂�ObzW���x�����An��LdCC�A����Q��
W�o��:�?= �ڄ�?s�|.�V�?�8�b(f��@��0/I[�i~he�u�O��G�}jQ�;ɗ�
��v5z�e��.��R��
J4O#WX�BK�D�j���I��
�ʋ�d�I6�&c��e9A��w9��|V���@��/�}N��Jr���ބՐ�'��䓞D����Z����`��>qU�}������"_�����!xg��7�W�������+�U��}���d5kj�U^�0HB%��i&p�z���f�	�pv�0NL�`�8���Zr����>�	�*�Ũߞ���[ӭ%�|ld���;l��)�<�K�k.V���J�Pvp�2Boͦ`p�����s)GG��x��(������s3�M�,u\Ϩ�^$�;+QJK�fL�oľ4��K�p3��"�S�Il�
�k[��/h%r%=����B��O+5f!4�x��c�~�r�9�n<Q����+�r����q���g�"�Mʘ�q���W�Ap��uW�)x�Q��`�&t��i�C��P�&
 ��.2��.��l�C��n4v�����ɘю|��3XbF�/��*��=��j)�Q_�\���K���I}����uxm$�}�5sƿҍzJ�7+b��W��<њ��]�k�$|���g!��aK	U�Oxy��N�wN��+f�j�4��&��nLX���ӼyCx����{��vw#�&��%���8E�C��~Yz<��+LY�m�Ə p{��P)Y�\"j�z�ka��,�$�7�T�Ɍ�q��J6,8���,�)Si��v���h�%�	r��Б �N�lHl��p�.EP)�}��P��`)��LI8k�%aM%jx�e�Z��1��͛��TRp+�f��L.D�≠�{�+�XB��`��[|ƻڛ�مq
��S�0�+$�1��~�&���=s���R��#����u�c# &�~C�XHJSg�r�����۵<�X#�
��n�����OT�Ŷ�p3��OiC���,��[�P�[�O� ����]w.��S]7�n����q)�99Gk\\\��ƿ����H9*�R?�Fk�(c=��$h}���v��6��1�K��?���d�eƨ�ȕa �+�&Q�M���Х��7�T�;��@����$[z}��U8L\�V*y�4vU ���"�l����P��}��w�ؖ�&.��I���F�L����Zk=�
=��̴���U��>1�W)�c�e9$\��	�p�����X~S	�x�J}٢&�w/�$3��P"�2��D?o�S�$�/b�'X�K?3�^�������.�9�x�`�/���"Z�*I}�+��N-��Je�簎��کm�w��΋&tnqT��+�Օ�́k�/�`�%nDN&8�>͍
�5;d�ų�B��sJkK/{�����F��ۨJ.L�Qé(��m#���2m����K1�\m�� �:��_(6�S>9 �`��4�W���R������[�6���K�?�;��naF������O�m�kC�a��po/<�	�����J>���urQL�-�-�4z���4�x��_ ���Yӿ�Fo���,e���z]s�;F�'i�+ޠ*2M��4q��lG_u{�~$6֥L���cfo�����*Ռ\Ht�,P�k�A�e�����n�P.r��R6L��s�����<��$���c��5$b}7䐃ʏV?��T&��9������u
d�G�c��%n�<(7�l�u��(�cb�O|+X9+']�v}R�e�:C-���kMs���F����֐�x���Q�&Kb��l	��{`菬��l$��h�{��^e)���l\��QB$��
f�͐� K@IŶ<JA=ک�J^r"�ץ:R`����O�Pk�L3qz=lk�(nبɂ�|r��K?�еt���e��m���HK6���b1��Px�G����c� �=G6��86�o/{\�d�R����B��Z�E���7�T�� =����$k�<s��)���[��|��F~�c�L�G�rب�p2n."���E�k��9��vL�Ʉ���n�X
�����,��M�o�N�5���n�0�1�BVp��z:g�	�����i�����#R8'�?:~ݨJ�]��$�±"
	[��O��0��^�č	�6
	�2��[� �D�F�}�e!�7�B��93���w���0,��-���d�uS���=,r�Ԁ�c�2�;��Øc��Z�z/X�������D�lRZ�I�>J�����-���H�8�j��p��)�Ɯj�}-He��I�~�H|�IC(��LB��aQ��i0��*,��D��+����| L1@E<��ݦ��R�9Z[�U[�Jvz�S��'J+h��ײ�ؙ�B)�������07�7�p�=ǎ�9��y��	�7i��<���g7��٩�C"a��$�j��J������*��ϖO "H_�^w �a+$�\!4j���v35&�ac����ze�g�-�T�mJ`۔�V(U���|�Y��S�p����8�L:#���F������+|CH�YX����l����|������J����OS�'wN��yK	?��Tfn��r�!���˒!*S�铔���� ����ҩC�!_�{�u��N�d���+ok/�/��֬o�נ�1�U���.�����<�=�H��+���C��pEzki&EQ��@�A8����n�ŝh��2Д�s
Mo�H�p�Grx��oZ�ۨ�)цZ���UEe4{5��\E���r��� j@ݼ�m�vUI�Z�5^i&\R�T������E�V�Z��t�$��a����%��j�h���}�΃����Sk��\�nm���bW��)�^p��_�V�s�u�Wȝ�/��Ĵ���[+E��WA<5���&˖+�֊�D��9$�R��;��}s�In[j�i��1Gh<+V���K*x��{���y��i����G��ڙ	�Q�D�5дr9�� H����M��n\Z��K�gƭ�ap��+��0d���n�K�-/b8���67�#������师;�=�1�7�S��DTr����0�b]"�[+R_�pO�o�P>}*�{����9�������+.�plE�J� Ua<�&�u�È��&���]c]�@�g�4�(d-��A�p�֍u�9/�v|��'�(�����/�6��Al��^�μ�3��������]��K
v;�~�ƃ��w	G��L��� �6I�j�^6W�K<�)`�|���N�� }�B*��v"��+���_����6�0&tF{/�;w�?��\�Y�j��SXj?�j Ԃ�.a��uM����P�a��*��!�'�c�lH���涫�/إ��+x�a�3��~���m��K+7t�>fԮڒ��4�F���ߝ,U�%��]��0%%�n��wy�,����b��783IC�Y	宣�&�N�V�[���K!v��M��?��&K�x]?79ۖ_%!�oN�b�"fVڴ6t�~�ZQ��X;��E�4�Mb�-w��[����|���}2Ӄ���[:?v����J�0#N�I4XK��2�]c�1����`��;h�ںTM��m���y���3�GH�;Z�R�M���6%�*@L"�}\�tj~���/�u�e����!�?ɻ�?xx�Ψj3څ�np�~�E��*�o���&����*نū�(�	�P�"���= N��᫇I%>ឣ*������0�>]��]\�|,?��)�2ڀ��v�+�
�������Қ9�$u&K�o,4%z���t&�#�|���%�&U�9A#6�8���i�p�F�vl�� ����r:���clM�$�8�<
E��L�LJ�Y���F��O3� ��ᜟ]�v�e!��{�5pߧ��RgU
�3�-�Pȗ9����f��kׯ50���F�5�h*ʋ�q\��NAY���?DZ���k*9�|������l�
;��<�o���N�	L���LkKW��ȏY���(��e��c8�����{����icv�!3|ثgL�����6�K!��Dq�O?c��� �\w@S�N��
�d��-�Z�M '�]�9䎥vU��)�ȷ�G�r"(���Շ�|�춬8kZoE<��6�2GF#�Q\j�y���@�TdnZ��
��AB-|���2�����BSl���(��!��{�ZV,OI�P�	�VA�����7�؟c0O+zꀼ6�MM ��1mD_���,{ZD��1i\���V��q������NFv��@���ݵ>�sl�Os�JW��mv�b�0gRծZ��w�N@ڪK8*�8M�v���z�?m/GWǿN���+Y��<�w�T���9�òq�goA���y�8Y�8�	����q/�{�����c�Β�44mN��HY%����;D44o��v�3jFa��	g���+���_$��&�2 �!�
�E�Ы��LP�0���+
������w�p�^�]�%�����X�W~X�ϛO�.�Jb�h�
Aٔ�,a��Y����v�5��"�����P��ٶ.�n�3�ÚAA@D��SI[���c �����f'5'�+e���ۉ�4z�"|�A�~
:������d~��(�V�x��F"������D�^��T#��P��,m�q.�s�o�f �H.�:�-g���]����t�R� ����%UssɌ�����"6�6�����|��!�>Қ��i󽗬u�a��}?[�K�L8�z���-��<3�R�~��P�Ƴ.���J��8�ZF0I��J-�Y��TY�e(��3B
Ӱ�PA�Մ�l���b
,jY�V���_9̹0�G��sW1pr�CL>���ũ'N�<-��~��a��M;e��-v�_���g��ю8�� �b#So-�M���1+Y���$D���7��|���s��;?':9�p;�ە�\qKIh��ӫ.8�s�Uֵ��F�/�1u;�X疹���:�͆�C�nu��A�����j��ظ>İ�uABl gM�I�c��"#3����iۍ��r�𗗎㪃HY|��*A�R�� 0� O*��\?�~���e�;��Գm���F��nq[��p�_�^�PL�U�&�g��5�ɋ���x3\Zi��?l�!˟� ��?�*1~4��o�������8����C"z��UU4��?��I����Ç^fy�))*��3����+ �s�U�߹.���0��t�{?�Q��f�1M�G���~ԟ$�H[+�%C�~Z�mZ�>Ⱥ�P{ǟ�A���e8�h�NZ��kR�+�[8S:]Oԝ]>��^V��4W#n_���&n]S���+�Yx�	���T�A[1�+�j��-���[�x��8�L���ے!ܯLZ���쉩�zȈdU����@69M����:�����RMq�Fm!t��j�8�\��2�Z;�P��:(�!�O�.���usd1o����f�&2��r�P����V.gy��P3��~�l����T��U��膧� �tmL�P��NΈY?��u�'�
g#+��v�dQږ� ��\酏�\%~����Aj_�i��r���ױ��--P�,�/��sH�Y�Ҷ#��cR-��g�h�h�o�J����)ڠ��a�PÒ��cP����]{��J�^��;9O}t(:�t+A玲*�\���2����>qj�TD,�������:0۫1�gB�>2��������"Gv}Օy-�*�aH~DZ�57����W��D�KP�$��[	976vw,w�Lm�/�k����-=���ҁ�WdyK=g�
�e��h	�@�Zhڽ��,*�(�����ʼ�!�u�
�(����@4
v��W��-m�i*ffC��%9G������!2�Ԙ����f�1%DFEW R���\Ma��u9��:�@H���|��5w��k�(v���M�[�����_�L�;2���b�z�21����U���%��O0��Rsb����֤�Dq��3ÀdZz���r�ҘU܏��5���l� :l��a���z�
PO;�=�}F�2��|�R<� Z�_��Xu����b7q0qtx�Xx����~�i:Mnߞ���Wb��j��������a��j�tE��k��,M�)s��M���Wa���:S#�4D��1�
0�c�`�A��ډ�ֻ!`�B6�[��01���/lK��#�ӟ�x���+�"[�Z���$/��~C��/�ˢ�����X.��a�]��5�LhU����� �U+�`��Y��A�X����Z�);넩�x����oF,��OF�i|�]��j%�x(O���#��)~ԩ4�&�L(p7��q�H�^n��ϵ�?��O5�QkHƚ|��0u �t\�h�2I�F3O��m�v\��կsZ�m��E��	��Ѧ
>΁<A!}{6�F����\��x80 ���Dl���?�Y��J�y�J� �2�}UH��]�;�1�����\BŞA���U��TPs�.����<� ����!�]!�K���N�U���r_���h�B���#SI�J^�~��*����b�-�,n����n/�K�Z��[9��`���2��Y&�;b�;�/�D`����-�D����ý�eV�TЉ���"r;+qC6bD 豗��������y	H)h�F���g25E�D_oq��t�̢�����5�E�Z��ƒ2	�
)�G�	Բ0��C'J8��HǢ�IQ1j������ϒ�E�(�I?!or�6?2��֫��R�pN��v�ۨ�	����Z�6�\�7�/2C1	�M����T�����PU�o��g��x9�	TN����ߚ�j�ȉ�y	�Ce9��
ܹ��{u):�l�)i�Ӛ! alI�ew��g?����̖ғH���mv��
M��n̖��vW�^�[iy>U)
�`�'��	�=h�@��xE��Sh|uj�B�����Cw��Pj��I��69�O����nk�W��|C�����"����(��ʣ�J��кu���n��?\�h`2i�{
*C����*?m�͋l�^������tV��\#���H�2s�ZV x�U�*��.ˏ�4�����gx�c�Lw���%��xT
P�Y�)��Z�9������@q���7.��tѰL���t:(���D��7��3��B�Ԭk�_[�V���h9nǥ�w�u{�>�=Zx����n���\��ώ:�hvU���<��+4�u��|u�\��G/ �f����?�a�+��= �/���R�0�0��m(>ӑE��+���P>�j�JI3UF���H��R0�H�[;�!���`���V��(��ZL�%M�_�{�ڢR� �q\ ������8��_��3>R]OζA.�������@�}�lۂ�������d�4&���sJOi�c�: ���{r�uk��������y���n�Sw�ȗ�O�Y�Eo�  ��z��.��5�> ����{W�敾u%�|Y��G%�_k�M�Xڠr��Խ��?|��q`B�f�V����p��97�>��4�L?5�r��W�a(\F���秢�;���;^\rX�~�&;	q��K7�'7�9�,����0�5':|�}･v��^�[ ����YQ�������R�Je�ލ�A��'���kO��r��цs��|^VoA]l�?�w���g���RqZ��-�gϡ�`\66"55�>f���|�Q~+&rO~���DX�r\=~k�E?���~^|w��f$j0��e�*{)�M��o��5��$�
��&7�����k���\�6�-�e(�����[�t�;���f��/1z�_��z�o�����BR*b�0�^O(]a��mZy4MZ�i���K�	#������\�~�{��xJr��R
߰4 �8^���)�9�R9���Y˿Q(�zh�͒Hl^�=[�����4�K������{	�qO����I�*.N���{� `�Á�Q��N�f[��oS�<�4����̈��V�G�	��?_z�a��iu9��d��PHo X�fy�GW�cp���N�2U�84���kW��@�j�q��|����֤'��k�J��r�c��ۻ���@09����HkV|��܎`��+�"�-� ^LŷrY9J�l�kXރǶ~��g	�7
H&�k�h(7�*8.Ӻڨ�Y!d�;%��"*Q�c�ʗ�u�?$��V9�E+q��C��4��7,ͪ�C�X	���B�g?���T_�?�;�H�K�;!n���*v��и�rwh2�A~:�;�cm�2<Z�s�rNJ�dj5۩=I`�6#�71�ַe��x�I�_�iD���HC:J�.E�f���3[R� 9	bR򱅺��~Ek���0n׌\ <}is�����{���o4k�
��2����uu�!$j�M�_����>���Ђ{�����v�%�����0S���EFtc�ҫ�i9rD���<�:ͽ׹����o��C�M|��9ǲlYڏ7�&!x�Vp41�h����a-ُ�˻�׾�b�@t��U�Y��y�U	ʞ���{��~�rQ�
Pu����e7������\!si�;�'P6�MƑ��X��1\��:o'�6���t��c��%ؑIӆ��\�Vg��2I�X/�C	�^�3�(�����6_��/�(:A�M��N��.uZ2!;p�h5�XC1s�WPN��;�{����\d)W�h�U��7�Z�~����>�S��F)�a*Xv�j��L��f�:(�b����)(p�7�z����o^F��.�^)�:A�(�5�S�;M��O2�ͷ������}vu_�w���e1$�o�p�#&~	�����w?��KWOP�<Ηݍۍ���U��3ʝ	Hr�M~�[6��@���E_�ɺ���8>Bq��T��N�.tv����6���۫�� �A[R�dK�D��/�7(�k��D�j������*:�8�*6^���b$�|m�K�]�öa��+�u0�@��D�xBM�H~���g�$d+�)G7X��!���ݓ�.�:��r'��=�dwZ��4SQsZ�:u(��S �-;$��j:B�CaC���NO޼��C8]�]ɜ܍�}���{	���?
�8v�		ې�xD�hSd�t�|����{d�u[,K�^=�H�Tq����`�av��ɹ/>��k�>����uDt����t�s�� ��yp^Z~�RK0d�@ �[1,梙�%�d�B�]vc��J�$WN����5g" d����0�ݿc��leUpi��UY^�U�H��ea���煰�j��Y��[���ɭ�� �|ģ�[�LQn�+�+�hU����wzg_�Q�VR�1�5��|l��ӊ�\�X��J�o*ᆨ@?�1a��u��F��RN���x[R�Uo*��Yb�F�~}2�\삌�C�ѡz�s��LM��r/��iL�3K��Cs��x�:.���b��P�'z��fq�,���KF��T��ɵ�/��=`��{F���e4w�\RO�~�6۫O�cB:bn�1;�[�7,S'��61����SQ튧�0�'�q~�a>�$��o�QWق�����U�Ԟ��D��#��2<��#*�����%�?�� =�O�Y;wq���N
�1}��1��M}�N����~{�mS�ת������^����(�Ԣ7�=y��$)��o�x�� } +��<�����n{��/��/"@�{�ޯ6���
�0%�M�2��x�eX�t��	�� �ƴ�.���UԵ�&��Y��AoJL[��s��Y	�
E�la���sA=e��{ha,�V�\����h���iz9���S7,5�����00���C�D���vj��X�<�D��N��\�eq@u�D7�L��86/�rF��U�{0l��*?+���u�_��m�!�hW�=��C<3������+���.ǀꦑ#ؘڦxm�b�w�;�I	�߫��j�l����c�����|�:�C�Z���K�8���Ky�l�Vh�����s�/����J�O�&��b�R�)�u*z�*s$�to�6���fv�?!��&�$��҇6�7h�^٨������ʆ�X\��kU��n�p����֓*ɶo�jHA�n�Op�k1"�ٴ�M��)�%}�m�Ç��	�����D���ŉ2Fx�4��v����k*��ud3B<��d�"q��b��Y)��-Or�ne"@ԁ M-�:��K����L�n�يI#L,�X�H�m�s�U+/��m�]`�+��Vu�d+[��Y`x�j�4WV�^JQ冽�9J�1�t���B���w�J�Y�p�A���k���Gc{E,ߚH�G��H�*lB��CջI�u�rs�I%{&���Z��Gm��k���+[���`��z���%�#&2�v]u0�Y�Eu�>�e(�L��F��f�]N;���-�G>Ը�EN~x(��w�hL�dKw�^� ���X)�N��=��2����MOr�N��AR?��6ɃAE��[p����'�.��|3��LC[�f^�� �I��!�܁[e������LȮ�{���e��s����Au�b�A(z�d\����UH���ï����0��������e�K��!��=������L,�ל2����6�`�����Ք�nР�kfG���rC��Hf2�So��c�#X�v�\�G��1�foA�MZzSe�֑6# {4�R���Y����9��E�����d^�\g��n��a�Y���"���R嗤>;\�+Ϗ�#l�����)�j�闹�e	��#�8C0�J�^��u%�[2�9�R
N��(�u��g��`쏳}�p;�0�#_��.��cZ�_&L$���+��7S�֛ϝ�A)>��O���"��@�C|�:n�B]Z�~qѰ�j��P�1�_K�^W;��3Ai�� ����a�޻�����{P�3��BA}�\J=m��@X����$�|ǀ��ԕ�p�,�=�p�l5����0D���k�x��S�7�M۸��5����������9*We-杦��=YX	�J���_�����B��pwo��"������w����u��g��]j���H��ؑaIje>���8���V07{������s�-��ʑ���R���KH]i�<��Y	����g����$:��6�ma�&":����$��Iv]�!d������|�^Z_/#/��J�':p�:�`tvq���<��PB��lxg��./������3k�v;#�r=�ҸMj�l��<�`�tSY�w��z�.#�V��g|��ټx{$�I`s'lr�J��R ;N++[��Akڴ5J9�#��k�Ѱ*i-��'ST�?�{ɹ�o���=$2n���Q��}��w�#jH�w&����A7���R���;(�l�`J֥��#)��3�D�����Z�`��_�2�H.�4s+Q:א��49��O�R��VU�Q�8bmo�0�����s���q7�sn�!Z�Љ��8⎷)�k���,��"��޲g���ÿ�`��}�2��J��>�}�,,��/h��"��/V1��j{������O�Ն��-�8!ߎ23����	�\����ՃF�iY�Q�a�g�9�55���S?�c^S���ac9�&����σ��'g���{� @ˀ���a���*��;���ϧc7'���i�ՠhE��k���8�Z1�jI��ͿB00*y.�k����(-q���ӈ2���E��~4�}��t��)�y<#�K��R��f��%t����U7Ȟ������B:��%>�n�2�7GpgN7�"�Sű�e�oն��u$�2RY�aodO���̧Tނ���4�}ϭ(E���V�9,}j'�v)��3b>�D��s���Z/�Gի��Z\f�����G�u=� �oE�:�p����fӋ��@�����Z�i�w����\K�c윥�3�N,�6^?5�A��:���u_�pL氠a>xCh��ܥ 	l>��G�>z)�ۆ�{@A<��-��uꩧ֍�4��3��g9����=恀���|�D*���������Y�:]`��&�(�Ѕ8��-=�?���8����9��<=2ɩG��\���u|A�tf���tp���(=��T��5#ϓ�upr�( `.+�O�*+b��=�&|xs���Kɔb;9��T������q���6a�5Ϋj7��g)�m!��3��~F��x���N����&?�/����XJ��zu�zF��������Z'=}�[~�~md5�/7�knKZ�r���/P����0��ye�NW[�\+&�yLh�~�c�(�m���2���H���O��k�1r�+"v���֬`S�̱���gdM;=b�m�E���W6Y��fЃ�L�/~�&�0Uk�q��n<��T$DӶ[��*����`'xf��}��e�E*��,!g��`8��nĢ�e%���35�x�ALa{�� ����Bd�G��G|0�x�v�6��x�Q����@)S
,�~_Is���#0�%lАZ1ݢ�q��~W�$����σ��5#�h�`N�0�tx�r�f���� �^�f*����ćT}%�r�L���x�7��\�+�:t��\`Qb`�Ut!/g��؝��t�/�-~����/�x�p�M�X���5(��;Q��Xu� ���{u�Q�tsM��%��gS�&^zx]A�C7Ǩ��M����]�u�O(��sY|���e|�{OVM���P����j�󟁳����H��P��!�+�-V7�nN!�U�-"K��M&���r�8y:��P(�*��P�����x5�_��˗���^�XƧ�*�F�~SS�xS,�26�l���"FaP�̟����.P%���޶(�xj\�Ɵ-��*��^�8/�����p����(�u��I�y��,���Pu���9w!p�l$Y�@E�e5��^�/��xDH�	�_��l����i�,��;
�]48����{�{�B�m%A%���@��
^��cȠp[���:czѤ$� ��6m|`�{΂q�{)�����JD!��%��,� ���&�����Pk�Snl`���}=
�<	����_0D�	��H�h�;����ɴw\��Z.�<GFNZ��w�#B�(:smz{�o�WUڼ+���CR��Z�����y�o�2
�޸��~���x�5s�S�ECf�o���/�x���m��������k�w�J�8��2e���P���*����JD�f�{"B����T�b+�=w�G�+.�qon�u��qo�0M� jqŴ�p	���@^Yx�&EVFEw��cL�R0E0W?�W; Ccާ�<���Pӏ�L�tIh�(bNB��n���g.{���a摳���,�2�I��Ժ%�
��뛀�_��B�h8��?�<�囶����r[ß��\F������߼�������կ4���I _�#��C��g0"bB�b�]��V����j����YF�BS�.�[����}���W�����yM`#��C?��|�h	��Ew�DVF)�Ÿ@(ZuL�x�����wS/��Dt�C�]���%2@�h@�4��dv�d�vnbd�<j�A����t�}]4����;`�ڠ�n���u���=ja�$R`K���$0L���.�B;���0
`�Ki�����מ��q� ��H�&�ߔ� 7n>�42�.�P���RC�M;c};�/�k�y�U����s�?��\����T�:'��nڄ����0W3�f�D|������7�O�s�#�W�T�a�K���vw](�~��
+�����|�ty�Q�47��ȟ09��dºu��7+_��06��E��������HN�1ne~pL�;�
�٪��A���݉:����}q6�V]hK��YB�f��������&�!��g9f��h=c,�9{��$c^&�x�,�']Z~C5�mL����{&9��:���#�E�ϱ��cgK�qB��T��3ڲb^�?���A�ֳGb5@0�@�Y�Nq�#�MXϽ�-Þ~
�����1�cl�ޟ3|�fY��놊-��z�	��4��0]����ȗQ-�/ڠ2����s����?5H�R����zc8������g��jT��!�"�l��{,�z_&�π���ߴKݐ8�L�B����Ͷ��U��J��K6i\Z����p�<�g-���i��1�Q:?!Z�'2���!��O��q؜s��xs̛SJ ��e��{y�?�kP?��, p��1�enL�������p�<�9��{1��Z
z,���F�F��W�o�.�x2�����e�l���6O�����evD�Ɯ�Ǳ�s���p����Fi�q�&�]v�,�ٶ�Lx���(�:FA1�ӓ򞋯�$Ǟ ;"��!��e��pЉ�;���@⑫�I��A]��qƇſ��������3�x��.��������J5y���?�E��F<����Z1E�xy{�5I6�W�4Ӗ��O��!8̃�j���!�];�S>�%L�>�ΐ�:ɐ|��N��S`���@��4*�%Y�������h!#Ҕ���f5Zԡ ��Hd�B�5�ײ\��NŲ��y��xkᅽ��2�$��'.4���h(�8ޫ�](�o���p ip]�,8eJ#���(�S�3m�P������o�NGԍ��_w4RK���֨G#��C��9mF�@� �q{��l���	k�%B9�lJ95����}$���S{�q؊��`�l��d��[�� [q� ��Y5/�濷gX�qۚ���$�iK���d%�;?�?F�J��H�2�Mԟ�
䡹L�Z+��︤��w��'h��Mʚ��QVu<��)*!���%���;O��,���>�+�K����^��� ����g���xٺ��|�s�#{��Zz�¤KT�=��3OVT�s�r�Mi«`D��M��?8{�yV
��� ����IA��L��S�=3��ӈ,@ܑl@7G�H4�٦l��H![�H�? �UY�x��3E���>,�dF��c簣ϑV�W��Y��NM�������I��w�nҬ������A?��r�;8:�|�'t=�~��$�q��s��J����� b��w�yt��+��� ���RH��#�A�vm��hG'4�ӉX78J��X3_���Wh��^mR�6~o�o���)�f+э:�����(�{��Iʃ��Tc(־BpxЋ��f��Bp�{�� I��R[�0����������WPt�53ݻ�����'�5��y�[��W�0�^���E?�<�0X��9>̦b/��l�]�h������<X��Tw��צO��ۉ���I�V��h7ܻI3��L��N�� �w{�|
Ue�e�T�A$R����%!d��s:�@+$�;�����X�Lb0��`��o>� ��'�6��tF�H:%y~Q�軀pPZ��&+�������R>t��Ja�	)s�����Y���H�l�-�(e��"cZ�{LW������I&���`��p�P��<���|<��NϚ�K[k����Q�5�y�es��t�!���f��>��H��۰�t��Q��$ʓ?�ê�Kh�:(n6Ԛ��|�̅�dG��Ưh�cu𜌙1��ef��P��R��a��X��2�|/5`�YG<�V�=��`���e+~@��Np�������WO�D���@�t,�<�n�bL�S.�#�O/��=��sd?��%�ll��v�9����ٙ��G�4�ـ�a��Օp����2y��#�s��3�A?7ME��ᢎ�bX,�2��<�ܳmF�e3����x'��F}�4f�˒*�*+v]�̚d/����wh�i�����mꞻ�}0�/�A�h^�{��@���n�ݼ<����� bD����s�� 7ǒ�K �IHAو�t�1��Te�����a�*��2=γ41cG��f�1�� �9�:}2=���#,�y�9 O�&�k|;2>�a�ѐ�� �F)�s�)�ϳ�+a�&���iD��	4+�
�L�.�Q��nɒ.�qs�؜���E�Ln\M'M�w���|���t�����C6���$��hT�Zcu�^��F9��~�C��?`�ο�i�h��ľ[��W!���>~��o'�E$�An�ZA�G77�PL ߃6��໾�fu��
Q�e���:�!К{K����G�\�Ч�q�A��WQ~�\�i	���s24]�9�M��Ƌ��~�m �9���F:�C��O4����G������3������P���z?�F��InH�Ɵ
�n>1��F)^��x�� �>��6�|~!U�F���i}��^#�����6��*�NXPD�9anl��d�Y�V0��i7wł��������D�����^F*�X&v~V���4�l�p]?]����q/�O>NX��:�X�J���#��g�n������Q5�<��B�@0�M���e�d�j4)o]����0��[Z-UC�����iʇ:�x`���԰*�_l���4Z0ΩI#�-P�N�EDM��^u�zj��bI�����@��"�peڈo��g� W�����3�	x�+~u�Y[K���L�u˱�9;V}[�/�F����ܠ�fK&N��К�D͉�tQ�N���zhϞ�J���N��pkW��6yL}�uq�������m
`W6�y�*x�T���V�p>4�m����V��a	�k�7.|Z��p(����nf=�����
<�coi��\ض��ޣ�=����<:��3.,{�(��/h�r�mʤ��x��#zs����c2����D@h���h������D8<{���vKwQV�.�����b�.�b�9@���[����8���6��`�I�Zl����!���w"(��i�`]�Q�%0�GI�	�������X\X�p�+���:wJ"�b���Gm���-\�����'��Ëk"���kD��:!����v,l�M�<��iJ��،F�$<����*;:�d����9�G!Le��ƠYܧ�rEO���N�߮>U%��<m��a�Tu��6�c���C��3��+���3lV���L�7 �{�����-Q#�6L��!K��^EY�Yn�F��~�d�.� ��Up����Ǚ����!t�h��ՊN`��Z�ƹG�W����7��2~�m��w:g�3��	~ɟ !u���%+φ�h�9cx��m��������nIfk��(uܙ�z@������]���k��"�D%�,�F��?Ŕ��*�ނ�Ô~|z��9c����k^%�56g�@ Ko���p3^P5�X$.�̀ar��F�@�p!�~��i[��5�0r���|�c�U�1�!Q۔�2��#��(����%�;
�}�`=�>��
G�Z�]���Vs�TB�6V��o�����_�	���)k�olSg;GV�t�?6���TV }��=9�e{e�M8�*�Uq5�|��N. ������D^VS6����+��x`Bqu�X.�"�p3فU�?�!��Z����J=/�_���|X���pak֣"l����Bv�Bw�����wU�|Ƹ�����>*#g��fFn.2�oá�N��#
����X���n�v�^b=�~��8�\��2�j�� ~P���FfL8)��[�>�b��%���ʮ�E�=<��d4N�G���0�lQrZ��)i[(m�m9��߉X�
�d����t�W�0��D���+�ۏ;��NU&dw�i�6�x�&����@���u��͘�L��-o��]Mb�i�&x�3���'��rO���97F֬����+f3[�Ip����fo������*��?4t�~q�������T��%N6���O�MY�9	BRV~h��:�*�5>�y�X�͇
��A��\j����sv_�'#!�c$�K0��?M��X�5��b�UŘj�	��]԰�0tγ��d5����D0ROB�$�n�<��M,u�#J^8�P�߿�{8�.��WQ�?�t�9(�'p�P��Q&�߹?������8th3���e}J��jY�b�����w�"�Oy�Kp�h�/���`L�D����v
4��'q	� � �l��#+���C��9����ɞ����pe����������d4B���A�D�(�M&���=�����l��Y]h�`�$*�2׷R:����J��?gQ�h!� ��+͝i�e�u��`3p &f����%�_j]��yz!�&��it�n&Bz�8|�H���^,�e���ۭ�=��2��S�gB�ol�6!�G�3���b�+�qf�h��Gx<�<3\iYbN����[]Y�mo�w3�FP������,H����J�Y��
	��2w;��f��0�	(��"/m�5 F��W�*5��0s��ܿ+��h�(�+�6��
�@���Ju�:m-�ڝh`��"O�k1$Q-���!���<�/�C���blr���B\����j��dg^�6W9F9��}D7K����/w�op������*#�ʮ4�`����k*���*��C/!�p��=B�����2[Ǫiȕ]˰x�����S�ڲt�|ɔ|�ZH8�书�>����BQϬ�k�F�	k'��5%C>&z���ſ��+�^�-V��Rchd~�"5//!��ْK����
��U��2MGf�o�1QG�` p���}���xӕ:$��`�nx�2��Wy0lE���+��WBH�q�g��1'�>,{ZՏ�!�[M�O(��G��� =�U���1`blʴ_�v;�t~�.Gv-�Z�0�M��`pw�ɮk~���S���
qN�01��C�;h���I�P�PrQt�iuN32(��XX�۰�m#�#�T:j8�����Ħ[�����S�h����BH�'^�)"�|�g�e���o��/��4��V����a ��2u��vi�f��K��SZ����t���.4 ֕uS=�ZTЉ !M_���e]�a��Q�^�X
�DS��|�؄T����p�կ�GiW848eRE�-a���+�b�c5��K(悂A�c��}�
��l:Ei��]�G<�!|+���S�NIR��j�F\���66,/���`�d��˼������F}
�W�ם��װ>ƜOٵW�'���u;� ����ʦ��.����^q?O{�;D>�\��Z5ڼ�+��_Dv�$���}Ne}(y�}TyIT����KO`��q�0���ջWOp�ߔ�!�$�b"����k�������<%���G]^��C�@f6 ���1���V�F
g��C�Wk!q[�ب���7м�z]&���� @ŹT_���� Zi�T�Q`�\L�%O�^��	�и_z|o�^�4O�k��jfz�Cu�{��1�(�\�]����z���#���M�TĤ�8�AY��n�3�X���T�9�V�)�@��u�̧�r��M��V���Ţ|5�q:XD��[]�|yQw=�Vٟ����on8/�C��2o�꫓�-/�� '�Ԭs[Q�S\�����h|�k���R�}�ӡxX�+��9h���>P������iH�~��0��C'~'�����G@(��u�IU�i+h�BdETv%%��?�3
 >�ʴ
��N�ĦQw�>箃4D�<`���W��;�WX�r�h\��`^xG�j��<L�{�����S��nR�Q?d9�ג׆x�嗢�\��0�9c��^Uiv'��L<us�R`�y��q���J������h���_hTG6�~q�}�0.<�`m�@�F�Q���r������5%7{�WIr	Z�(�t&�O��$���޷n�_�R�V�Cȅ(u��[K�u����o�	 �ػ��%����n��
9r|m��!-�֯-)�G�ϕ�`Yd�f��e���]���e*Ty�͎��A�WA�=��&#�ª/*�����*���?�i	��K[</�K�daͨ��i�ݻ�\D"��*h�:��=�l��^�Uz��R�Q���(�
Jކ�de �}����s��Ʈ�55��oZ�Y3��]����R�_['V���Y��4U������(���w����_���މNh8�$��V>���9���:'�����/ �	Z�AZ7fA���X�Se���]6Ç�JM��4�5	�p2������6|T����R��P?$PM���2���XO����_`�z�`	X�;
����ۿa�YHU���N��{� gLd����͕H7�#Qd��j*�ʜ�Zn|I๢�zd�ܧ�g���}T=9������q�C8��������h����5��jq-��*�(~Ӂ����^�� ˑ"P�C[w�˸X�q;_�\��
�,~l0��)c6h��r��L2�U%kp��ϧd���
9f7���<����t��'�N6�w~�E�5YY�Y�͐
�+��Qt`*v�}2{��5lYz��Dy+�ff��|�y�Kj?H�[��
��:2; ���?�&��L�R�6�ҔR�8�U�[���ّܦj^P��w^�$�jI5z��[h���	{�dp'M:{Ϩ��z ŕRM�Lc�5w�=��F5Y��jg�Cp�x[�q�O�)���.W� x��8ȠV@4�<�uYJ�H+@qr��u=�� LN.�x������Ns�6���͸�i�dO1l�:�`Sb�-���˳���Sl�*�F�,�B�#&�)JE�f��huv��N�%e^yO��_��u�螷<~+l	F�L�����}fTX^�s������9����ɤ�U��Arc֮��p���Ӆ5�$�(�ZO��~�Tm?Q���_�?Ke!�-!X�^e)�7{8�v�=bf��@�?����6$P���'2=�!��L��W���q�/Zŏ����Q5{+,)Evc"*S��e��K���8g/An���=���lz�TR�sp��*]��FV���=�*Q���4i���A�$ph��Da�� ���:��D`/1Ӧ&֋))8a6+x�Y!(�YH�������|�H���`h1I0b��~u���y�o���{C��^�5p�Vx�W�L�:�zF��)Y3W=23��`�����[�Z$�ψ7b�f��.&�ٛBm?_yN@TRŮ�4$����ώ��>����OO��)�c���y�I?<R��j7~ċ,�t�tB��샇>��!A�F��xڲ��j����Z�Q6���y��� G(��wU2��:-�SSD��.��Ք���_�e��*��df��O�qd���7��d���u�t6ڔ�d�f���ll0����{�sZ]@s�W��Y��B��n�|C4�E��#�EE�-�[�s�5��	�a}��� �蟦�(�H��?f	�}�9K�{�W��^�S�Ʉ:'&�����F��y���*��\�-xG��l��)�ĩ��X�lJ�h���V�����7���Iꋧ��+'��0��nj읕�>���f0�m�{���*�T����5�ϙ_�dəྲRqq���Ä*�f:��q�������n;t�&����I���$�U�S����·��{�HE����|�O���Os5+��]P�H���Ros��zۛ1�5�:��ps�����F�q�/"O��7�z�1�� �N����B�iL��NV/K�$�"��'&$4�V�� x��@~P�f��YG�U����o�{�KQϋw�7��z����}ae�� ��1x�3���6�H�kU�jw���VǠ�&��tFt����5�֢.>b��R,��g*0����]�Ar�������N* 񾍒����m��L�b�6�d⇸hIQ��V�-,iÚkNL�Ϳ�ꔖ���Qq�����"Ǎp:��W�r�N�M�1h���NA� ��c�д�R�z	2�Ձ^v��?�[���N���ĲA��ϯȥ�qV��B��d�yh����x�~̮k�&rtC��e ����;P�G R��(��a��F�������y_��H�/�.�G���=��C�0T���]o�@��L�57����&�^�*A6�i5-/Ŵ^O!xj�G��Ғv4���e�P�m��= � ���RxV���I���/�8>���_F'�B���Um�0���*����W�ξ��9.U��=��/8��6������T�(�4��v���`�r]X}s�m�������� �=�X��&�q^���8"w��N!�����&�Z�ץV�`�$]CyL<^������s���h�� [h<8�rS��^��i���W\m�"���ޔ�a���%{Y��D
�u��� !\@�~���(H��}Wz�9>g�E�-4ߝx|�-������P~ƴ�dJ����ԉ�Μ>
[o����x��@p��*�Q�W�ea�aZ�h���FN�����3,a6q� q*����?���Fӫ��a$"b$���&��0>���L��/w�0�6�J�h�x�������>S��;��	�!����ca�#��Hb�י��\0��D�(����M~Q4s�j
��`<���s��<���Y�c\F�S,�(�P���oz�/�ē�!����k9NW͊ ����g�D�կ����wz������҈�9���wx�=���g���
�� :��n����+N�)b�!�.�z��D0��'�d�?u"�,�,��=qZe��q%��\����S�I����i{�*G�l@c˗�YC�@l�D~�+�
5{�#\�y߰M��ܦ��"�G�����b�l���!��g���Wh�k�ep��K��mefފ	�O����]�b�sT�����#���9k������@OPm�ӂ,�h���Ӧ,g�|���
=�k���.a�h�@�������Ɉry��It��-Mr�r�e���V���ʛݶ*I��9SuE���h�Z�� ��z���SkG?5�\�|c3_���~���܄��:�������ű+�x�����[�)���{�#�Jp�á#q9I����n�#^K���S^6���K%%�hA5�I%�j�M3�K�B��|Ki��;a��"<A$?���J]ʝ��T�K�h���z��ǹ�I��A�ۇ��!W~��MO�����n Q��1��y���N�2|W�L�D�Zŵ\T�r�tp�r�x��+�@3��E�NJ�`���O&�RcZ�8ߛ3��
H����k3�!�IVΕ�������.�bm��!
��̜����Pb�莋:�ŨZ	�l�/�{TG�תc�ן	� 4(�'�}�E;Q�Y�$r\��qB5�g��P�^�o��+a�����KP��������?̌���o}᠅%M���{?E�߿W���SRf,��J8�!� �/,�m�}:�JcEGw]����Ż�B,���i��,<�6��3�������N�T8��&�s�j���&���y3郼uDݑV�=I����]h��[lm�1�|X�/:"�C'�<Zg;�J�E�Ƌ�u΍V��G��8wH��i���)4���&�8��)1�`i��0�9�Լ�҄	r�E#�d~*2�����7�|��oei��v=�Лr���a�u�<�G���bl.ۓ��C���O�Cj���Wy/����O�e=�j�*
��X���fW<��͚$;�V;�_ ���E�̬��ԓ�U�lx
b#� ��0eK���[N�������l��Ӈ嫮�L�Q��׌�w��T����4Y�B}$��1-�w�����bDi���$�JD&\�f_�R�؛��wɝ�<�����_��ľ7j ������a���h�"N�OsX�"x�3b���i҆�_&g)G�B�_��׶��e4��`������-	^�vz��"oʍw]m��/�� fld�h %2N��J�A�ouق"f���N��/SKD�������|��,�H?B�B<�d�=�z}��\Yɹp@3��w(�[�-LO=U��6�vSѤ�B_+R`�AOQ����ԛt�M��g���ZPz�Ճ2I2�Vc��#
���p�!W$���$�Z]���qʛP~g/=<�TPlf��G����c�%�3�*Wm>��+��>��U��Y�XiP����[e4}lgV9��$��<r�T�%7��W�2��I�Q��\k����%���e���cn���)�/r8E��`���y!2)�c�z�S!l.�������&�����Y���"���:g�˦�_���:�u�o:f��z�ɤ`ni��-K�_!,>����2�-|��?�B��*|PTkΝȺ�`O�P(+�2D����u�VX�|�0�Z;�[��nu�^N�w2q��yD*�b�ۈ�,E�3�n�䳞C ď�V���6��	��/�x*�3��I=ʬ0m/���(S�9��#oڡ���|jü�h� �})XuwN6�d�b��t���5���Ha���.G�LV��P����S$M���X�W�В!��֭וa��Z�t@2=�}�o\&�A��������T��!#�\��u ,�������<�7��Lؾ�D3�B���׍[筞�z��*s�`Ӏr���P}�����ӂm��2c���ݲ5���X)�S��.�sӲg厾�,�4���j0B~+��*H�u~�U���|���M���Em�r�`���8���g*���?�\WI�'d7�{��ٓ]�f��AR0�-�c�94����Ɩ��^T��f>�
��t`CI�Az��|�G㓢z������5cb]�=����$��Y+"����z�և�~o�9ʀu۷��c�apʰ�~�E�B��6,�݂me��VX2�gv��Pzm��7r�U�?�S<&�:禚E�Z���3-{2*�`R�SD5wʅ�ǊUG6d$�r
�p��D��`r�FJ@W��c7p7tz��u�'ƌ�� f���F|�k�%�Ɯ.<���O�_�B5�pbE�Ot��{�7o�H��13��&�i����T�D�)�'��J#W�t��<%��-�Mp�B~f��_~^.�B�h����׹,���# Q��u�|����ҩb�/ 5��	�W�1�����%�=�?�Yؓ�ٓx�sPJ���~#�,SM� �*��P֞E1������	��NP3V���
����>y8�x<MIpz��@��}�����P-��էo>�l�~	sv=K��7ӐÉ2�D���_:Le@�J�$%ܞA�k���I��j*�-r�w7:n0��f��d��]|�]����h´]q�d�yX�BG����Y\~�TԺ��n�3���=z��=��U>q U]%��yb����)�����N�Փ���s�W���{�]�$��~���Ig�l�ӽsc?|8�eO5*�"�.1��H/�
�s�Y��p�fA5�mN=�u\H��.��1.�Sc��v^���Ju�eN��m��=�٤<V���جt������Ґ��af�
�݆�F���M�]�;�ډL�1|M�g�7����C�x'}����z�~�7�D�%Tn��I1훒�*fR�/;�j��Q�/��Ň'' ��w�D6\3A�j]u��ZW�c�k���d�K-E��K7�5��
)_Z�W�M���#U��u�����@M�Iw7��I��N�6�'e!m(S��v�&ݿ��v.t����Y��K0���9d���{%
73t}`v!j.�%�h�Q1W5駠��Ha��8��'��`�ƫ+�U��4��i A1��|X��!PE����A�B|V��BK�C����w
|�X�Hi,f���y�f����MQ�*/ÿ��R�Y����v��d˲BJ���ؾ�V6���4�fܕ��f����:g�u|.�7�z��t��îv�bP��'� L������J�o+��L���*�O��%�|3uӠ�4Bk���絯�P���9��	��qt˱Asy	�ay��.�S�J�1@���q�B3\!��Kv�P��̖0��� g8��uM��76�I�]o'!���-��Ѿ>��͌�F�Q2?nJA,2��q\�V�9ȫ�-�\��K<��[��S�ɮ�1M)�۟��lFWy��'wP�by��/6{��՜1w��G;`�dh��e)��<k��Q�"ؠk�z>]�l�dj�Tg�2d��ԁ��q���.� �0��X�a�N�"s�ش֏��6�E���-��Z��1C�H-M���z��Ÿ�)�x�ۆ!��c��!���)*����a{�[�X��j�����$��G���^m�$�`��g��X�Ś�h���R��5c({�ѽ\+N5�3��dd���eA9p6Y�W�T5p0�giX�Ɋ0k�}�f�_hYU��%`S%^Q�a�{�Y�5 =�I���n7�<�9���3�Nhj8����-�e+F�P���%&�� �F���6�1�5W�
�[v�d��^}ͧ��&��V^�G�:�@F�h�#�Bu���@�R"�����q�q/��A�Z"-ڼ���hl�H�P��Q(�'��+u�f�R�<�y�1�"%��~k�'�����0H�y�-�Y�b)ߴ8��:�ʧ�~��&O*�9����`!U�`y���B-�k$��#���x�Ú���%rG��AT�(".��cXg{D޿���f�SX〙.+Qh{�(�@��a�I����,@�~¡�k�`�l/���)�>�<���]�e� t�\0���b9�BvbY�/ k@�)ʄ+)�+��O=1�*����{5Ws�\L�tL�wݳ"ȼ����p.6�p�x�h����>D��,��}��SS�:W:�m���S��״!���̙��d�R���V=��G�"��q@�0P���O�����G ��٠����=��t�-$����������R;�\�*Wq��.�
�bi�9�]Ґ9�ʧ�L{uA�<�[���t��5T���&cI�N�s��!�E�.�UP�q��
�-����8%zb����"^�p��f���7k4@
{�V�ϴ�-h�rɴו�q]em W�7}���M4���BY�H��t9~R��!Y�����{��w���w�U�m�ɫ,�);�}4\q9��!��WU�*��J���*��n�� ��]��S+�Fr�I�$��J0=U��!�1$BV�y�
^��ٞ��A �ج�A%e���[��K(	A΢UI� �S�rQ���x�+�&���iL��_Rm���J��������2K�v�P���S�nʾ)+�I?^ CZ-�G�ݨ
���M��S݇������Aq���8�T�ږ���l�����{�����i�'p���F�)������[���t��*�ϻ��Q���$��Yt��H��'�*\�>k�?!ǩ�"y�j=R5���g�04�u{V�\�Г1y��;r
�5�׫�J�w�����	���Rb���c~.��٢L�egt�ZC� W��bp��%�M��� N}��x�`Jd
�z1`O��3�X�Y�.	!���h�[��+�@.����WEbk�=�T����}�mL�w��w�n`d�#�X��QK��{Z�1���<m��+�@S%MPB�3�Kt���]�֤�[!G+u�є��Z�%☉����Q�Tk$��l@xw�)�.u2IG��sW{����!eUE�	�/U��W�:�#�p��Q�RV����L�a�I��8�ݚ�й��N5���mqcF�06%%�������0��ը���j�l]yfzVW�ø�Ξ��G[o;��u���o �s:K�ϚkI��.��K��{�# �����O�Pƛ{����lJ�v��2�9!�b�9���X�&i]m�bQ"۪���d�>��u@���S��JJ�%�S�U���]qc��ᑨX��w�yE����	��`��WC�� ݚ@��� K{j=7���gz�=���}!�5�1�f	��J[���:��?歂Q�Y�����B�pRL�C�,�uZ��|�&D����?�e�x�������jl/�Co7�)�q����i���Z��<`���E��߉c��6�y��$_�{��KdZ�WS��qCB�[�*�5�5XBFł˒˻{O?�PUiW@ ����	��0�(�0C��dAOl'�W��~t&!2�J/;��K�G��ݬ�0����;Q�"��RA(Ɓ� g�����,��۞qõٹذ�y���>�(�8B�]o��6s�J�L'���]�ل"]���B����!��w�`m�jp!����@�f�u�[3�ݕ����cA�Eȸ5��e�֒����NI���_�Ðh�j`L�^8Β��������mb"`��Ȓ���d%���r,R��>��zݺ
�<d�t"P 	�D�$G��!P�ϯ�@'K�P�2��4��>z�ԗ�/M�)���z�z~{�(ˑ���BmaVfY�*�N����ʇ]���M��o���
�!��'�I*t'�L�o�@��c��J{d��f�;s����%P�m�9�fM�L,��s@`���t5G���q)q'Q��t�u�#Fd���o��K�?Cr�m����X�
6�w��O-�աA����(h�Q��v�.���K�~�X"����~�$W��_q�W�=T�r�4�
 ϫ��+������ʘ��S�̿va'C��_Y$(^����z�^;�j]�;uf r'�k��9�������e���$��R�Z�>}�Z$����o{mt�ygc���2�\{e�6�.���@+�喓��:븂5ߴ�;�ڶ�l����<��@i/��F	};7:J�\���Q������*5�Ԙ��N�Xf���'z�%�c�A<�$0i�g��pN�i���;���]�����At����Pi�����P�]̻H����p�ˀa��ƠKq|�ʐ��8a6 HK���e�����Q�Lv�)Y�#����0	Tӷ�~��nΑF�b�S�J���(&����h4�T�cYk[,�Yj�r��,� �}�Ɍ��/�(��e|]�p�>M�♈�A�	� J�6t�od
q��|����`{��ݤK,[��˔
����^��t�����1� ��Ż#!4s2����n�w5��im
��k(�ƶ��$�]!^DŸ�_�	0�kK�n���9)^��i�&�����.a~V���������nnp]A])���MumW�	?���~��wK� �`27~-h{2q����������� I�� \���Co��5&GvȪN���p9�.V�3ś�gT�YV3��e}��	Яf��MJ��>�D{�i���L:�ޑ*>�Aa�+�݂��p�:��+�Se,ą����6]}D���JKH�*��dKtt\㐚�hoiDp/x FCÇ�I�~K���'�I{1Jʋ$��z��U�I��w��W"��!�<�C�&Ի�<	��cwH��4�К�����4��R2�ش�!�zu?�a�D��챤�Ǣ�	.S�k�Zd�]Pw
�D^ߓ'și�ђ'�����(�8FW-�&'��α2a�2z3Y�A�4��y5��y|�3Q)MXȕJ4�ɖ��9��3=ఱ⁂�֨�4�ߴ��]���[�7���F�^���ݗ� �?|��֋�l�:@����۔V��<:���0ƪ@�O��[=<�7!��Gμ��*������f����F0wk�KY���t�i+�V��9xsxp:��5��A ��?�w50��p���py>��s���x�\�r�L���j��(q�k�%Hf��S����iZ�S��>Lu��jP.~SZ��h�'a���*O �⠼��<r��|l9����K���M�� +��G�)�Yhg�7��E>�V���c�W�y���qnS��%����#���`��z�C�����5L(�e����~����{��jG�(����UA�c�`&:�ϸ*f��7F��7�ŝL�'I�!������!&�=�%_H2�.v�J�]�N��O��g���vc%��������B֪~���m14k�� $W0�H�yX �4e�������A���@����5�{�wX# [������dn��=;o���2���?�uw	8�����1v<�J��:''�܎��F\�F�$���:>�2ɦ��������q��%,�+�����t�ix�1^m��z@��?d����3�Tw �+H��8W2�с��ZX8�n0�lZ�b�������U.e�D�]Nn��S�jLu�H��&M�����`K��@a�	�zBŴYVٳ�IR7=_���ǅ�Z�Bz۳�,��z�[����e6@��_1	#.�?�qa��ҳ���0X��'o�-���0HO��:r"�9��4�߫�sf�	�T��n�D�O��`UH۽DB�u���\�	GID�v�����	- ����v<�\�#�U�]%s<����������S�N��>9��N��d���|��ᯠ�e��0/R��H�6l��l)�Ks�i�B���(o��F�y�X+����Fݮ�y��C� �mVrXm�3凴D.l����������i��ޔ���i�Ӕ�1i_��Ab�.m��(�$o��R��SH#l��.�d
n����JscXK�[j���A��E�P+E�!��)w���{j��K�}F08�R����2N7��Zu��p]��l��aUu�TCbw}I���T��ň�B��&D2d����!E7��qUN`����}��J6)����!�]��`�+v��	6�� Q�	��p��C�{0����r��$\5�c�<��IC˂�8�ʆ�q�VL<V^��d���zR���"���<?U��vٔdd�_�:E�@%ˢ|�a��@kA�$�U��,�=��e���kMq0��z�u��A0r����=e��;ً_:��̋>C� ]vI��~���ړ�N�w��4	�܋�Z-5��+���ꋦ��d��(���_�<�9�
Q�~��I�RҦ����U��Ҏ�+3Yz��bo��C+O���r�6�ń[�o��MQ?���Cm��A��c/G���L߾&�g7�:����N�{�(B/3�B����R�qI�����Pgw�u6���ۿS�B�U6�!W̷�>>�hP�BWƌ73���j��O���F�ؚ����2Wj�d���y7�or��
��Øި�n	��T���=�i���ģ�y#~4���Z�c>�h��R9�I7b��3�2�@��Ci:�Rz�[+o|�,{7��3�?	42��HlN�R�{�]8��(<��wMX�s������r$O��)�j��BQ(�B}&�e�r�	S�l|��	H{��'� �����8�-��X�8�K#`t�D.��E����6	],)}�^N��oB-�犩s���E�F��c�����4��4��@z�2��lVy���c�X��>��OKB����׋�G�l���f��ݢw,��$e��TfP-19ćp�0-SŞp+f`$����r�U��aqz��:���>~| �#]����T$R����~eP��Q�����z��15��'�ܰ����.�|'�K@��* �a) ;UU�1�f�[`4l+�ؾʒ��h��aW����AMj����Y�粆�� u�GPIr�ήE����h���. ƽ���3�!�`AY����X3NMGFtN�,&��&�۞a�$�\}^ @�����e*0ȃ�G(�g,�� 7��MZ-B�n�䃵7BC�P"�`"}���E��Le%-��`�Um�=�X*�[|�H���'WCE�̀O�$��#ʒ�Ji���-I���E>B��w����n��kU6Ҕ�m/�E6�A��"r7{�v�?1%}��Ze�k5�B��K^�3��R��y=�,b�[�3 Fe�j�1�o�����ȶ� T	S�>"�k�����K�θf؀hz0�C"��Hm�,n�,)d���0mR)�sO���0���t:9���D닖w��L�tڎ����/F'QqM�y-S�Y�D�L�aw�P�A�3L#�n�2�\����EI��Ԟ�6hf�p7{��I��0��l� �-gJs{����X �9X������������1���5��h�B"��QNVy~)j�^7Q���������HRR�'Ó�]�`C�eW�0y�q�X���bdv�M0p}��0����/�ŗbŗE˻�����s�\X;��'���^�e!3�Sa��`s�I[]�;)��W8�Z`Ue����5�@7����-x+)t�}�������7Ğ����U������C��?+�Q���-.55{C�q}�Z=��`�����8&m�N�Oz���̎5�P��������yTlL��<֙}3���RFE5}#
��`�`%h����!ϐ��3����(����}�`ӑ��U�"��x���x	q�ͩ�,�C�7S���{�%�| �G}nZ�#b"	+D�|/n5ɤ�8���!�����H��I \2���!���f�Q�fD4�)}:�Q�+��j+���qzh�ʼ�20@���Rv����� ��~��c����?ƹ8�(�$�J@#\��PEx�j�!!^9>U��e�9PX�&�(��o<L��Ao�K��Ԓsbnrc���n����*7���ڛ�TM����f��▗��?��|U}�@�Q����曡؋�֤�J3𧡎�X;���
�X�N�r�-�����n
���z�K���%0�Vr��B�[{�h�t}��|�3v��	Q|��]����%��?�D}����һE��ڇMo-b8��ٚ	(�x"kRUc�]ul�ᒳH
��g�e�R����
3�(JXݳ���W�YH���9��U��ڲ�y�H���������v �I[�4����Y0�l���8f��M0ٜ2����x��[9���@����/Un��̗�i�	 g��%��Ħ�vU	��/�����7:^��m}Q��`j��	(Q� �шk���w��kU�S�N�^�*JBK+q U��G��)t�i���0EΈE�L�+�=�]r�~�hn/8h]�N���^��ғ��	E�5OhN���Q�A��cF�.W�lk��z��|$:0`-(X�&U{o�i���G�����I� ����`�S�˲צ�Gȇ��&�u���n����QJ����s=Mrj������˞R8R�n��"���Ai�=}̽y����rȉ�&��a>8��q�AI�6*���;�,����NHE@��:a��;%�N�,p��ǘuu�/GL�2���x5j@���a���ɸ �0�+^��׬�jz�T_Ѷ� ���Q�~���j5N���"��yEN�B��f"؃@��j�w�r~l;�O��֙vW�I��!��>Q�#xB��|J�Fry`�!\!�h������d��"�3����܄OL�㍤]�g���&9_r�������;]0�H7^s[�OS�>O�7���`��s��m��	�A3R	�%3��Vb�ߜ��O�7��rYV|�/*M>�'3�ߌH?K|(�J� ȹ1�
9�mi���ջ����Fo'������٫@�Q�QKG(8�ńlj�b�����z^��z���^�~�ūO/ڥE��ާ|�+p�-v�j�����
�c��%�S*�An�z�ɋ������X���=p�a�B���k��K�0r����uLZ0(��oq-��W��Y�G~�7+v7��7�5��:����j|j�z�1�����7/�xf���oj�Z��ֶb�u�x�����i�x��
9R��\��;4�P�N��ں�c5�D=f��{��OM�3��?�9A'������W��[;�g͝V7��9㎾xɝ���MT��r~�i��Ϭ�0�2�׽ę+�/�:���G&��W�c�'Տ<����aZ�;�p�B-�:������7o�����V��=R��ˀ`�J���b�db��k�Cke_	��nT�|Ǫ����]��ֲ]�U�xL.E����"_��cH����k{�5	*AYE�"�%��ʟ;O#��w�B��W;-G�X,܀a�5a�&n5u~k|<q���[~w�R��r*�~�	�Z���ۭ��l6����ˎ|9#<���pW���y�>Y��.v�;JaQ��2&EL<�0�E�_=��	cT�4:��­��%��x���B�_�`� b�G�x�yr����~[ؿ�j��'hxL��h߱Gٱ��'����.+8�8�p�ϗP����������������`��#z�t�
�_�z9��I�W���f���������ŗ�u��߱�6��t��	��R�&w��?*��j�?r(�-<sk�L@�T��WL��kOU�p� ����w�����N%�@m��y���A>��hBH\p�I��	@�D=�l�}[���*�K�2���g%���� e�O�i��G����^�fܕ�)t�|���b��P�q�pm���o3(1���������p �Z�a�2M����jw��JA�$� ��̋"=�ξy�₃���}u�+��șgz؍95F�Pj�鮹���h,�I�l�nD�>��"^XXrB�A��X`��<D_LfuP,^3R(�phm�_�I��݄�:�:�Y}zg�M7��
�6Q �O+��-���wh��:j�t9F�Zy<B�6*�a����c�"�~t��ï1J��C��~�E�R��}�1O���ne�%�ɠH����H�A^�����F��"�	�O�=Tp@G�L�'@�+?�T�; z����0h=U�����J�d.�x�.-�%(��$�έ��A�.�]�$��$c�*Ѩ��l#��W)4���hͬ )�����zy���г�[4�AT�lIZ4ɶ�H�����xk��	�Uo�8>?sӫ���~�����1�1��O{��|E�gvK:�$r�gG�s_��t�V+� ��65fyu�a��WK)9���o)�QO'9y��t"�������a	:!�X�Yh��Kg��e�_}�H|�r��C�!���T���������lW0B���l�Q�|��Kx$�;%|LC� �`�k�pҕ��tQ#���7ك�p�����]ͧ(
�F�.��٣h'D�?�0��}B0XS���	�!��g�z36�=y���۵J��r1�]m�'�[i).�˜ Iq]�5��e��_����5����VNp�tg�FS�_�/�����[<z� �2�{��V��>��Z{s��?R-�L�Uw�߃��x�Tt`����^��slҿ|�������Y�m}�n(��$hiĉ
�;C�a'�f���L��Z!���H��7蔐�@���k�&�mm3�|�=�V^?������v�G͹ͯ�+KTr��W�\7�6��M~RKա�Z8�2R���%�)c�����5�p��?�U�O�#�RAh�r@T��B�Y �= n�����bR\!"�uq\6�άœ��X��яIS�#��WQ�z,��o�O�;;2"
�\�J�;�SӢE2z�xao�lh��|M:H�aE�QOH࠹��/�[�!���b��(q�Z��n��]���Q�R4�����<P�|4�C;;l�no�`6�
�I��(��4|V�C��2�	F��ޡ�q#.D<`���,�R�� �ܰ��Cc��Z� K /|��<�6�s�G�������ٞ�H��$��>��e�H�pF����j��G��e�͋�_��-��I`���5!�?�C��%���c��M�:�7�����Oe͡�b����}v6�`,p�@�3dQ(��n�T�O�e��o>*���v��Q�ӂ<$д"Η��EY��g�c�*����:�?�g]���rfۏ`XR��J`��wH���n��&<�I��}=-��o����
C#��Q����G����gs�O)kk�n(I����D���'|'w1����&8c���)-=�z�.��	hj\�$�[�׋�8�4�L'}������"�lO0Gh\a����W�v`���o|�&�|���&�|vۥ�J`K����8��,ɩK{�3�g�5A!W%�":2���n�8����[��O���[�F(8���H效�����l��^�O�Om��v�^�-����`}��9X?�z�������`���RM̜�dl�K������-�!	<ig8蚳��c�&4�,����-a*8�-Øx�5܆�.o1E:/����U�����
0]:4�k�]x�[[��T���� �eB�h1V��K.������=[�=2���a���5Ǆ��-��J{$Z+������t�̘������ntQ$�<�z�`�� �ך��LI��n�\ V���!�0�j�c�t�:ا���?u��V�j̥(��Om���h�ΫW2w������w�@�R�Y���8萤W�v�rM�M���v�hG>2���g��������NH�����|iTWtU0E�|��6RҒ��ϊ�B���;J$�A���rp��;6���4 ��u�)+��=b�UT�Qs�*,6}%R�z�z"eS��_r�&�cD�n��pu�J�3$�ӲByF��H�p[<J��������!m�T�0�|�s���O���n?��������vk)�6N���O^�#nM�����7h/}���X�1k;(Q�D�$�o���*��� �D�GX�b�<D���$�?���*��Ȑ���w��j6d�ja�է��y��|	KGXYP֗D�\���
lU}Q�mԉ/���2�@��C��^\���X2������+��{ٗ����|w�I�3Kb��8�j�7c��T��bs�h�8�E;��
SJw&�'\p�0�J�h��SR`�-�W�:�ۃ�G�Q`�j�"�'4}�ef!:�W(5L;gZ�]Z������0����<K��$ׄ�ꌸAm�p!���;���R���^һ~�Y�1��P�JD^>/�����>�P�m��l�G�Az�Ve�%6�4���}vXvŴ����%��?��3�_t��%�kŞ)+).Tюrwgvc(�JE��Mq��Uh�4Vd��kPSe��#b<Md������WP��|�f�eʎ�6w����Q���+�D5��S�nu��e�An4�փ����G:
�S��<Pu�YO�8�l�b���OE\Q���ط��H�wk��>�g�k4����@R�`��X�84�j��t7�)=���]�]w���o���ʆbOSq=��$v%�Pt	Q3����VWq�Tx�cF���9�����ް�2����h��jU#:���u,���q������W�M�!Z�!D��΢ۮ��;�
�x_�����6���*5:��w}(�@���D̼��?�A,��;����� ��+%"�"�W��ǒ���?��P�JtH>��:~]Rk���Pl�f�/��;Y�:�r}�����M�f:�9���#�`T�w����>�UR��è��J�W��]y øC��kI3�W������������d�M�So�� _���ɷ�g*��)#Uj}d�t��}���K�zv@l,t^3G��W
��1�XhN��,6ɺ��e*��Y��%w`��O��Ӳ��K?�i�hՏ"T<���)\���%$���0d�~������0��9U�
�-�Y'���]̊C�nf'�6�3�z\���$��W��pq�Z'\�7.�,�������@�0��$��+��W�z�����]��g��I�zenӐNV��k㧤�#��-���_X$.M�L�i���MW�a!��u{�<N&�����>�1�>���7��"9�)�ۥ���Р$��Zb�!���j����.��_�x�E9��/m�}k;o��؆��%v]8�1<��4</�؉?��pW�o�A֛�-;3ArF�5i!*�f�2�,/�}P�P�zB=.�x������QK�;��&T>�x����`��������e�g�c�}y��p��P���d;�ɍ&��q�H�xGz!�qE�`Buf�B_�t�+۟��vS^�>���O�[Rtsug��0�ԋ�Y�f�1F�Gr@��HKCE�1�,nھ�6ݷ����N#��nZ������ca���ePl�Ã��ʋ�v��"�� ���gtj���ju���;���B���1�%B:��[,9��h4�at���A�Vzv�����>�%*(9��)s>K�5�8x�����&�0TeN@�/l#@�21X�����
�6E��a.=��7�2
��cja_rhŶM]��u�9�*j8�[�����4܊)�H^�q�.d")���^ʠ�W6��/W�B�~~7Fb�����U��ȃ��p80����F?�꼐����/]��Ȏر�:h|�v�}Rp��y[̙�A1���h;RL�z����p)�N�\����6uM��[�#Rn������\� Q�!��!X�JR)"�h��s���Q?�.�e0��6I�i�X@�R�ZnP>Z͏vv�n�݅���&8m�i,	�֗`_<�~R��\��լ�Eh�'ΩJ9^�\�K������~p	�ݼ�)~R@L��_6��ŭ+�Gm�4�5�2��cJ�������czm,������`)Aݗ���~]c,����H�-,�Tf���C����m\�B�K��|e#X;l��\d����S�eXs5���jU����?�Ļ��b�KP��c=��ȝٷ�)r!�YW�Ԙ���8,ևvo�"�4���~��!���+X�攖Bs�����Z(M�e�}�d��,X��^�t�
���Jy��P�+ڭ�=��Oe]{$�t��������:��HvJn���Db`�&!Q$����)$>�����2��g��y J�"[8�Xuyhh��u�/�9�}�7��������.��}��Q�
~���BKms��?�*{��q��Q��,R���2hB��&۫��JjZQ�mҳ��g����]?�1��v����ˬ��,�Fcx�I�E�\3���:��Qs���;�bO�4�Ce$�;���̑t���*�����{l��w�ĿC��q���t�9/*62�����芟<��<&�j��޸���<�R�,�=l^Y����OL1Y.����
J��՝�74������2)bI��:B%��#���~���ݘ�ϩ�Ki�eߕ�d[�iZ\��Z��n݃3a �s�l-q8���?t�Sǿ3G��O�kʗ.(zd��������]�8Ҹ�SK�_��P0'�qsך��=����]�x�8�x>����/Z�,Wv�J��BmPV�"�eF���2�����c���m��f�[`\j�v�"��L�;s��Xm����B�������.@�9��õu�.Vم��}��,;����	�9����]����N�:.�}H�(�?-�9��$& �&��ȝ��~�������9
1��Bh���4���0����Kp%GC�&�x�[��ߓ�OB�d'�r|�lP"�:���f���K|a�;����j�̊�(z���z[��`��1��A;��a�~�a���O]2s��;�[D�>�!�6��P4%+�5v��s��"��i���+�NuG^�4�bU�J{�2ju2~��H3�-\O���}���(b�a�_u�K�	��>�r#3���yǬ԰4�V��DOJ�t��?�]}P�ݙ0,UN]�Yo�*#l�B���&v�&���P�_�B�f�H�i�HZY>����@�GI���l��	����w�V�&��')یEF0-���ڙ�jf
�Lc���{��Z� ���f �Wnw�0�Nū�x��^� h \��/�c~�i���BkA�Ԏt���z�����b���}� ,�Z�.��.����/W��z��w��[�fǪ����Vw�4��v�;~��߸|���ʌ]�qG����>)F����}�r��zu�y������p��vU�����\J�$y��F*��6�9��_��$Z�Sp����c$=M*�l`��ty�����c9X��3���љ���\��\����*��n���;��r���>�d��F�ȉ�5�f���~
�@��U&���rmKu�G�hDŌ&��!���mԦ�P���	�e�j��(BV�a)�,���@�|�4���{�"�I�	7��EO?�kM�1�]���e�b%"�?w�\*�di�l�.3�T.-2%�U�8ʜ��,4��1��	�_��e��>��(����*�Yco�WB��^��Ҁp�I�R��r?�r��L�8�Ј�)��~:��6�UB0���'�a?3(�9��e"�C�q
-
��j���V�;�>�O��HS������_�g��4V� |Y��6���K�݃��R;�o�Bz�`����fD�[��("5�ַi�#!�n�?L^�{i������iD�q���!R�Df$�b��X�f*���a��/-�A0�Uٺc�_�5�g |F�6KQ��sb�5�ꯓ�	�r?�����r���Ps<���T Ѝ#�q́�^�nL2E�=�Xy�~��S[�I�ߓO0g�"��� )��Bߞ��'����������R���B E&�����<�f2-�� Ԣ;oK����k9�oޕ?�6�H@����D	W�6���R�z��0�Le��$)�ܐ��mx����YP�PDO���]@gYm�#y-�k�Z������]���->������B�э�G�m��}�˽�ۑ�B�-�����F���|R8R�^���}�;#���m�
�R�;G-L|�WIeX�]'bhY���z��_9�omz��Rx��ގKy���:�%�^��~�ݸEF�s�|qm���ߚ[�8�NRO4�=V�����Phu:;X����S8s]��ԗ�E��M��/^�y�4G�9[�� ^7Rjm^�Y��y���%�;P����[�S�'%��p�,���oT�-�u��{��r�u"#����ɕ� ���`��2Jq��*�g��-s����	��i����e��� ����˝���j�A|����Ի���5y��W	Mdz�\R�\��Yf���z$P�˙	j~x@sV�a?�J�/­�|b�f�f��М� ���@�m5#jt�G���L�;&�Q׫�]v��6���0��Hc"=��(#���C#{Mj^!�n*�.�ӘO/���S �� 7���Q�:��.G�>�n{���d~(S�T@-����
s����U&�dTJ��Cv?Ҧ��*q�xtf_R���el��F^$�c��R���"Uۊk������	�r�	��3����v��t�U�'c߀�{t����r�]����h&�
j�)>�[X��Ԁ-H�G����ů	M�U�����E��~�|�Sd�g���m���>��L�z17�hn"�*!g�C��I;Dv���r�_ދ�'V�dU�Ba�癞$����E��_㺚g�r�;��\��l���756�\!0rwr�5�I��s�P^�V�HO�x!�$��'����CbBZ��)=��)����hG(�.�Kr]��*��l�{N��
\	����[[�����Ë5e��b��S�KΓ�ˎLIecP�dH���c�o��ʿD���0A]�^r�j�QꔙJ/�+p<'�4�����I���VQ���Lz�I���5{��o���D�BB�P%�:�"1�X*<�����L͞���F%SU��U�x�'�
Q�������.:`����O��A:�6N�xPU	`�ݙ�G!fa�z^�+s��I� Б"C�!�Yِg8�au��*����X�6<Xr��gI��3@g ���Ɍ/m;�6����C�P.#h�&�p�j!s��M�U>�ۼƤ�� p*7	��%"R� o�6���!��`�R��!�k�8��9�h�/}!`��*�A��w�, QF'Z�@���'��6����b�񜷊���5Q�B�+�6�Jɯ�Ӈ@����"+�B�iU<����h��Fx���JY�P���hk�<�><+6�q���е��ʻ}/���lN9��R���Hm��1��Oɶ�6�BF�r�p��A�vp�*�2J��iBH����01�����(�d�Ռ����S�\<���us�Ʒ�'��EtH�^��WfӜLJ�I��#t3����H�Y��k��(,�h��(�V
_b��!gY��K��m���9�!G�"Z�<��6�������s���x�6��	�,��y������տ�k�1�Zs�;ƥ|�G�3�]�����%�8�p��zgA��2�vOтO��3{� B�A>iy��J��$ä�鴳���9p�{2,�7�7�Pj�}󅿔�K�wV'��%�_�����y��ɦ8?��m������D�]BRZ1;�3�������Qs+�ծ���X>�� v$Qؑ2Yz�xU7�~��Pp�V�A�B	�wR�*_i��U��	�(fb���G�E6V��XӨ�
�n鮵�{����:�/���w�V�Ư������������:Ywq˄m&h]�xX�
�vф4�@��7��a+&�U�!�'[���.܈�f���v�s�igo�	���0L_�m���<�Y�fz���}g!#����022K�n4�P��7Km���nO<2x��!�|>�=e�1�k�oj ��X��doe�ۏd*�X\��8}�6�}��ib�)�fZ��C���GU����/ Vȴ���ު����_M�vi�p�>��Ynj-��su���q{²�B��C0H`�z[��r��ǅ��c�KN��3F������!�*���c��Mq�����a��� �.,�� ��{}�����{�T��U�ǎ.��*��>'��SL8����%�M�QUӉ`�':���>2E|��E$�X�>�c}4ˡ�$�+VX39���7��:!OQ�q�|�ܒ�I����In���<*���;��o����h�6�(�p�_��Gɣ����U�@e��1�:=�f�%-���S�m��v���ay�]�O��*�i.�˒�qu>�=��[�]�j'd���8猐M�U^q�(u������6Y������P����H�b�py�&G2O��B:}� �\,ޫ�=H���P	2�F�5��q�)b�m��߷W���/6����?����KнQ�P@~d��i�t}.O� "���P�mڜ�IE�c��Hj�_fP��t��WA�J��tg+��"�tA��su��a��]�uT�v�����qU�g��Dk��VǒYLBQ�2���v��|4�77:�]Ggi��4=!f��|��-��&%0��D8,����V���e�0����o��y?����2.J-�k��7U"˖U:���gȓ=m4����(x!�T�"��������F].��Q�q�iTg����ۅe�%�;���i��-x�i���M`��)�`!�:�^�q,#����C�O�q�����h��M�YNz0L*Khh����/�n��h��{{�b��;S�p{6�g�6!N((v��9���oo��\O߬�~�"���R}�fF5,Fv��aݰ�����z{��fZ[%������xq`�OL�Ok�T�Z���j�~i��k)z�1Q���F̺���o"��s3>_[����7/�ʹ��c��(H�������x�]Y���O�C䫬���c�j�#W�BO�4D�m�������Q'}����"6�vnߥ��Y���k�����Y��)V��h����Rs�ْ���`6YD�ᮡ�fxܳ���Y-
����/4l� @H}g��>яY�I·�ib2� �,�=�m��ӭ=��/t�mb��|K,Vc;��R(�ٰ�[^$����%�F�����{��QlҞ��o0�Pg�� -�t�Ƕ����(��-�)�l�Cx=��܈����l�z�׋o�T��S�}#���� Άg��}�1�\��n�;�^c����P�yV�y7��Bk��z"���L��\���Q�יO+hy{3�	H�����?v������2q�|u���O��Z��l���ǰ��ЄTqz��ޓ��n�ڼ(F��*0���SC�I�>u�Up��B���C=@�@ d)�!�O�ch���Y�.+]��L �G�:K?b�����������`��oÿ��3�f��@�rU�\Ҍj�z&��x��U�����~[����H� zˬrf�j���{���Vg
���tօ7t5@����v�2v�����T�֘U|���E#[��`Σ��54o~.Ճ��㖠���2�V�BXF��-`�<k�)����Cȅ�̳a�ʂmon��o�_���.��Nu��~�� ;.w�T���ER�:�h�o��a���63X��W��V	��\�%�a� sT1�3�Έ	[��'I��b��ٔ>��g��;�_�&"[v�wv^�/�O�vk\��l�z��y%N1�/�F'⦟HLc~���$�&'BM��]���9��om#������D1����Ք�X�k������SӡC��C:^{�K�U��~ח��$������[[-,j�]�̭W+���� �D�|h4�1k
���u�yY)�9�S��
r5�Ω������榥*�_7��/��7f ������{Q1�.z%�1��V�,
ʯ���J��܉?��J0gS'Nl:����*FН��8*��C����������ה�(�/@�i�myx�-.���I=G��l1$�ɭ�͈� ����Iz��x���[9�hx1J��A:ǎ�7�[_l}`i�}/k�a�Q֎B"b���.� ��k<=���:z���] '� ���o<��ߏCד!a7/�D���U��VE�<���q��MNݝ���t��V�ܘ��,�Ns,�S��nL�>����6;L�\��ԡκ�Pj����dep9���$8� �9,�H�H�jY���3�U�p����1�B�A�+�����I��ܒ>2A5d�Y��#N��ʉ	Ooc%¯mi��(B�h���H��0�m�S4��]2T��c�@l�"8�uB�����-�pQj)=��h����r�^�wHR/.���U���1���SS�T����I��k���bX��>8S@�������p��n��u^'��i*�yU�^~��;��~w��ϐة��@$ϥ��3l��ǡ��Ev�Z$K`C`����[����
���H����T/�9I����4�hH������"�PI2_,��N}�'e����Wȷg�����){���,����O3�r�,��t[���p�&f��ۓ���g����C̷�������1�tJ�#2�s�kq/���jI�w؎B�~ѐҗX�dYz x��zc�ʑNF���_5R�).լ�D�D[�#�2̤Ǧ�@B�A^�0B�!j��NO~�߳W���1ڟ}�D����P?-7	���c�~[$� �Qj�G%�Cm�s�z���םhň���i�ڠ#�23s�g��=�+��S �|w="�9L�[��^�]�����h@a��!�����}l����ҁ	���u�Z�)MF���Q����~�@ZP�Ȏ�V9�8�cD����޶�"	�WƜ�ةr����M���c+B�73 �Dkt_ֹ���
�"�>����g�O��� s�C����mO�\��q;��]xLG���E�e%�c�PV+�/��ԣ�`�[ȡM�/��6�>Z��,����[F��Y�B��6���d&�d3@`jd�_ ��Vֈ�����l�����1	�&E�YKm:�Q��f����ZUe��]��e�h�Zi0i���f`-h��tJ	&3)H��g��|�Ot��<2&����)��ږ�ro$}�����HkIaϦ{�W������X�T�G��9�v�P��d�ַ�&@�W '��P�aZ�F�����74CK��*�v��Q�}�D'2�K�o���=C��-�Yq�weû،�9��U;Q��v-����!�o4̌�0F��j'1�}Q
��c{��8,�䝾��E4��.�q�ޏ�،�^�����$���$oпjr��գ[p`�����p'O�Bɒ������!����M��ا�}�F�=�s��y�r�DJ��d���Q��W�lnV���P�e�l�g��,K2H���dm5�O����G�=��b<t��U������ֿ��>�B��-gI9ohc�h�L�PV��C�>�b �+����/@B���d�e�����tb�qc	�^�@��#�}���@y:"���eE#G�\��#J�͡2���i�W��8���c����M�)7�l˹-����wO���5�S�մ��+j �l�ut,�yK���}Ȃ_��,�}�k���6���&�h.މO)q�Z�"�?��oO�)��I���]Mv�4��D�;�g��j�<F�ei��v��):���j�~6jy�@+.����CKũ���>;���{q9�8w.a-�`	s�Y(��Т讽�($�t���R��?�6�xc�?(G-�sZ��WU���E�jى�B �k��FH��@V�*��4��88���b����G�r�_�����W��Fd ��K��"�R@�{1f����z٫� >0L}"���9$���:�𤥤n�����Xh�t�^��D�ғ���!{��+�������{-[ӥ��J/!al��_b��sj��Tclp���'�EX>��U�#��]�J���9�d�s	3�{H_5������l�L�vw[�=���]h.an����U�;��˴��<x�'����_�w~�Y7�����m�l���݅����U������z@7S}Qs�_�/u$� @$�kΰ�wy��")2��	���CҚ6��S���×����YC���ُ���x�����2y(*踖�!��O�K�Oh��^<=w��< ���2���{��Ud������mm ~8z	�MI�v�wbJ�\��Q����\Ez����S�^
>0�}���������%n�a@ъ�899i�>9���0Dh�����b�8�\~oT��*V|�_L���]�&�uV-i�����VF��=.�7�	\��Ex?�_'Ty�ԓ��CL�n;��P��1��v<%���{}y*ia �69?�1٘N��
螙�j�x�<O��W�x���\�I�c���̾�TM�KGH"4���~廒I�%d��T�aC��QJ�j��k6�+6o�����ս��Z� ��R��q�:��1�3�G��:[�}�����;��Zc�J�v�t���%�𘺶��ۍ`�M�_B���D���ܻ�O�5��e���EL�l�O���q�`��7@������V���7]{no���f������e4*�/&���C;G����u�y����C�6S���M*j�e�>l��A�y7��\r%"4���	�R�V����9��>gҠY_Z��_�ԩҐXDMxiYAhf+��{.�xY��){	�N�����s�$��s��Ce�+̶x��q��*����̞�w�C;x�a�i9q`����׫��h��6�Z�҃z�R��x�T�ޗҁ�[q�ۅ�֗i4m�@uV����D�q��@�4���-��]�I{o��ǫ��.��Sb\\(/1 ?AU8O�G��v�I-.Y����]�bA*��޾�
u�I�A���h��nuU���	s�&�<Ju����%F����j�{'����BҼv����oQ�+'[��"��ho�
�zn����=��D����VB����Gk��$�މo�Q��߮����~3�����`�Z�H4*"��^��)[�,��&9)	P��\=�� v3�〷Gl�3A�98�7�@���r�u|�3� ����Ҙ֊���/�-�bV�aH{���Ȁ��G ��ȳ��@�s(9�
�n�n.����Q:�O��z��,n����W9�5����wfO��Sk0�1_�IE�C���p��L���������\&���I����'��؈�]�|:�xZ@����2,p5Ö�25|@��6�ۙ�h���^De��f��k�W�X�TI�z�@&��4r��-nc�2�.���`6�u�%]6�M�B���v@�k�9d�Ļ_H{�������*���֡��aS�Q�Ҷ���&Ky�j(Z)�ej�k�5������!ȗդVb��w���c*���0)4��������
q(��v&���%\��AN��i��1�oe^��aɦ���Z�?]����E%ǃ�RdyD���ď��Ǜ�e9��xҶx8������C���na�'� D���k�Oc���Df�X���kZ������ � <�J$��Gp�d�}�8"̀iX�W��j���p�m~3On;P64��BK$_Z��&Lǘ�f��,` O��rg\_�p��9�l��5!H%�t0�_*6߶M����7��$J!0�	o��Ũ�GL :d��Z�D��p����U{��58b�MQ��K�`Rn�$��6�B-ҘYL�y�g��"�c+x�X�UYB P3ݢ���r�ϓ�i�f�T�#\ժU��N�#���������4ʢX���P�y��Rw���Lⶆ�^���ٟ�N��1�r1O��WF97��DDnx�}�[��SF��3�h�zs�=����m:?��ݝ�Z�Lo�h��>Ǯ���e�1�k��z���3;I���W��=���K�<8!q����y.b]Tu�َ��ۯ�`�w���QhEY�e��<���(�6Z&t�Z�v1]m��+��\ ��Um��,����WZ��h|U�q7������IH�:<A?�g�|��^�l�|�i�wQ��ꊠ(R�1�n�ۊ�;��ڤ���]I!�s������� ��ox7�yP%���Qn\J|lK�  gԽL�?�z�����ސZг�v����T�g����L����Lx� �R���XO���I�u@��D�9��w\�\rT�Y͐ܥZ��|����&\*5��;�&J{o��*��U�p�p��>t6��P~N��D�3�A��D��4��I[4����� |4��-��Q��<��T����e�����Beּ5�|�w~���}6�G6Z�'_�e\��-�Z�p���#Jح��7�tc��`Ǭ�?��&d�)8��en}�!P!z]�wu�i3�3yJt>)K�47ME@���Z��r�ұ��z����R�v,47�f�끖�0��E��?��2a��t�d�5(�S9K�h�Ϭ��~�tT_9�=Dw>��r�@��4��-�k(��su