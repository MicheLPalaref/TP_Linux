��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�q���4]oHe��zL!��Qo���r���d�Lݠ��%yl�/�1 oJ�'�nT��ָ��T�:p>c�Y�-�2b�x��(@�KH6�fH5yM���m��ljr@�Gu�<7�t�I��M�MX�9����˺��G��q��	%���q��m4�N�ˠ����� q�s�e޶����y��	'���u
lc0�Ӓ�Ŧ��}�.睩�1r�ry8��[w=��4�J �m�s��:��G����x�_����t�G��!�.��IBp�8cx�eK�C}4d�J��,�꺊,��К%X�@a,�:�{o
�In��)x>������������U�;/�_�Ng�:!�w2�U�A<�C��^>/���$;���Dx�6��ROZ�+m_\��񫃧Ƕ�(y�'2χ���C6��V^ۑ�H!C]��T\�B�9x��������3���R���BG�%��_�n�,�R��/��u�k*h:�r��TE~�B�	���\%7�!P�P��JToyE���wYZ�ܭH,c켝vz�R��݅�6v�e�xJI�����>#��X����c���?Bt�R?�N6y��9�vAA�Svl��Xk,��f���6�i���'��F���Op��+Vlקjö&�Z�}IQ�6,"�UD0_�K�Cl{�l�Wkkz��/bG��<�������"X����j�F^f��cf"���r��}���Cr��|T�����,�;X�&n:\: