// DE10_Standard_Qsys.v

// Generated using ACDS version 16.1 200

`timescale 1 ps / 1 ps
module DE10_Standard_Qsys (
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_clk,            //      alt_vip_cl_cvi_0_clocked_video.vid_clk
		input  wire [7:0]  alt_vip_cl_cvi_0_clocked_video_vid_data,           //                                    .vid_data
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_de,             //                                    .vid_de
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_datavalid,      //                                    .vid_datavalid
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_locked,         //                                    .vid_locked
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_f,              //                                    .vid_f
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_v_sync,         //                                    .vid_v_sync
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_h_sync,         //                                    .vid_h_sync
		input  wire [7:0]  alt_vip_cl_cvi_0_clocked_video_vid_color_encoding, //                                    .vid_color_encoding
		input  wire [7:0]  alt_vip_cl_cvi_0_clocked_video_vid_bit_width,      //                                    .vid_bit_width
		output wire        alt_vip_cl_cvi_0_clocked_video_sof,                //                                    .sof
		output wire        alt_vip_cl_cvi_0_clocked_video_sof_locked,         //                                    .sof_locked
		output wire        alt_vip_cl_cvi_0_clocked_video_refclk_div,         //                                    .refclk_div
		output wire        alt_vip_cl_cvi_0_clocked_video_clipping,           //                                    .clipping
		output wire        alt_vip_cl_cvi_0_clocked_video_padding,            //                                    .padding
		output wire        alt_vip_cl_cvi_0_clocked_video_overflow,           //                                    .overflow
		input  wire        alt_vip_itc_mtlc_clocked_video_vid_clk,            //      alt_vip_itc_mtlc_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_mtlc_clocked_video_vid_data,           //                                    .vid_data
		output wire        alt_vip_itc_mtlc_clocked_video_underflow,          //                                    .underflow
		output wire        alt_vip_itc_mtlc_clocked_video_vid_datavalid,      //                                    .vid_datavalid
		output wire        alt_vip_itc_mtlc_clocked_video_vid_v_sync,         //                                    .vid_v_sync
		output wire        alt_vip_itc_mtlc_clocked_video_vid_h_sync,         //                                    .vid_h_sync
		output wire        alt_vip_itc_mtlc_clocked_video_vid_f,              //                                    .vid_f
		output wire        alt_vip_itc_mtlc_clocked_video_vid_h,              //                                    .vid_h
		output wire        alt_vip_itc_mtlc_clocked_video_vid_v,              //                                    .vid_v
		output wire        audio_avalon_controller_conduit_end_CLK,           // audio_avalon_controller_conduit_end.CLK
		output wire        audio_avalon_controller_conduit_end_LRCIN,         //                                    .LRCIN
		output wire        audio_avalon_controller_conduit_end_DIN,           //                                    .DIN
		output wire        audio_avalon_controller_conduit_end_LRCOUT,        //                                    .LRCOUT
		input  wire        audio_avalon_controller_conduit_end_DOUT,          //                                    .DOUT
		output wire        audio_avalon_controller_conduit_end_BCLK,          //                                    .BCLK
		output wire        av_i2c_clk_pio_external_connection_export,         //  av_i2c_clk_pio_external_connection.export
		inout  wire        av_i2c_data_pio_external_connection_export,        // av_i2c_data_pio_external_connection.export
		input  wire [3:0]  button_pio_external_connection_export,             //      button_pio_external_connection.export
		input  wire        clk_clk,                                           //                                 clk.clk
		output wire        clk_mtlc_clk,                                      //                            clk_mtlc.clk
		output wire        clk_sdram_clk,                                     //                           clk_sdram.clk
		output wire        clk_sys_clk,                                       //                             clk_sys.clk
		output wire [3:0]  led_pio_external_connection_export,                //         led_pio_external_connection.export
		output wire        pll_0_locked_export,                               //                        pll_0_locked.export
		input  wire        reset_reset_n,                                     //                               reset.reset_n
		output wire [12:0] sdram_wire_addr,                                   //                          sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                     //                                    .ba
		output wire        sdram_wire_cas_n,                                  //                                    .cas_n
		output wire        sdram_wire_cke,                                    //                                    .cke
		output wire        sdram_wire_cs_n,                                   //                                    .cs_n
		inout  wire [15:0] sdram_wire_dq,                                     //                                    .dq
		output wire [1:0]  sdram_wire_dqm,                                    //                                    .dqm
		output wire        sdram_wire_ras_n,                                  //                                    .ras_n
		output wire        sdram_wire_we_n,                                   //                                    .we_n
		output wire        td_reset_pio_external_connection_export,           //    td_reset_pio_external_connection.export
		inout  wire        touch_i2c_opencores_export_scl_pad_io,             //          touch_i2c_opencores_export.scl_pad_io
		inout  wire        touch_i2c_opencores_export_sda_pad_io,             //                                    .sda_pad_io
		input  wire        touch_int_n_external_connection_export             //     touch_int_n_external_connection.export
	);

	wire         alt_vip_vfr_0_avalon_streaming_source_valid;                      // alt_vip_vfr_0:dout_valid -> alt_vip_cl_mixer_0:din1_valid
	wire  [23:0] alt_vip_vfr_0_avalon_streaming_source_data;                       // alt_vip_vfr_0:dout_data -> alt_vip_cl_mixer_0:din1_data
	wire         alt_vip_vfr_0_avalon_streaming_source_ready;                      // alt_vip_cl_mixer_0:din1_ready -> alt_vip_vfr_0:dout_ready
	wire         alt_vip_vfr_0_avalon_streaming_source_startofpacket;              // alt_vip_vfr_0:dout_startofpacket -> alt_vip_cl_mixer_0:din1_startofpacket
	wire         alt_vip_vfr_0_avalon_streaming_source_endofpacket;                // alt_vip_vfr_0:dout_endofpacket -> alt_vip_cl_mixer_0:din1_endofpacket
	wire         alt_vip_cl_vfb_0_dout_valid;                                      // alt_vip_cl_vfb_0:dout_valid -> alt_vip_cl_crs_0:din_valid
	wire  [15:0] alt_vip_cl_vfb_0_dout_data;                                       // alt_vip_cl_vfb_0:dout_data -> alt_vip_cl_crs_0:din_data
	wire         alt_vip_cl_vfb_0_dout_ready;                                      // alt_vip_cl_crs_0:din_ready -> alt_vip_cl_vfb_0:dout_ready
	wire         alt_vip_cl_vfb_0_dout_startofpacket;                              // alt_vip_cl_vfb_0:dout_startofpacket -> alt_vip_cl_crs_0:din_startofpacket
	wire         alt_vip_cl_vfb_0_dout_endofpacket;                                // alt_vip_cl_vfb_0:dout_endofpacket -> alt_vip_cl_crs_0:din_endofpacket
	wire         alt_vip_cl_crs_0_dout_valid;                                      // alt_vip_cl_crs_0:dout_valid -> alt_vip_cl_csc_0:din_valid
	wire  [23:0] alt_vip_cl_crs_0_dout_data;                                       // alt_vip_cl_crs_0:dout_data -> alt_vip_cl_csc_0:din_data
	wire         alt_vip_cl_crs_0_dout_ready;                                      // alt_vip_cl_csc_0:din_ready -> alt_vip_cl_crs_0:dout_ready
	wire         alt_vip_cl_crs_0_dout_startofpacket;                              // alt_vip_cl_crs_0:dout_startofpacket -> alt_vip_cl_csc_0:din_startofpacket
	wire         alt_vip_cl_crs_0_dout_endofpacket;                                // alt_vip_cl_crs_0:dout_endofpacket -> alt_vip_cl_csc_0:din_endofpacket
	wire         alt_vip_cl_mixer_0_dout_valid;                                    // alt_vip_cl_mixer_0:dout_valid -> alt_vip_cts_0:din_valid
	wire  [23:0] alt_vip_cl_mixer_0_dout_data;                                     // alt_vip_cl_mixer_0:dout_data -> alt_vip_cts_0:din_data
	wire         alt_vip_cl_mixer_0_dout_ready;                                    // alt_vip_cts_0:din_ready -> alt_vip_cl_mixer_0:dout_ready
	wire         alt_vip_cl_mixer_0_dout_startofpacket;                            // alt_vip_cl_mixer_0:dout_startofpacket -> alt_vip_cts_0:din_startofpacket
	wire         alt_vip_cl_mixer_0_dout_endofpacket;                              // alt_vip_cl_mixer_0:dout_endofpacket -> alt_vip_cts_0:din_endofpacket
	wire         alt_vip_clip_0_dout_valid;                                        // alt_vip_clip_0:dout_valid -> alt_vip_scl_0:din_valid
	wire  [23:0] alt_vip_clip_0_dout_data;                                         // alt_vip_clip_0:dout_data -> alt_vip_scl_0:din_data
	wire         alt_vip_clip_0_dout_ready;                                        // alt_vip_scl_0:din_ready -> alt_vip_clip_0:dout_ready
	wire         alt_vip_clip_0_dout_startofpacket;                                // alt_vip_clip_0:dout_startofpacket -> alt_vip_scl_0:din_startofpacket
	wire         alt_vip_clip_0_dout_endofpacket;                                  // alt_vip_clip_0:dout_endofpacket -> alt_vip_scl_0:din_endofpacket
	wire         alt_vip_cl_csc_0_dout_valid;                                      // alt_vip_cl_csc_0:dout_valid -> alt_vip_clip_0:din_valid
	wire  [23:0] alt_vip_cl_csc_0_dout_data;                                       // alt_vip_cl_csc_0:dout_data -> alt_vip_clip_0:din_data
	wire         alt_vip_cl_csc_0_dout_ready;                                      // alt_vip_clip_0:din_ready -> alt_vip_cl_csc_0:dout_ready
	wire         alt_vip_cl_csc_0_dout_startofpacket;                              // alt_vip_cl_csc_0:dout_startofpacket -> alt_vip_clip_0:din_startofpacket
	wire         alt_vip_cl_csc_0_dout_endofpacket;                                // alt_vip_cl_csc_0:dout_endofpacket -> alt_vip_clip_0:din_endofpacket
	wire         alt_vip_clip_1_dout_valid;                                        // alt_vip_clip_1:dout_valid -> alt_vip_cl_vfb_0:din_valid
	wire  [15:0] alt_vip_clip_1_dout_data;                                         // alt_vip_clip_1:dout_data -> alt_vip_cl_vfb_0:din_data
	wire         alt_vip_clip_1_dout_ready;                                        // alt_vip_cl_vfb_0:din_ready -> alt_vip_clip_1:dout_ready
	wire         alt_vip_clip_1_dout_startofpacket;                                // alt_vip_clip_1:dout_startofpacket -> alt_vip_cl_vfb_0:din_startofpacket
	wire         alt_vip_clip_1_dout_endofpacket;                                  // alt_vip_clip_1:dout_endofpacket -> alt_vip_cl_vfb_0:din_endofpacket
	wire         alt_vip_cl_dil_0_dout_valid;                                      // alt_vip_cl_dil_0:dout_valid -> alt_vip_clip_1:din_valid
	wire  [15:0] alt_vip_cl_dil_0_dout_data;                                       // alt_vip_cl_dil_0:dout_data -> alt_vip_clip_1:din_data
	wire         alt_vip_cl_dil_0_dout_ready;                                      // alt_vip_clip_1:din_ready -> alt_vip_cl_dil_0:dout_ready
	wire         alt_vip_cl_dil_0_dout_startofpacket;                              // alt_vip_cl_dil_0:dout_startofpacket -> alt_vip_clip_1:din_startofpacket
	wire         alt_vip_cl_dil_0_dout_endofpacket;                                // alt_vip_cl_dil_0:dout_endofpacket -> alt_vip_clip_1:din_endofpacket
	wire         alt_vip_cl_clp_1_dout_valid;                                      // alt_vip_cl_clp_1:dout_valid -> alt_vip_itc_mtlc:is_valid
	wire  [23:0] alt_vip_cl_clp_1_dout_data;                                       // alt_vip_cl_clp_1:dout_data -> alt_vip_itc_mtlc:is_data
	wire         alt_vip_cl_clp_1_dout_ready;                                      // alt_vip_itc_mtlc:is_ready -> alt_vip_cl_clp_1:dout_ready
	wire         alt_vip_cl_clp_1_dout_startofpacket;                              // alt_vip_cl_clp_1:dout_startofpacket -> alt_vip_itc_mtlc:is_sop
	wire         alt_vip_cl_clp_1_dout_endofpacket;                                // alt_vip_cl_clp_1:dout_endofpacket -> alt_vip_itc_mtlc:is_eop
	wire         alt_vip_cts_0_dout_valid;                                         // alt_vip_cts_0:dout_valid -> alt_vip_cl_clp_1:din_valid
	wire  [23:0] alt_vip_cts_0_dout_data;                                          // alt_vip_cts_0:dout_data -> alt_vip_cl_clp_1:din_data
	wire         alt_vip_cts_0_dout_ready;                                         // alt_vip_cl_clp_1:din_ready -> alt_vip_cts_0:dout_ready
	wire         alt_vip_cts_0_dout_startofpacket;                                 // alt_vip_cts_0:dout_startofpacket -> alt_vip_cl_clp_1:din_startofpacket
	wire         alt_vip_cts_0_dout_endofpacket;                                   // alt_vip_cts_0:dout_endofpacket -> alt_vip_cl_clp_1:din_endofpacket
	wire         alt_vip_scl_0_dout_valid;                                         // alt_vip_scl_0:dout_valid -> alt_vip_cl_mixer_0:din0_valid
	wire  [23:0] alt_vip_scl_0_dout_data;                                          // alt_vip_scl_0:dout_data -> alt_vip_cl_mixer_0:din0_data
	wire         alt_vip_scl_0_dout_ready;                                         // alt_vip_cl_mixer_0:din0_ready -> alt_vip_scl_0:dout_ready
	wire         alt_vip_scl_0_dout_startofpacket;                                 // alt_vip_scl_0:dout_startofpacket -> alt_vip_cl_mixer_0:din0_startofpacket
	wire         alt_vip_scl_0_dout_endofpacket;                                   // alt_vip_scl_0:dout_endofpacket -> alt_vip_cl_mixer_0:din0_endofpacket
	wire         alt_vip_cl_cps_0_dout_0_valid;                                    // alt_vip_cl_cps_0:dout_0_valid -> alt_vip_cl_dil_0:din_valid
	wire  [15:0] alt_vip_cl_cps_0_dout_0_data;                                     // alt_vip_cl_cps_0:dout_0_data -> alt_vip_cl_dil_0:din_data
	wire         alt_vip_cl_cps_0_dout_0_ready;                                    // alt_vip_cl_dil_0:din_ready -> alt_vip_cl_cps_0:dout_0_ready
	wire         alt_vip_cl_cps_0_dout_0_startofpacket;                            // alt_vip_cl_cps_0:dout_0_startofpacket -> alt_vip_cl_dil_0:din_startofpacket
	wire         alt_vip_cl_cps_0_dout_0_endofpacket;                              // alt_vip_cl_cps_0:dout_0_endofpacket -> alt_vip_cl_dil_0:din_endofpacket
	wire         alt_vip_cl_cvi_0_dout_0_valid;                                    // alt_vip_cl_cvi_0:dout_0_valid -> alt_vip_cl_cps_0:din_0_valid
	wire   [7:0] alt_vip_cl_cvi_0_dout_0_data;                                     // alt_vip_cl_cvi_0:dout_0_data -> alt_vip_cl_cps_0:din_0_data
	wire         alt_vip_cl_cvi_0_dout_0_ready;                                    // alt_vip_cl_cps_0:din_0_ready -> alt_vip_cl_cvi_0:dout_0_ready
	wire         alt_vip_cl_cvi_0_dout_0_startofpacket;                            // alt_vip_cl_cvi_0:dout_0_startofpacket -> alt_vip_cl_cps_0:din_0_startofpacket
	wire         alt_vip_cl_cvi_0_dout_0_endofpacket;                              // alt_vip_cl_cvi_0:dout_0_endofpacket -> alt_vip_cl_cps_0:din_0_endofpacket
	wire  [31:0] alt_vip_vfr_0_avalon_master_readdata;                             // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire         alt_vip_vfr_0_avalon_master_waitrequest;                          // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire  [31:0] alt_vip_vfr_0_avalon_master_address;                              // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire         alt_vip_vfr_0_avalon_master_read;                                 // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire         alt_vip_vfr_0_avalon_master_readdatavalid;                        // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire   [6:0] alt_vip_vfr_0_avalon_master_burstcount;                           // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                             // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                             // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                                 // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                              // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                    // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                   // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                               // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                         // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                          // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                             // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         alt_vip_cl_vfb_0_mem_master_rd_waitrequest;                       // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_waitrequest -> alt_vip_cl_vfb_0:mem_master_rd_waitrequest
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_rd_readdata;                          // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_readdata -> alt_vip_cl_vfb_0:mem_master_rd_readdata
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_rd_address;                           // alt_vip_cl_vfb_0:mem_master_rd_address -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_address
	wire         alt_vip_cl_vfb_0_mem_master_rd_read;                              // alt_vip_cl_vfb_0:mem_master_rd_read -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_read
	wire         alt_vip_cl_vfb_0_mem_master_rd_readdatavalid;                     // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_readdatavalid -> alt_vip_cl_vfb_0:mem_master_rd_readdatavalid
	wire   [6:0] alt_vip_cl_vfb_0_mem_master_rd_burstcount;                        // alt_vip_cl_vfb_0:mem_master_rd_burstcount -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_burstcount
	wire         alt_vip_cl_vfb_0_mem_master_wr_waitrequest;                       // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_waitrequest -> alt_vip_cl_vfb_0:mem_master_wr_waitrequest
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_wr_address;                           // alt_vip_cl_vfb_0:mem_master_wr_address -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_address
	wire   [3:0] alt_vip_cl_vfb_0_mem_master_wr_byteenable;                        // alt_vip_cl_vfb_0:mem_master_wr_byteenable -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_byteenable
	wire         alt_vip_cl_vfb_0_mem_master_wr_write;                             // alt_vip_cl_vfb_0:mem_master_wr_write -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_write
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_wr_writedata;                         // alt_vip_cl_vfb_0:mem_master_wr_writedata -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_writedata
	wire   [6:0] alt_vip_cl_vfb_0_mem_master_wr_burstcount;                        // alt_vip_cl_vfb_0:mem_master_wr_burstcount -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_burstcount
	wire         alt_vip_cts_0_master_waitrequest;                                 // mm_interconnect_0:alt_vip_cts_0_master_waitrequest -> alt_vip_cts_0:master_waitrequest
	wire  [31:0] alt_vip_cts_0_master_address;                                     // alt_vip_cts_0:master_address -> mm_interconnect_0:alt_vip_cts_0_master_address
	wire  [31:0] alt_vip_cts_0_master_writedata;                                   // alt_vip_cts_0:master_writedata -> mm_interconnect_0:alt_vip_cts_0_master_writedata
	wire         alt_vip_cts_0_master_write;                                       // alt_vip_cts_0:master_write -> mm_interconnect_0:alt_vip_cts_0_master_write
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                 // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                 // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata;            // alt_vip_vfr_0:slave_readdata -> mm_interconnect_0:alt_vip_vfr_0_avalon_slave_readdata
	wire   [4:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address;             // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire         mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read;                // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire         mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write;               // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire  [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata;           // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire         mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_chipselect;  // mm_interconnect_0:touch_i2c_opencores_avalon_slave_0_chipselect -> touch_i2c_opencores:wb_stb_i
	wire   [7:0] mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_readdata;    // touch_i2c_opencores:wb_dat_o -> mm_interconnect_0:touch_i2c_opencores_avalon_slave_0_readdata
	wire         mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_waitrequest; // touch_i2c_opencores:wb_ack_o -> mm_interconnect_0:touch_i2c_opencores_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_address;     // mm_interconnect_0:touch_i2c_opencores_avalon_slave_0_address -> touch_i2c_opencores:wb_adr_i
	wire         mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_write;       // mm_interconnect_0:touch_i2c_opencores_avalon_slave_0_write -> touch_i2c_opencores:wb_we_i
	wire   [7:0] mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_writedata;   // mm_interconnect_0:touch_i2c_opencores_avalon_slave_0_writedata -> touch_i2c_opencores:wb_dat_i
	wire  [31:0] mm_interconnect_0_alt_vip_scl_0_control_readdata;                 // alt_vip_scl_0:control_readdata -> mm_interconnect_0:alt_vip_scl_0_control_readdata
	wire         mm_interconnect_0_alt_vip_scl_0_control_waitrequest;              // alt_vip_scl_0:control_waitrequest -> mm_interconnect_0:alt_vip_scl_0_control_waitrequest
	wire   [6:0] mm_interconnect_0_alt_vip_scl_0_control_address;                  // mm_interconnect_0:alt_vip_scl_0_control_address -> alt_vip_scl_0:control_address
	wire         mm_interconnect_0_alt_vip_scl_0_control_read;                     // mm_interconnect_0:alt_vip_scl_0_control_read -> alt_vip_scl_0:control_read
	wire   [3:0] mm_interconnect_0_alt_vip_scl_0_control_byteenable;               // mm_interconnect_0:alt_vip_scl_0_control_byteenable -> alt_vip_scl_0:control_byteenable
	wire         mm_interconnect_0_alt_vip_scl_0_control_readdatavalid;            // alt_vip_scl_0:control_readdatavalid -> mm_interconnect_0:alt_vip_scl_0_control_readdatavalid
	wire         mm_interconnect_0_alt_vip_scl_0_control_write;                    // mm_interconnect_0:alt_vip_scl_0_control_write -> alt_vip_scl_0:control_write
	wire  [31:0] mm_interconnect_0_alt_vip_scl_0_control_writedata;                // mm_interconnect_0:alt_vip_scl_0_control_writedata -> alt_vip_scl_0:control_writedata
	wire  [31:0] mm_interconnect_0_alt_vip_clip_0_control_readdata;                // alt_vip_clip_0:control_readdata -> mm_interconnect_0:alt_vip_clip_0_control_readdata
	wire         mm_interconnect_0_alt_vip_clip_0_control_waitrequest;             // alt_vip_clip_0:control_waitrequest -> mm_interconnect_0:alt_vip_clip_0_control_waitrequest
	wire   [2:0] mm_interconnect_0_alt_vip_clip_0_control_address;                 // mm_interconnect_0:alt_vip_clip_0_control_address -> alt_vip_clip_0:control_address
	wire         mm_interconnect_0_alt_vip_clip_0_control_read;                    // mm_interconnect_0:alt_vip_clip_0_control_read -> alt_vip_clip_0:control_read
	wire   [3:0] mm_interconnect_0_alt_vip_clip_0_control_byteenable;              // mm_interconnect_0:alt_vip_clip_0_control_byteenable -> alt_vip_clip_0:control_byteenable
	wire         mm_interconnect_0_alt_vip_clip_0_control_readdatavalid;           // alt_vip_clip_0:control_readdatavalid -> mm_interconnect_0:alt_vip_clip_0_control_readdatavalid
	wire         mm_interconnect_0_alt_vip_clip_0_control_write;                   // mm_interconnect_0:alt_vip_clip_0_control_write -> alt_vip_clip_0:control_write
	wire  [31:0] mm_interconnect_0_alt_vip_clip_0_control_writedata;               // mm_interconnect_0:alt_vip_clip_0_control_writedata -> alt_vip_clip_0:control_writedata
	wire  [31:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_readdata;            // alt_vip_cl_mixer_0:control_readdata -> mm_interconnect_0:alt_vip_cl_mixer_0_control_readdata
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_waitrequest;         // alt_vip_cl_mixer_0:control_waitrequest -> mm_interconnect_0:alt_vip_cl_mixer_0_control_waitrequest
	wire   [6:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_address;             // mm_interconnect_0:alt_vip_cl_mixer_0_control_address -> alt_vip_cl_mixer_0:control_address
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_read;                // mm_interconnect_0:alt_vip_cl_mixer_0_control_read -> alt_vip_cl_mixer_0:control_read
	wire   [3:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_byteenable;          // mm_interconnect_0:alt_vip_cl_mixer_0_control_byteenable -> alt_vip_cl_mixer_0:control_byteenable
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_readdatavalid;       // alt_vip_cl_mixer_0:control_readdatavalid -> mm_interconnect_0:alt_vip_cl_mixer_0_control_readdatavalid
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_write;               // mm_interconnect_0:alt_vip_cl_mixer_0_control_write -> alt_vip_cl_mixer_0:control_write
	wire  [31:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_writedata;           // mm_interconnect_0:alt_vip_cl_mixer_0_control_writedata -> alt_vip_cl_mixer_0:control_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                   // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                    // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;          // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;       // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                    // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                      // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                       // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                         // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                     // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_led_pio_s1_chipselect;                          // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                            // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                             // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_write;                               // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                           // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_0_button_pio_s1_chipselect;                       // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                         // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                          // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_write;                            // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                        // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire         mm_interconnect_0_av_i2c_clk_pio_s1_chipselect;                   // mm_interconnect_0:av_i2c_clk_pio_s1_chipselect -> av_i2c_clk_pio:chipselect
	wire  [31:0] mm_interconnect_0_av_i2c_clk_pio_s1_readdata;                     // av_i2c_clk_pio:readdata -> mm_interconnect_0:av_i2c_clk_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_av_i2c_clk_pio_s1_address;                      // mm_interconnect_0:av_i2c_clk_pio_s1_address -> av_i2c_clk_pio:address
	wire         mm_interconnect_0_av_i2c_clk_pio_s1_write;                        // mm_interconnect_0:av_i2c_clk_pio_s1_write -> av_i2c_clk_pio:write_n
	wire  [31:0] mm_interconnect_0_av_i2c_clk_pio_s1_writedata;                    // mm_interconnect_0:av_i2c_clk_pio_s1_writedata -> av_i2c_clk_pio:writedata
	wire         mm_interconnect_0_av_i2c_data_pio_s1_chipselect;                  // mm_interconnect_0:av_i2c_data_pio_s1_chipselect -> av_i2c_data_pio:chipselect
	wire  [31:0] mm_interconnect_0_av_i2c_data_pio_s1_readdata;                    // av_i2c_data_pio:readdata -> mm_interconnect_0:av_i2c_data_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_av_i2c_data_pio_s1_address;                     // mm_interconnect_0:av_i2c_data_pio_s1_address -> av_i2c_data_pio:address
	wire         mm_interconnect_0_av_i2c_data_pio_s1_write;                       // mm_interconnect_0:av_i2c_data_pio_s1_write -> av_i2c_data_pio:write_n
	wire  [31:0] mm_interconnect_0_av_i2c_data_pio_s1_writedata;                   // mm_interconnect_0:av_i2c_data_pio_s1_writedata -> av_i2c_data_pio:writedata
	wire         mm_interconnect_0_td_reset_pio_s1_chipselect;                     // mm_interconnect_0:td_reset_pio_s1_chipselect -> td_reset_pio:chipselect
	wire  [31:0] mm_interconnect_0_td_reset_pio_s1_readdata;                       // td_reset_pio:readdata -> mm_interconnect_0:td_reset_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_td_reset_pio_s1_address;                        // mm_interconnect_0:td_reset_pio_s1_address -> td_reset_pio:address
	wire         mm_interconnect_0_td_reset_pio_s1_write;                          // mm_interconnect_0:td_reset_pio_s1_write -> td_reset_pio:write_n
	wire  [31:0] mm_interconnect_0_td_reset_pio_s1_writedata;                      // mm_interconnect_0:td_reset_pio_s1_writedata -> td_reset_pio:writedata
	wire         mm_interconnect_0_audio_avalon_controller_s1_chipselect;          // mm_interconnect_0:audio_avalon_controller_s1_chipselect -> audio_avalon_controller:avs_s1_cs_n
	wire  [31:0] mm_interconnect_0_audio_avalon_controller_s1_readdata;            // audio_avalon_controller:avs_s1_readdata -> mm_interconnect_0:audio_avalon_controller_s1_readdata
	wire   [2:0] mm_interconnect_0_audio_avalon_controller_s1_address;             // mm_interconnect_0:audio_avalon_controller_s1_address -> audio_avalon_controller:avs_s1_addr
	wire         mm_interconnect_0_audio_avalon_controller_s1_read;                // mm_interconnect_0:audio_avalon_controller_s1_read -> audio_avalon_controller:avs_s1_read_n
	wire         mm_interconnect_0_audio_avalon_controller_s1_begintransfer;       // mm_interconnect_0:audio_avalon_controller_s1_begintransfer -> audio_avalon_controller:avs_s1_begintransfer
	wire         mm_interconnect_0_audio_avalon_controller_s1_write;               // mm_interconnect_0:audio_avalon_controller_s1_write -> audio_avalon_controller:avs_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_avalon_controller_s1_writedata;           // mm_interconnect_0:audio_avalon_controller_s1_writedata -> audio_avalon_controller:avs_s1_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                            // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                              // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                           // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                               // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                  // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                            // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                         // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                 // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                             // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_touch_int_n_s1_chipselect;                      // mm_interconnect_0:touch_int_n_s1_chipselect -> touch_int_n:chipselect
	wire  [31:0] mm_interconnect_0_touch_int_n_s1_readdata;                        // touch_int_n:readdata -> mm_interconnect_0:touch_int_n_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_int_n_s1_address;                         // mm_interconnect_0:touch_int_n_s1_address -> touch_int_n:address
	wire         mm_interconnect_0_touch_int_n_s1_write;                           // mm_interconnect_0:touch_int_n_s1_write -> touch_int_n:write_n
	wire  [31:0] mm_interconnect_0_touch_int_n_s1_writedata;                       // mm_interconnect_0:touch_int_n_s1_writedata -> touch_int_n:writedata
	wire  [31:0] mm_interconnect_0_alt_vip_cts_0_slave_readdata;                   // alt_vip_cts_0:slave_readdata -> mm_interconnect_0:alt_vip_cts_0_slave_readdata
	wire   [4:0] mm_interconnect_0_alt_vip_cts_0_slave_address;                    // mm_interconnect_0:alt_vip_cts_0_slave_address -> alt_vip_cts_0:slave_address
	wire         mm_interconnect_0_alt_vip_cts_0_slave_read;                       // mm_interconnect_0:alt_vip_cts_0_slave_read -> alt_vip_cts_0:slave_read
	wire         mm_interconnect_0_alt_vip_cts_0_slave_write;                      // mm_interconnect_0:alt_vip_cts_0_slave_write -> alt_vip_cts_0:slave_write
	wire  [31:0] mm_interconnect_0_alt_vip_cts_0_slave_writedata;                  // mm_interconnect_0:alt_vip_cts_0_slave_writedata -> alt_vip_cts_0:slave_writedata
	wire         irq_mapper_receiver0_irq;                                         // alt_vip_vfr_0:slave_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                         // alt_vip_cts_0:status_update_int -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                                         // button_pio:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                         // jtag_uart:av_irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                         // sys_clk_timer:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                             // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver2_irq;                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                    // touch_i2c_opencores:wb_inta_o -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver6_irq;                                         // irq_synchronizer_001:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                // touch_int_n:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver7_irq;                                         // irq_synchronizer_002:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                // audio_avalon_controller:avs_s1_irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [alt_vip_cl_clp_1:main_reset, alt_vip_cl_cps_0:main_reset, alt_vip_cl_crs_0:main_reset, alt_vip_cl_csc_0:main_reset, alt_vip_cl_cvi_0:main_reset_reset, alt_vip_cl_dil_0:av_st_reset, alt_vip_cl_mixer_0:main_reset_reset, alt_vip_cl_vfb_0:main_reset, alt_vip_cl_vfb_0:mem_reset, alt_vip_clip_0:main_reset, alt_vip_clip_1:main_reset, alt_vip_cts_0:reset, alt_vip_itc_mtlc:rst, alt_vip_scl_0:main_reset, alt_vip_vfr_0:master_reset, alt_vip_vfr_0:reset, av_i2c_clk_pio:reset_n, av_i2c_data_pio:reset_n, button_pio:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_0:alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram:reset_n, sys_clk_timer:reset_n, sysid:reset_n, td_reset_pio:reset_n]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                           // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [audio_avalon_controller:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, mm_interconnect_0:touch_i2c_opencores_clock_reset_reset_bridge_in_reset_reset, touch_i2c_opencores:wb_rst_i, touch_int_n:reset_n]

	DE10_Standard_Qsys_alt_vip_cl_clp_1 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (3),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_IN_WIDTH                 (800),
		.MAX_IN_HEIGHT                (480),
		.CLIPPING_METHOD              ("RECTANGLE"),
		.LEFT_OFFSET                  (0),
		.RIGHT_OFFSET                 (0),
		.TOP_OFFSET                   (0),
		.BOTTOM_OFFSET                (0),
		.RECTANGLE_WIDTH              (800),
		.RECTANGLE_HEIGHT             (480),
		.USER_PACKET_SUPPORT          ("PASSTHROUGH"),
		.RUNTIME_CONTROL              (0),
		.LIMITED_READBACK             (0)
	) alt_vip_cl_clp_1 (
		.main_clock         (clk_sys_clk),                         // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cts_0_dout_data),             //        din.data
		.din_valid          (alt_vip_cts_0_dout_valid),            //           .valid
		.din_startofpacket  (alt_vip_cts_0_dout_startofpacket),    //           .startofpacket
		.din_endofpacket    (alt_vip_cts_0_dout_endofpacket),      //           .endofpacket
		.din_ready          (alt_vip_cts_0_dout_ready),            //           .ready
		.dout_data          (alt_vip_cl_clp_1_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_clp_1_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_clp_1_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_clp_1_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_clp_1_dout_ready)          //           .ready
	);

	DE10_Standard_Qsys_alt_vip_cl_cps_0 #(
		.BITS_PER_SYMBOL     (8),
		.USER_PACKET_SUPPORT ("PASSTHROUGH")
	) alt_vip_cl_cps_0 (
		.main_clock           (clk_sys_clk),                           // main_clock.clk
		.main_reset           (rst_controller_reset_out_reset),        // main_reset.reset
		.din_0_data           (alt_vip_cl_cvi_0_dout_0_data),          //      din_0.data
		.din_0_valid          (alt_vip_cl_cvi_0_dout_0_valid),         //           .valid
		.din_0_startofpacket  (alt_vip_cl_cvi_0_dout_0_startofpacket), //           .startofpacket
		.din_0_endofpacket    (alt_vip_cl_cvi_0_dout_0_endofpacket),   //           .endofpacket
		.din_0_ready          (alt_vip_cl_cvi_0_dout_0_ready),         //           .ready
		.dout_0_data          (alt_vip_cl_cps_0_dout_0_data),          //     dout_0.data
		.dout_0_valid         (alt_vip_cl_cps_0_dout_0_valid),         //           .valid
		.dout_0_startofpacket (alt_vip_cl_cps_0_dout_0_startofpacket), //           .startofpacket
		.dout_0_endofpacket   (alt_vip_cl_cps_0_dout_0_endofpacket),   //           .endofpacket
		.dout_0_ready         (alt_vip_cl_cps_0_dout_0_ready)          //           .ready
	);

	DE10_Standard_Qsys_alt_vip_cl_crs_0 alt_vip_cl_crs_0 (
		.main_clock         (clk_sys_clk),                         // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_vfb_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_vfb_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_vfb_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_vfb_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_vfb_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_cl_crs_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_crs_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_crs_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_crs_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_crs_0_dout_ready)          //           .ready
	);

	DE10_Standard_Qsys_alt_vip_cl_csc_0 alt_vip_cl_csc_0 (
		.main_clock         (clk_sys_clk),                         // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_crs_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_crs_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_crs_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_crs_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_crs_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_cl_csc_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_csc_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_csc_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_csc_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_csc_0_dout_ready)          //           .ready
	);

	DE10_Standard_Qsys_alt_vip_cl_cvi_0 #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (2),
		.COLOUR_PLANES_ARE_IN_PARALLEL (0),
		.SYNC_TO                       (0),
		.MATCH_CTRLDATA_PKT_CLIP_BASIC (0),
		.MATCH_CTRLDATA_PKT_PAD_ADV    (0),
		.OVERFLOW_HANDLING             (0),
		.USE_EMBEDDED_SYNCS            (1),
		.USE_HDMI_DEPRICATION          (0),
		.GENERATE_VID_F                (0),
		.USE_STD                       (0),
		.STD_WIDTH                     (1),
		.GENERATE_ANC                  (0),
		.ANC_DEPTH                     (1),
		.EXTRACT_TOTAL_RESOLUTION      (1),
		.INTERLACED                    (1),
		.H_ACTIVE_PIXELS_F0            (720),
		.V_ACTIVE_LINES_F0             (288),
		.V_ACTIVE_LINES_F1             (288),
		.FIFO_DEPTH                    (2048),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0)
	) alt_vip_cl_cvi_0 (
		.main_clock_clk                   (clk_sys_clk),                                       //    main_clock.clk
		.main_reset_reset                 (rst_controller_reset_out_reset),                    //    main_reset.reset
		.dout_0_data                      (alt_vip_cl_cvi_0_dout_0_data),                      //        dout_0.data
		.dout_0_valid                     (alt_vip_cl_cvi_0_dout_0_valid),                     //              .valid
		.dout_0_startofpacket             (alt_vip_cl_cvi_0_dout_0_startofpacket),             //              .startofpacket
		.dout_0_endofpacket               (alt_vip_cl_cvi_0_dout_0_endofpacket),               //              .endofpacket
		.dout_0_ready                     (alt_vip_cl_cvi_0_dout_0_ready),                     //              .ready
		.clocked_video_vid_clk            (alt_vip_cl_cvi_0_clocked_video_vid_clk),            // clocked_video.vid_clk
		.clocked_video_vid_data           (alt_vip_cl_cvi_0_clocked_video_vid_data),           //              .vid_data
		.clocked_video_vid_de             (alt_vip_cl_cvi_0_clocked_video_vid_de),             //              .vid_de
		.clocked_video_vid_datavalid      (alt_vip_cl_cvi_0_clocked_video_vid_datavalid),      //              .vid_datavalid
		.clocked_video_vid_locked         (alt_vip_cl_cvi_0_clocked_video_vid_locked),         //              .vid_locked
		.clocked_video_vid_f              (alt_vip_cl_cvi_0_clocked_video_vid_f),              //              .vid_f
		.clocked_video_vid_v_sync         (alt_vip_cl_cvi_0_clocked_video_vid_v_sync),         //              .vid_v_sync
		.clocked_video_vid_h_sync         (alt_vip_cl_cvi_0_clocked_video_vid_h_sync),         //              .vid_h_sync
		.clocked_video_vid_color_encoding (alt_vip_cl_cvi_0_clocked_video_vid_color_encoding), //              .vid_color_encoding
		.clocked_video_vid_bit_width      (alt_vip_cl_cvi_0_clocked_video_vid_bit_width),      //              .vid_bit_width
		.clocked_video_sof                (alt_vip_cl_cvi_0_clocked_video_sof),                //              .sof
		.clocked_video_sof_locked         (alt_vip_cl_cvi_0_clocked_video_sof_locked),         //              .sof_locked
		.clocked_video_refclk_div         (alt_vip_cl_cvi_0_clocked_video_refclk_div),         //              .refclk_div
		.clocked_video_clipping           (alt_vip_cl_cvi_0_clocked_video_clipping),           //              .clipping
		.clocked_video_padding            (alt_vip_cl_cvi_0_clocked_video_padding),            //              .padding
		.clocked_video_overflow           (alt_vip_cl_cvi_0_clocked_video_overflow)            //              .overflow
	);

	DE10_Standard_Qsys_alt_vip_cl_dil_0 #(
		.MAX_WIDTH                        (720),
		.MAX_HEIGHT                       (576),
		.USER_PACKET_SUPPORT              ("PASSTHROUGH"),
		.USER_PACKET_FIFO_DEPTH           (0),
		.PIXELS_IN_PARALLEL               (1),
		.BITS_PER_SYMBOL                  (8),
		.NUMBER_OF_COLOR_PLANES           (2),
		.COLOR_PLANES_ARE_IN_PARALLEL     (1),
		.IS_422                           (1),
		.IS_YCBCR                         (1),
		.DEINTERLACE_ALGORITHM            ("BOB"),
		.MOTION_BLEED                     (1),
		.RUNTIME_CONTROL                  (0),
		.MOTION_BPS                       (7),
		.CADENCE_DETECTION                (0),
		.CADENCE_ALGORITHM_NAME           ("CADENCE_32_22_VOF"),
		.CLOCKS_ARE_SEPARATE              (0),
		.MEM_PORT_WIDTH                   (256),
		.WRITE_MASTER_FIFO_DEPTH          (64),
		.WRITE_MASTER_BURST_TARGET        (32),
		.EDI_READ_MASTER_FIFO_DEPTH       (64),
		.EDI_READ_MASTER_BURST_TARGET     (32),
		.MA_READ_MASTER_FIFO_DEPTH        (64),
		.MA_READ_MASTER_BURST_TARGET      (32),
		.MOTION_WRITE_MASTER_FIFO_DEPTH   (64),
		.MOTION_WRITE_MASTER_BURST_TARGET (32),
		.MOTION_READ_MASTER_FIFO_DEPTH    (64),
		.MOTION_READ_MASTER_BURST_TARGET  (32),
		.MEM_BASE_ADDR                    (0)
	) alt_vip_cl_dil_0 (
		.av_st_clock        (clk_sys_clk),                           // av_st_clock.clk
		.av_st_reset        (rst_controller_reset_out_reset),        // av_st_reset.reset
		.din_data           (alt_vip_cl_cps_0_dout_0_data),          //         din.data
		.din_valid          (alt_vip_cl_cps_0_dout_0_valid),         //            .valid
		.din_startofpacket  (alt_vip_cl_cps_0_dout_0_startofpacket), //            .startofpacket
		.din_endofpacket    (alt_vip_cl_cps_0_dout_0_endofpacket),   //            .endofpacket
		.din_ready          (alt_vip_cl_cps_0_dout_0_ready),         //            .ready
		.dout_data          (alt_vip_cl_dil_0_dout_data),            //        dout.data
		.dout_valid         (alt_vip_cl_dil_0_dout_valid),           //            .valid
		.dout_startofpacket (alt_vip_cl_dil_0_dout_startofpacket),   //            .startofpacket
		.dout_endofpacket   (alt_vip_cl_dil_0_dout_endofpacket),     //            .endofpacket
		.dout_ready         (alt_vip_cl_dil_0_dout_ready)            //            .ready
	);

	DE10_Standard_Qsys_alt_vip_cl_mixer_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_WIDTH                    (800),
		.MAX_HEIGHT                   (480),
		.IS_422                       (1),
		.USER_PACKET_SUPPORT          ("DISCARD"),
		.USER_PACKET_FIFO_DEPTH       (0)
	) alt_vip_cl_mixer_0 (
		.main_clock_clk        (clk_sys_clk),                                                // main_clock.clk
		.main_reset_reset      (rst_controller_reset_out_reset),                             // main_reset.reset
		.din0_data             (alt_vip_scl_0_dout_data),                                    //       din0.data
		.din0_valid            (alt_vip_scl_0_dout_valid),                                   //           .valid
		.din0_startofpacket    (alt_vip_scl_0_dout_startofpacket),                           //           .startofpacket
		.din0_endofpacket      (alt_vip_scl_0_dout_endofpacket),                             //           .endofpacket
		.din0_ready            (alt_vip_scl_0_dout_ready),                                   //           .ready
		.din1_data             (alt_vip_vfr_0_avalon_streaming_source_data),                 //       din1.data
		.din1_valid            (alt_vip_vfr_0_avalon_streaming_source_valid),                //           .valid
		.din1_startofpacket    (alt_vip_vfr_0_avalon_streaming_source_startofpacket),        //           .startofpacket
		.din1_endofpacket      (alt_vip_vfr_0_avalon_streaming_source_endofpacket),          //           .endofpacket
		.din1_ready            (alt_vip_vfr_0_avalon_streaming_source_ready),                //           .ready
		.dout_data             (alt_vip_cl_mixer_0_dout_data),                               //       dout.data
		.dout_valid            (alt_vip_cl_mixer_0_dout_valid),                              //           .valid
		.dout_startofpacket    (alt_vip_cl_mixer_0_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (alt_vip_cl_mixer_0_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (alt_vip_cl_mixer_0_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_0_alt_vip_cl_mixer_0_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_0_alt_vip_cl_mixer_0_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_0_alt_vip_cl_mixer_0_control_write),         //           .write
		.control_writedata     (mm_interconnect_0_alt_vip_cl_mixer_0_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_0_alt_vip_cl_mixer_0_control_read),          //           .read
		.control_readdata      (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_alt_vip_cl_mixer_0_control_waitrequest)    //           .waitrequest
	);

	DE10_Standard_Qsys_alt_vip_cl_vfb_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.READY_LATENCY                (1),
		.MAX_WIDTH                    (720),
		.MAX_HEIGHT                   (480),
		.CLOCKS_ARE_SEPARATE          (1),
		.MEM_PORT_WIDTH               (32),
		.MEM_BASE_ADDR                (16777216),
		.BURST_ALIGNMENT              (1),
		.WRITE_FIFO_DEPTH             (512),
		.WRITE_BURST_TARGET           (64),
		.READ_FIFO_DEPTH              (512),
		.READ_BURST_TARGET            (64),
		.WRITER_RUNTIME_CONTROL       (0),
		.READER_RUNTIME_CONTROL       (0),
		.IS_FRAME_WRITER              (0),
		.IS_FRAME_READER              (0),
		.DROP_FRAMES                  (1),
		.REPEAT_FRAMES                (1),
		.DROP_REPEAT_USER             (1),
		.INTERLACED_SUPPORT           (0),
		.CONTROLLED_DROP_REPEAT       (0),
		.DROP_INVALID_FIELDS          (1),
		.MULTI_FRAME_DELAY            (1),
		.IS_SYNC_MASTER               (0),
		.IS_SYNC_SLAVE                (0),
		.USER_PACKETS_MAX_STORAGE     (0),
		.MAX_SYMBOLS_PER_PACKET       (10),
		.NUM_BUFFERS                  (3)
	) alt_vip_cl_vfb_0 (
		.main_clock                  (clk_sys_clk),                                  //    main_clock.clk
		.main_reset                  (rst_controller_reset_out_reset),               //    main_reset.reset
		.mem_clock                   (clk_sys_clk),                                  //     mem_clock.clk
		.mem_reset                   (rst_controller_reset_out_reset),               //     mem_reset.reset
		.din_data                    (alt_vip_clip_1_dout_data),                     //           din.data
		.din_valid                   (alt_vip_clip_1_dout_valid),                    //              .valid
		.din_startofpacket           (alt_vip_clip_1_dout_startofpacket),            //              .startofpacket
		.din_endofpacket             (alt_vip_clip_1_dout_endofpacket),              //              .endofpacket
		.din_ready                   (alt_vip_clip_1_dout_ready),                    //              .ready
		.mem_master_wr_address       (alt_vip_cl_vfb_0_mem_master_wr_address),       // mem_master_wr.address
		.mem_master_wr_burstcount    (alt_vip_cl_vfb_0_mem_master_wr_burstcount),    //              .burstcount
		.mem_master_wr_waitrequest   (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),   //              .waitrequest
		.mem_master_wr_write         (alt_vip_cl_vfb_0_mem_master_wr_write),         //              .write
		.mem_master_wr_writedata     (alt_vip_cl_vfb_0_mem_master_wr_writedata),     //              .writedata
		.mem_master_wr_byteenable    (alt_vip_cl_vfb_0_mem_master_wr_byteenable),    //              .byteenable
		.dout_data                   (alt_vip_cl_vfb_0_dout_data),                   //          dout.data
		.dout_valid                  (alt_vip_cl_vfb_0_dout_valid),                  //              .valid
		.dout_startofpacket          (alt_vip_cl_vfb_0_dout_startofpacket),          //              .startofpacket
		.dout_endofpacket            (alt_vip_cl_vfb_0_dout_endofpacket),            //              .endofpacket
		.dout_ready                  (alt_vip_cl_vfb_0_dout_ready),                  //              .ready
		.mem_master_rd_address       (alt_vip_cl_vfb_0_mem_master_rd_address),       // mem_master_rd.address
		.mem_master_rd_burstcount    (alt_vip_cl_vfb_0_mem_master_rd_burstcount),    //              .burstcount
		.mem_master_rd_waitrequest   (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),   //              .waitrequest
		.mem_master_rd_read          (alt_vip_cl_vfb_0_mem_master_rd_read),          //              .read
		.mem_master_rd_readdata      (alt_vip_cl_vfb_0_mem_master_rd_readdata),      //              .readdata
		.mem_master_rd_readdatavalid (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid)  //              .readdatavalid
	);

	DE10_Standard_Qsys_alt_vip_clip_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (3),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_IN_WIDTH                 (720),
		.MAX_IN_HEIGHT                (480),
		.CLIPPING_METHOD              ("RECTANGLE"),
		.LEFT_OFFSET                  (0),
		.RIGHT_OFFSET                 (10),
		.TOP_OFFSET                   (0),
		.BOTTOM_OFFSET                (10),
		.RECTANGLE_WIDTH              (720),
		.RECTANGLE_HEIGHT             (480),
		.USER_PACKET_SUPPORT          ("PASSTHROUGH"),
		.RUNTIME_CONTROL              (1),
		.LIMITED_READBACK             (0)
	) alt_vip_clip_0 (
		.main_clock            (clk_sys_clk),                                            // main_clock.clk
		.main_reset            (rst_controller_reset_out_reset),                         // main_reset.reset
		.din_data              (alt_vip_cl_csc_0_dout_data),                             //        din.data
		.din_valid             (alt_vip_cl_csc_0_dout_valid),                            //           .valid
		.din_startofpacket     (alt_vip_cl_csc_0_dout_startofpacket),                    //           .startofpacket
		.din_endofpacket       (alt_vip_cl_csc_0_dout_endofpacket),                      //           .endofpacket
		.din_ready             (alt_vip_cl_csc_0_dout_ready),                            //           .ready
		.dout_data             (alt_vip_clip_0_dout_data),                               //       dout.data
		.dout_valid            (alt_vip_clip_0_dout_valid),                              //           .valid
		.dout_startofpacket    (alt_vip_clip_0_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (alt_vip_clip_0_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (alt_vip_clip_0_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_0_alt_vip_clip_0_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_0_alt_vip_clip_0_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_0_alt_vip_clip_0_control_write),         //           .write
		.control_writedata     (mm_interconnect_0_alt_vip_clip_0_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_0_alt_vip_clip_0_control_read),          //           .read
		.control_readdata      (mm_interconnect_0_alt_vip_clip_0_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_0_alt_vip_clip_0_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_alt_vip_clip_0_control_waitrequest)    //           .waitrequest
	);

	DE10_Standard_Qsys_alt_vip_clip_1 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_IN_WIDTH                 (720),
		.MAX_IN_HEIGHT                (576),
		.CLIPPING_METHOD              ("RECTANGLE"),
		.LEFT_OFFSET                  (0),
		.RIGHT_OFFSET                 (10),
		.TOP_OFFSET                   (24),
		.BOTTOM_OFFSET                (10),
		.RECTANGLE_WIDTH              (720),
		.RECTANGLE_HEIGHT             (480),
		.USER_PACKET_SUPPORT          ("PASSTHROUGH"),
		.RUNTIME_CONTROL              (0),
		.LIMITED_READBACK             (0)
	) alt_vip_clip_1 (
		.main_clock         (clk_sys_clk),                         // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_dil_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_dil_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_dil_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_dil_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_dil_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_clip_1_dout_data),            //       dout.data
		.dout_valid         (alt_vip_clip_1_dout_valid),           //           .valid
		.dout_startofpacket (alt_vip_clip_1_dout_startofpacket),   //           .startofpacket
		.dout_endofpacket   (alt_vip_clip_1_dout_endofpacket),     //           .endofpacket
		.dout_ready         (alt_vip_clip_1_dout_ready)            //           .ready
	);

	alt_vipcts131_cts #(
		.BITS_PER_SYMBOL               (8),
		.NUMBER_OF_COLOR_PLANES        (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.TRIGGER_ON_WIDTH_CHANGE       (0),
		.TRIGGER_ON_HEIGHT_CHANGE      (0),
		.TRIGGER_ON_IMAGE_SOP          (1),
		.DISARM_ON_TRIGGER             (1),
		.MAX_INSTRUCTION_COUNT         (10)
	) alt_vip_cts_0 (
		.clock              (clk_sys_clk),                                     //       main_clock.clk
		.reset              (rst_controller_reset_out_reset),                  // main_clock_reset.reset
		.slave_read         (mm_interconnect_0_alt_vip_cts_0_slave_read),      //            slave.read
		.slave_readdata     (mm_interconnect_0_alt_vip_cts_0_slave_readdata),  //                 .readdata
		.slave_write        (mm_interconnect_0_alt_vip_cts_0_slave_write),     //                 .write
		.slave_writedata    (mm_interconnect_0_alt_vip_cts_0_slave_writedata), //                 .writedata
		.slave_address      (mm_interconnect_0_alt_vip_cts_0_slave_address),   //                 .address
		.master_address     (alt_vip_cts_0_master_address),                    //           master.address
		.master_writedata   (alt_vip_cts_0_master_writedata),                  //                 .writedata
		.master_write       (alt_vip_cts_0_master_write),                      //                 .write
		.master_waitrequest (alt_vip_cts_0_master_waitrequest),                //                 .waitrequest
		.status_update_int  (irq_mapper_receiver1_irq),                        // interrupt_sender.irq
		.din_data           (alt_vip_cl_mixer_0_dout_data),                    //              din.data
		.din_valid          (alt_vip_cl_mixer_0_dout_valid),                   //                 .valid
		.din_ready          (alt_vip_cl_mixer_0_dout_ready),                   //                 .ready
		.din_startofpacket  (alt_vip_cl_mixer_0_dout_startofpacket),           //                 .startofpacket
		.din_endofpacket    (alt_vip_cl_mixer_0_dout_endofpacket),             //                 .endofpacket
		.dout_data          (alt_vip_cts_0_dout_data),                         //             dout.data
		.dout_valid         (alt_vip_cts_0_dout_valid),                        //                 .valid
		.dout_ready         (alt_vip_cts_0_dout_ready),                        //                 .ready
		.dout_startofpacket (alt_vip_cts_0_dout_startofpacket),                //                 .startofpacket
		.dout_endofpacket   (alt_vip_cts_0_dout_endofpacket)                   //                 .endofpacket
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (800),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (8000),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (4000),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (30),
		.H_FRONT_PORCH                 (210),
		.H_BACK_PORCH                  (16),
		.V_SYNC_LENGTH                 (13),
		.V_FRONT_PORCH                 (22),
		.V_BACK_PORCH                  (10),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_mtlc (
		.is_clk        (clk_sys_clk),                                  //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),               // is_clk_rst_reset.reset
		.is_data       (alt_vip_cl_clp_1_dout_data),                   //              din.data
		.is_valid      (alt_vip_cl_clp_1_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_cl_clp_1_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_cl_clp_1_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_cl_clp_1_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_itc_mtlc_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_mtlc_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_mtlc_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_mtlc_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_mtlc_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_mtlc_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_mtlc_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_mtlc_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_mtlc_clocked_video_vid_v)          //                 .export
	);

	DE10_Standard_Qsys_alt_vip_scl_0 alt_vip_scl_0 (
		.main_clock            (clk_sys_clk),                                           // main_clock.clk
		.main_reset            (rst_controller_reset_out_reset),                        // main_reset.reset
		.din_data              (alt_vip_clip_0_dout_data),                              //        din.data
		.din_valid             (alt_vip_clip_0_dout_valid),                             //           .valid
		.din_startofpacket     (alt_vip_clip_0_dout_startofpacket),                     //           .startofpacket
		.din_endofpacket       (alt_vip_clip_0_dout_endofpacket),                       //           .endofpacket
		.din_ready             (alt_vip_clip_0_dout_ready),                             //           .ready
		.dout_data             (alt_vip_scl_0_dout_data),                               //       dout.data
		.dout_valid            (alt_vip_scl_0_dout_valid),                              //           .valid
		.dout_startofpacket    (alt_vip_scl_0_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (alt_vip_scl_0_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (alt_vip_scl_0_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_0_alt_vip_scl_0_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_0_alt_vip_scl_0_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_0_alt_vip_scl_0_control_write),         //           .write
		.control_writedata     (mm_interconnect_0_alt_vip_scl_0_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_0_alt_vip_scl_0_control_read),          //           .read
		.control_readdata      (mm_interconnect_0_alt_vip_scl_0_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_0_alt_vip_scl_0_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_alt_vip_scl_0_control_waitrequest)    //           .waitrequest
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (3),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (800),
		.MAX_IMAGE_HEIGHT               (480),
		.MEM_PORT_WIDTH                 (32),
		.RMASTER_FIFO_DEPTH             (1024),
		.RMASTER_BURST_TARGET           (64),
		.CLOCKS_ARE_SEPARATE            (0)
	) alt_vip_vfr_0 (
		.clock                (clk_sys_clk),                                            //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (clk_sys_clk),                                            //            clock_master.clk
		.master_reset         (rst_controller_reset_out_reset),                         //      clock_master_reset.reset
		.slave_address        (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (irq_mapper_receiver0_irq),                               //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	audio_avalon_controller_top audio_avalon_controller (
		.clk                  (clk_clk),                                                    //       clock_reset.clk
		.reset_n              (~rst_controller_001_reset_out_reset),                        // clock_reset_reset.reset_n
		.avs_s1_write_n       (~mm_interconnect_0_audio_avalon_controller_s1_write),        //                s1.write_n
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_controller_s1_writedata),     //                  .writedata
		.avs_s1_read_n        (~mm_interconnect_0_audio_avalon_controller_s1_read),         //                  .read_n
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_controller_s1_readdata),      //                  .readdata
		.avs_s1_begintransfer (mm_interconnect_0_audio_avalon_controller_s1_begintransfer), //                  .begintransfer
		.avs_s1_addr          (mm_interconnect_0_audio_avalon_controller_s1_address),       //                  .address
		.avs_s1_cs_n          (~mm_interconnect_0_audio_avalon_controller_s1_chipselect),   //                  .chipselect_n
		.avs_s1_readyfordata  (),                                                           //                  .readyfordata
		.avs_s1_dataavailable (),                                                           //                  .dataavailable
		.avs_s1_irq           (irq_synchronizer_002_receiver_irq),                          //            irq_s1.irq
		.audio_CLK            (audio_avalon_controller_conduit_end_CLK),                    //       conduit_end.export
		.audio_LRCIN          (audio_avalon_controller_conduit_end_LRCIN),                  //                  .export
		.audio_DIN            (audio_avalon_controller_conduit_end_DIN),                    //                  .export
		.audio_LRCOUT         (audio_avalon_controller_conduit_end_LRCOUT),                 //                  .export
		.audio_DOUT           (audio_avalon_controller_conduit_end_DOUT),                   //                  .export
		.audio_BCLK           (audio_avalon_controller_conduit_end_BCLK)                    //                  .export
	);

	DE10_Standard_Qsys_av_i2c_clk_pio av_i2c_clk_pio (
		.clk        (clk_sys_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_av_i2c_clk_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_av_i2c_clk_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_av_i2c_clk_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_av_i2c_clk_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_av_i2c_clk_pio_s1_readdata),   //                    .readdata
		.out_port   (av_i2c_clk_pio_external_connection_export)       // external_connection.export
	);

	DE10_Standard_Qsys_av_i2c_data_pio av_i2c_data_pio (
		.clk        (clk_sys_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_av_i2c_data_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_av_i2c_data_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_av_i2c_data_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_av_i2c_data_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_av_i2c_data_pio_s1_readdata),   //                    .readdata
		.bidir_port (av_i2c_data_pio_external_connection_export)       // external_connection.export
	);

	DE10_Standard_Qsys_button_pio button_pio (
		.clk        (clk_sys_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                    //                 irq.irq
	);

	DE10_Standard_Qsys_jtag_uart jtag_uart (
		.clk            (clk_sys_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                   //               irq.irq
	);

	DE10_Standard_Qsys_led_pio led_pio (
		.clk        (clk_sys_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)       // external_connection.export
	);

	DE10_Standard_Qsys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_sys_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	DE10_Standard_Qsys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_sys_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	DE10_Standard_Qsys_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (clk_sdram_clk),       // outclk0.clk
		.outclk_1 (clk_sys_clk),         // outclk1.clk
		.outclk_2 (clk_mtlc_clk),        // outclk2.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	DE10_Standard_Qsys_sdram sdram (
		.clk            (clk_sys_clk),                              //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	DE10_Standard_Qsys_sys_clk_timer sys_clk_timer (
		.clk        (clk_sys_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                       //   irq.irq
	);

	DE10_Standard_Qsys_sysid sysid (
		.clock    (clk_sys_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	DE10_Standard_Qsys_av_i2c_clk_pio td_reset_pio (
		.clk        (clk_sys_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_td_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_td_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_td_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_td_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_td_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (td_reset_pio_external_connection_export)       // external_connection.export
	);

	i2c_opencores touch_i2c_opencores (
		.wb_clk_i   (clk_clk),                                                          //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (touch_i2c_opencores_export_scl_pad_io),                            //           export.export
		.sda_pad_io (touch_i2c_opencores_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_receiver_irq)                                     // interrupt_sender.irq
	);

	DE10_Standard_Qsys_touch_int_n touch_int_n (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_touch_int_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_int_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_int_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_int_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_int_n_s1_readdata),   //                    .readdata
		.in_port    (touch_int_n_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)            //                 irq.irq
	);

	DE10_Standard_Qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                               (clk_clk),                                                           //                                             clk_50_clk.clk
		.pll_0_outclk1_clk                                            (clk_sys_clk),                                                       //                                          pll_0_outclk1.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                    // alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.touch_i2c_opencores_clock_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                                //  touch_i2c_opencores_clock_reset_reset_bridge_in_reset.reset
		.alt_vip_cl_vfb_0_mem_master_rd_address                       (alt_vip_cl_vfb_0_mem_master_rd_address),                            //                         alt_vip_cl_vfb_0_mem_master_rd.address
		.alt_vip_cl_vfb_0_mem_master_rd_waitrequest                   (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),                        //                                                       .waitrequest
		.alt_vip_cl_vfb_0_mem_master_rd_burstcount                    (alt_vip_cl_vfb_0_mem_master_rd_burstcount),                         //                                                       .burstcount
		.alt_vip_cl_vfb_0_mem_master_rd_read                          (alt_vip_cl_vfb_0_mem_master_rd_read),                               //                                                       .read
		.alt_vip_cl_vfb_0_mem_master_rd_readdata                      (alt_vip_cl_vfb_0_mem_master_rd_readdata),                           //                                                       .readdata
		.alt_vip_cl_vfb_0_mem_master_rd_readdatavalid                 (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid),                      //                                                       .readdatavalid
		.alt_vip_cl_vfb_0_mem_master_wr_address                       (alt_vip_cl_vfb_0_mem_master_wr_address),                            //                         alt_vip_cl_vfb_0_mem_master_wr.address
		.alt_vip_cl_vfb_0_mem_master_wr_waitrequest                   (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),                        //                                                       .waitrequest
		.alt_vip_cl_vfb_0_mem_master_wr_burstcount                    (alt_vip_cl_vfb_0_mem_master_wr_burstcount),                         //                                                       .burstcount
		.alt_vip_cl_vfb_0_mem_master_wr_byteenable                    (alt_vip_cl_vfb_0_mem_master_wr_byteenable),                         //                                                       .byteenable
		.alt_vip_cl_vfb_0_mem_master_wr_write                         (alt_vip_cl_vfb_0_mem_master_wr_write),                              //                                                       .write
		.alt_vip_cl_vfb_0_mem_master_wr_writedata                     (alt_vip_cl_vfb_0_mem_master_wr_writedata),                          //                                                       .writedata
		.alt_vip_cts_0_master_address                                 (alt_vip_cts_0_master_address),                                      //                                   alt_vip_cts_0_master.address
		.alt_vip_cts_0_master_waitrequest                             (alt_vip_cts_0_master_waitrequest),                                  //                                                       .waitrequest
		.alt_vip_cts_0_master_write                                   (alt_vip_cts_0_master_write),                                        //                                                       .write
		.alt_vip_cts_0_master_writedata                               (alt_vip_cts_0_master_writedata),                                    //                                                       .writedata
		.alt_vip_vfr_0_avalon_master_address                          (alt_vip_vfr_0_avalon_master_address),                               //                            alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                      (alt_vip_vfr_0_avalon_master_waitrequest),                           //                                                       .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                       (alt_vip_vfr_0_avalon_master_burstcount),                            //                                                       .burstcount
		.alt_vip_vfr_0_avalon_master_read                             (alt_vip_vfr_0_avalon_master_read),                                  //                                                       .read
		.alt_vip_vfr_0_avalon_master_readdata                         (alt_vip_vfr_0_avalon_master_readdata),                              //                                                       .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                    (alt_vip_vfr_0_avalon_master_readdatavalid),                         //                                                       .readdatavalid
		.nios2_gen2_0_data_master_address                             (nios2_gen2_0_data_master_address),                                  //                               nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                         (nios2_gen2_0_data_master_waitrequest),                              //                                                       .waitrequest
		.nios2_gen2_0_data_master_byteenable                          (nios2_gen2_0_data_master_byteenable),                               //                                                       .byteenable
		.nios2_gen2_0_data_master_read                                (nios2_gen2_0_data_master_read),                                     //                                                       .read
		.nios2_gen2_0_data_master_readdata                            (nios2_gen2_0_data_master_readdata),                                 //                                                       .readdata
		.nios2_gen2_0_data_master_write                               (nios2_gen2_0_data_master_write),                                    //                                                       .write
		.nios2_gen2_0_data_master_writedata                           (nios2_gen2_0_data_master_writedata),                                //                                                       .writedata
		.nios2_gen2_0_data_master_debugaccess                         (nios2_gen2_0_data_master_debugaccess),                              //                                                       .debugaccess
		.nios2_gen2_0_instruction_master_address                      (nios2_gen2_0_instruction_master_address),                           //                        nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                  (nios2_gen2_0_instruction_master_waitrequest),                       //                                                       .waitrequest
		.nios2_gen2_0_instruction_master_read                         (nios2_gen2_0_instruction_master_read),                              //                                                       .read
		.nios2_gen2_0_instruction_master_readdata                     (nios2_gen2_0_instruction_master_readdata),                          //                                                       .readdata
		.nios2_gen2_0_instruction_master_readdatavalid                (nios2_gen2_0_instruction_master_readdatavalid),                     //                                                       .readdatavalid
		.alt_vip_cl_mixer_0_control_address                           (mm_interconnect_0_alt_vip_cl_mixer_0_control_address),              //                             alt_vip_cl_mixer_0_control.address
		.alt_vip_cl_mixer_0_control_write                             (mm_interconnect_0_alt_vip_cl_mixer_0_control_write),                //                                                       .write
		.alt_vip_cl_mixer_0_control_read                              (mm_interconnect_0_alt_vip_cl_mixer_0_control_read),                 //                                                       .read
		.alt_vip_cl_mixer_0_control_readdata                          (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdata),             //                                                       .readdata
		.alt_vip_cl_mixer_0_control_writedata                         (mm_interconnect_0_alt_vip_cl_mixer_0_control_writedata),            //                                                       .writedata
		.alt_vip_cl_mixer_0_control_byteenable                        (mm_interconnect_0_alt_vip_cl_mixer_0_control_byteenable),           //                                                       .byteenable
		.alt_vip_cl_mixer_0_control_readdatavalid                     (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdatavalid),        //                                                       .readdatavalid
		.alt_vip_cl_mixer_0_control_waitrequest                       (mm_interconnect_0_alt_vip_cl_mixer_0_control_waitrequest),          //                                                       .waitrequest
		.alt_vip_clip_0_control_address                               (mm_interconnect_0_alt_vip_clip_0_control_address),                  //                                 alt_vip_clip_0_control.address
		.alt_vip_clip_0_control_write                                 (mm_interconnect_0_alt_vip_clip_0_control_write),                    //                                                       .write
		.alt_vip_clip_0_control_read                                  (mm_interconnect_0_alt_vip_clip_0_control_read),                     //                                                       .read
		.alt_vip_clip_0_control_readdata                              (mm_interconnect_0_alt_vip_clip_0_control_readdata),                 //                                                       .readdata
		.alt_vip_clip_0_control_writedata                             (mm_interconnect_0_alt_vip_clip_0_control_writedata),                //                                                       .writedata
		.alt_vip_clip_0_control_byteenable                            (mm_interconnect_0_alt_vip_clip_0_control_byteenable),               //                                                       .byteenable
		.alt_vip_clip_0_control_readdatavalid                         (mm_interconnect_0_alt_vip_clip_0_control_readdatavalid),            //                                                       .readdatavalid
		.alt_vip_clip_0_control_waitrequest                           (mm_interconnect_0_alt_vip_clip_0_control_waitrequest),              //                                                       .waitrequest
		.alt_vip_cts_0_slave_address                                  (mm_interconnect_0_alt_vip_cts_0_slave_address),                     //                                    alt_vip_cts_0_slave.address
		.alt_vip_cts_0_slave_write                                    (mm_interconnect_0_alt_vip_cts_0_slave_write),                       //                                                       .write
		.alt_vip_cts_0_slave_read                                     (mm_interconnect_0_alt_vip_cts_0_slave_read),                        //                                                       .read
		.alt_vip_cts_0_slave_readdata                                 (mm_interconnect_0_alt_vip_cts_0_slave_readdata),                    //                                                       .readdata
		.alt_vip_cts_0_slave_writedata                                (mm_interconnect_0_alt_vip_cts_0_slave_writedata),                   //                                                       .writedata
		.alt_vip_scl_0_control_address                                (mm_interconnect_0_alt_vip_scl_0_control_address),                   //                                  alt_vip_scl_0_control.address
		.alt_vip_scl_0_control_write                                  (mm_interconnect_0_alt_vip_scl_0_control_write),                     //                                                       .write
		.alt_vip_scl_0_control_read                                   (mm_interconnect_0_alt_vip_scl_0_control_read),                      //                                                       .read
		.alt_vip_scl_0_control_readdata                               (mm_interconnect_0_alt_vip_scl_0_control_readdata),                  //                                                       .readdata
		.alt_vip_scl_0_control_writedata                              (mm_interconnect_0_alt_vip_scl_0_control_writedata),                 //                                                       .writedata
		.alt_vip_scl_0_control_byteenable                             (mm_interconnect_0_alt_vip_scl_0_control_byteenable),                //                                                       .byteenable
		.alt_vip_scl_0_control_readdatavalid                          (mm_interconnect_0_alt_vip_scl_0_control_readdatavalid),             //                                                       .readdatavalid
		.alt_vip_scl_0_control_waitrequest                            (mm_interconnect_0_alt_vip_scl_0_control_waitrequest),               //                                                       .waitrequest
		.alt_vip_vfr_0_avalon_slave_address                           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),              //                             alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                             (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),                //                                                       .write
		.alt_vip_vfr_0_avalon_slave_read                              (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),                 //                                                       .read
		.alt_vip_vfr_0_avalon_slave_readdata                          (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),             //                                                       .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                         (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata),            //                                                       .writedata
		.audio_avalon_controller_s1_address                           (mm_interconnect_0_audio_avalon_controller_s1_address),              //                             audio_avalon_controller_s1.address
		.audio_avalon_controller_s1_write                             (mm_interconnect_0_audio_avalon_controller_s1_write),                //                                                       .write
		.audio_avalon_controller_s1_read                              (mm_interconnect_0_audio_avalon_controller_s1_read),                 //                                                       .read
		.audio_avalon_controller_s1_readdata                          (mm_interconnect_0_audio_avalon_controller_s1_readdata),             //                                                       .readdata
		.audio_avalon_controller_s1_writedata                         (mm_interconnect_0_audio_avalon_controller_s1_writedata),            //                                                       .writedata
		.audio_avalon_controller_s1_begintransfer                     (mm_interconnect_0_audio_avalon_controller_s1_begintransfer),        //                                                       .begintransfer
		.audio_avalon_controller_s1_chipselect                        (mm_interconnect_0_audio_avalon_controller_s1_chipselect),           //                                                       .chipselect
		.av_i2c_clk_pio_s1_address                                    (mm_interconnect_0_av_i2c_clk_pio_s1_address),                       //                                      av_i2c_clk_pio_s1.address
		.av_i2c_clk_pio_s1_write                                      (mm_interconnect_0_av_i2c_clk_pio_s1_write),                         //                                                       .write
		.av_i2c_clk_pio_s1_readdata                                   (mm_interconnect_0_av_i2c_clk_pio_s1_readdata),                      //                                                       .readdata
		.av_i2c_clk_pio_s1_writedata                                  (mm_interconnect_0_av_i2c_clk_pio_s1_writedata),                     //                                                       .writedata
		.av_i2c_clk_pio_s1_chipselect                                 (mm_interconnect_0_av_i2c_clk_pio_s1_chipselect),                    //                                                       .chipselect
		.av_i2c_data_pio_s1_address                                   (mm_interconnect_0_av_i2c_data_pio_s1_address),                      //                                     av_i2c_data_pio_s1.address
		.av_i2c_data_pio_s1_write                                     (mm_interconnect_0_av_i2c_data_pio_s1_write),                        //                                                       .write
		.av_i2c_data_pio_s1_readdata                                  (mm_interconnect_0_av_i2c_data_pio_s1_readdata),                     //                                                       .readdata
		.av_i2c_data_pio_s1_writedata                                 (mm_interconnect_0_av_i2c_data_pio_s1_writedata),                    //                                                       .writedata
		.av_i2c_data_pio_s1_chipselect                                (mm_interconnect_0_av_i2c_data_pio_s1_chipselect),                   //                                                       .chipselect
		.button_pio_s1_address                                        (mm_interconnect_0_button_pio_s1_address),                           //                                          button_pio_s1.address
		.button_pio_s1_write                                          (mm_interconnect_0_button_pio_s1_write),                             //                                                       .write
		.button_pio_s1_readdata                                       (mm_interconnect_0_button_pio_s1_readdata),                          //                                                       .readdata
		.button_pio_s1_writedata                                      (mm_interconnect_0_button_pio_s1_writedata),                         //                                                       .writedata
		.button_pio_s1_chipselect                                     (mm_interconnect_0_button_pio_s1_chipselect),                        //                                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),             //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),               //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),            //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),           //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),         //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),          //                                                       .chipselect
		.led_pio_s1_address                                           (mm_interconnect_0_led_pio_s1_address),                              //                                             led_pio_s1.address
		.led_pio_s1_write                                             (mm_interconnect_0_led_pio_s1_write),                                //                                                       .write
		.led_pio_s1_readdata                                          (mm_interconnect_0_led_pio_s1_readdata),                             //                                                       .readdata
		.led_pio_s1_writedata                                         (mm_interconnect_0_led_pio_s1_writedata),                            //                                                       .writedata
		.led_pio_s1_chipselect                                        (mm_interconnect_0_led_pio_s1_chipselect),                           //                                                       .chipselect
		.nios2_gen2_0_debug_mem_slave_address                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),            //                           nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),              //                                                       .write
		.nios2_gen2_0_debug_mem_slave_read                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),               //                                                       .read
		.nios2_gen2_0_debug_mem_slave_readdata                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),           //                                                       .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),          //                                                       .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),         //                                                       .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),        //                                                       .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),        //                                                       .debugaccess
		.onchip_memory2_0_s1_address                                  (mm_interconnect_0_onchip_memory2_0_s1_address),                     //                                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                    (mm_interconnect_0_onchip_memory2_0_s1_write),                       //                                                       .write
		.onchip_memory2_0_s1_readdata                                 (mm_interconnect_0_onchip_memory2_0_s1_readdata),                    //                                                       .readdata
		.onchip_memory2_0_s1_writedata                                (mm_interconnect_0_onchip_memory2_0_s1_writedata),                   //                                                       .writedata
		.onchip_memory2_0_s1_byteenable                               (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                  //                                                       .byteenable
		.onchip_memory2_0_s1_chipselect                               (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                  //                                                       .chipselect
		.onchip_memory2_0_s1_clken                                    (mm_interconnect_0_onchip_memory2_0_s1_clken),                       //                                                       .clken
		.sdram_s1_address                                             (mm_interconnect_0_sdram_s1_address),                                //                                               sdram_s1.address
		.sdram_s1_write                                               (mm_interconnect_0_sdram_s1_write),                                  //                                                       .write
		.sdram_s1_read                                                (mm_interconnect_0_sdram_s1_read),                                   //                                                       .read
		.sdram_s1_readdata                                            (mm_interconnect_0_sdram_s1_readdata),                               //                                                       .readdata
		.sdram_s1_writedata                                           (mm_interconnect_0_sdram_s1_writedata),                              //                                                       .writedata
		.sdram_s1_byteenable                                          (mm_interconnect_0_sdram_s1_byteenable),                             //                                                       .byteenable
		.sdram_s1_readdatavalid                                       (mm_interconnect_0_sdram_s1_readdatavalid),                          //                                                       .readdatavalid
		.sdram_s1_waitrequest                                         (mm_interconnect_0_sdram_s1_waitrequest),                            //                                                       .waitrequest
		.sdram_s1_chipselect                                          (mm_interconnect_0_sdram_s1_chipselect),                             //                                                       .chipselect
		.sys_clk_timer_s1_address                                     (mm_interconnect_0_sys_clk_timer_s1_address),                        //                                       sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                                       (mm_interconnect_0_sys_clk_timer_s1_write),                          //                                                       .write
		.sys_clk_timer_s1_readdata                                    (mm_interconnect_0_sys_clk_timer_s1_readdata),                       //                                                       .readdata
		.sys_clk_timer_s1_writedata                                   (mm_interconnect_0_sys_clk_timer_s1_writedata),                      //                                                       .writedata
		.sys_clk_timer_s1_chipselect                                  (mm_interconnect_0_sys_clk_timer_s1_chipselect),                     //                                                       .chipselect
		.sysid_control_slave_address                                  (mm_interconnect_0_sysid_control_slave_address),                     //                                    sysid_control_slave.address
		.sysid_control_slave_readdata                                 (mm_interconnect_0_sysid_control_slave_readdata),                    //                                                       .readdata
		.td_reset_pio_s1_address                                      (mm_interconnect_0_td_reset_pio_s1_address),                         //                                        td_reset_pio_s1.address
		.td_reset_pio_s1_write                                        (mm_interconnect_0_td_reset_pio_s1_write),                           //                                                       .write
		.td_reset_pio_s1_readdata                                     (mm_interconnect_0_td_reset_pio_s1_readdata),                        //                                                       .readdata
		.td_reset_pio_s1_writedata                                    (mm_interconnect_0_td_reset_pio_s1_writedata),                       //                                                       .writedata
		.td_reset_pio_s1_chipselect                                   (mm_interconnect_0_td_reset_pio_s1_chipselect),                      //                                                       .chipselect
		.touch_i2c_opencores_avalon_slave_0_address                   (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_address),      //                     touch_i2c_opencores_avalon_slave_0.address
		.touch_i2c_opencores_avalon_slave_0_write                     (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_write),        //                                                       .write
		.touch_i2c_opencores_avalon_slave_0_readdata                  (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_readdata),     //                                                       .readdata
		.touch_i2c_opencores_avalon_slave_0_writedata                 (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_writedata),    //                                                       .writedata
		.touch_i2c_opencores_avalon_slave_0_waitrequest               (~mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_waitrequest), //                                                       .waitrequest
		.touch_i2c_opencores_avalon_slave_0_chipselect                (mm_interconnect_0_touch_i2c_opencores_avalon_slave_0_chipselect),   //                                                       .chipselect
		.touch_int_n_s1_address                                       (mm_interconnect_0_touch_int_n_s1_address),                          //                                         touch_int_n_s1.address
		.touch_int_n_s1_write                                         (mm_interconnect_0_touch_int_n_s1_write),                            //                                                       .write
		.touch_int_n_s1_readdata                                      (mm_interconnect_0_touch_int_n_s1_readdata),                         //                                                       .readdata
		.touch_int_n_s1_writedata                                     (mm_interconnect_0_touch_int_n_s1_writedata),                        //                                                       .writedata
		.touch_int_n_s1_chipselect                                    (mm_interconnect_0_touch_int_n_s1_chipselect)                        //                                                       .chipselect
	);

	DE10_Standard_Qsys_irq_mapper irq_mapper (
		.clk           (clk_sys_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (clk_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (clk_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (clk_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_sys_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
