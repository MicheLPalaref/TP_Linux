��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U������Qܻ�#VQ�ٍ�BQm<CA��}q��Э�d����i�����U$^�\��o!�gu�Db#��e���)�؍�IAV��:��G��&B&{n�C��bBR�E���|��E3_}׳�`w���w��1US���Z�X6�����\�S���:����s;x,շ�v)a��!��l�X��3��K7��I������O�1@F�R��ܥ�[�/���1����_h��	�����8,B�6�q�9���W���������	��Z��'9]/͔�Nꓹ���b���O��q@�hDp�:� }fCQ� ͗A�4�ۿ���>)hB�osɑO_sˬ�0���Z�2�ye�㭗��	�4���?�74�y��A����l��O'�9I܉�h��O�sZ����ck?���]5o��ç������+��G	!r�X�3g��pK�W9�m.���� ��'�<�G �;)���6�_ŏ6@6(�3���2�j��֮�������K��p��o �܆P�����9�О�#�ϸ��]���'̒�C����ΟT7��߲� �#J]2܉����;�r��z�d�Y�*dG��K��Ӝ��+oWÂ�t�F¬�ћB�����-.�M���vف� �R2���_T�|��S�T5��7��L�(��X@�݌��-j� F��K �%���.�)Zt~�8�ތ���J�ێ�;��Ȥ�[��s�c(K2m�;�v�&B��J�'惜֓ks�2���:IL��B�4���qvW�� �LPDt�f�KQ8E�9~��A�[TPg\_۸c�y)\��|�J	l�+a�X�P?�����D������(�:֒�M�����ǒ�����b0�0����s{�GZk��%�{�s;;���"y��r��}�oWz��Q�����?�W�����޻�����B����K�UB2�1�����X�?,j"�H9�Iy�*&�����q���od9��*@ȯ���|]�\�ܞ�jk�