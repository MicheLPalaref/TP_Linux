��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����`��B�㓪F:��ew���@�C�k�.U6�vά1�xrl9��Sr?$R�t��M��~3pwd��<�i��w_�)4ޟo$#)����4F�1s[�p;��Q�!q��i�u�k�
rw���b�Q�G�Et���M��%�b�1��L����%Y�{pI �sW=��߁ޏt��`��/�M!���=Y;t�~����4���S_��2�NQ}]W`o��ϽL�{׸;��'9<�!�	��p���[3��J�?d���Z�׶��v�GT�H<5Y�Ցu�Xc[�1^�#�7��eq���=sY�W������Y��y��@62�E�{G��к�3B�UZ	qnI<#{�w[U���(#Jk���qϽit[��^�"OE��0&&�'k���VQܢKr�<%�����)D���LnE&�g���iR�I�.��0��C�WQ)���K�:�͊�q�X�J�=X� �^�B=^�'i���b͸���-�q�{�����ω���.��;c�$FS�?d?�DR8�
i�+1(t6���%��7���b�-/�� D.��<��!�h��AB
^��1��hO/��l����V�B��"����N��3��!�%y{�	��1x�Х���w1NL<�Е0,�(�plL�v�vp��K����f�)�����A�����d���U���C;1��g�Q>x�*�������������@�{vO)�H>;���a������Ajgw�m(L56&>9�
I����z�i�������Q/����1��3T�BO�.%��
�C(+��J�R�s��ݾ$)#y��,,8�$pS�v�R�s!��۹ђUݟ-���S	�H'�ia|E���>X<�7��Zy֥��Ȱ5\��C��*>$X�D��	kG���>�4� �Ut��b�>�Ą�X?byƔ���On�ޜ^�j���ZBǵs��{��4/�л����:�����>��R/lNN��-OzX}��]����`eZ��mh��S=�7^���P�I3����6:�
��O�pO#�������\t킄;ۭ��	�+ZE>>��Aww������jp���\�5�۱>�Z�8�^۷������Qs**Ep�_���V��ϕ8y�b�
�� 5dU��w�T�Z�?��I��m�u�g ��Aj&:9!5L��4���yQƅM�z�����aˈ	�:�x�YZC\T�q��]Cod(U�K��>�4�s�M|@c�w�>��n�[!h��lO�%ގ����-�_�(���Ӗ�� ��jB[zh�g.`ԙ�9��ɛ����-@3S��ԵX�b�U]=B�4�Ӽ�E�c�,*�!���})>E��Л�!����L&�M]���l�d{ �_жs�̞��1c;h��G)2��v��#�*88�ĝ#�4J���z;|~��}�f����/6`O�Zd�N{�P8����e�ݟ��x���,���o��c�HP?&p�B����831���/a/�E�!qV�֍k�	�V0`៵A�D��7�&��E��bQ�_:�)�cq�6������&�7�e2��E������4�q�`%��zƯ�z}��>�����wZ6�ABۮ�?.g}��f� gg�pM�d��p!�C"�H2Li���h3_{�v4��a�u�=�W<g��(Y���V0{>Os�D=�M�ߔ��Rklu�&�f$�IC@LW/ْ�2�����R�I���T�x�&]}i�ڏ��U���R��L�[G^�џ���,�
�{� `�Wz�ĉ9d=O���:"��cʩS;dc%���=�~`��#=��/W��s隋e(n	���Z��>�l��ry���~]?@��}�%�dR�
�[�D�[O�w����� �brڹɳ��1������ ���BX�qGy��-kz�t�$[z�^9&��]ހS��}�[���,���m�*�c�B@�2E��ɛ9d5�yf�r�0?��4�pb����N����=CjY�=+��g�|�kA�3#�
L� i���pБ�1�)p���(�"W�����i�t����ˈ�L�sn��n'�_
W�1�t�u!��1���ֆ3��u�Д��"�V�yc���2�A����s�,� ��ge|}�ţ�RR��R�(dVM���U�w���S�q,im��b�̤N��!-�ܗb���&��c�v��zU�X�n^[s��Z��|\^$i��6=l�JB҉^)���NY�D���r�~ެ�(h�?���� ���_�C�*�}�6���;dI�8 R��$E�{۲��H�o\�"�,	���kz��u�{����G�f� ۗ�s��Y$�|���ʢȳ���O��i�O�7g_��
���2m͜��W�N��y�W��'�T�f~V;�,�{��k'�Kj���k\���*�:��BQJ�r�O�e��@�����M��5���xs�I���W/�q9�/
0B�[�~]���L��#�-��&�Qt��j(PkntbQ�_�c���듘������ȱ����Dj$��:;v�N�2_S[R���"(#+���V�'Zj��o �V�}k��;��أ^r����i>�mA9(�_lX��o���1�C�w?���pƥ����>|Wh;�*]���W�Y�{��.@�1���d6����EV�v�{�����SI��X��@�-���t��j��p���Ʈ��hC^�$<���Kϵ��7��Ґ7q����������{��3�&&r�̩S4����?&&�xuZ?�zۖ����Y��l���������',+CL4��w�g+Uܖf`�)y��	`�e؟v���^#ɜ7�tsg6H��y��C�^���G�F�Mנ�)�^'�i��(��i$�Τ�;�p��8q�3�ݬ�&�� /�&}�ZU�C���{�Y=Ч|�<�7㶈��.�{�d	3nI�/�f�74�A�T�uw~WM\�u��#\ɚ�h�8���7&�����Q���'O/��Z��=��G�x�'�)yC�_�$��rS�^X�D�f2���D�q[���<�e-ϑko݊�`�qŔL��ܞ��^��C@�ՙ��}Ot-���IΙ�u�,���z��g�0W���A��~,z��{��eA0��6��B�j>��B�!
�|O˰���ԩk=4�ݲ_P��tګ��wN��3�I*4T�
�$�?t'��N<Bc��^XX�ٗ�E���3�{�Ò�Z\��{B�H�0������z�G���E����a0���(�9�Y�d���Z+�$iHe-_81Ս�AdL��8�bщX�����q�}:6�óڭ��B�E�:폀�ٛTQ���P��nh�����~A�LU��RQj��F��v3!� �Xr5%[���,~!H�Ψ�/�
�1�7�ks�,�w��W�9�Hn�	�9QDA.O(
�V�]FM�ܣ��ME��]u)�N�i����{S�q��=O���KГU�8���U�}V�}��9�~Tg�0B|�;0�������Wb�>՛s�篝C@V�y~n�Z�Vgq���ӌg�����/���-Q4�Z*Wſ��PS��3��.�0b�8	5*��)D�ѩ�]�4���ưt�P���V�"�"�2�Ig�d��K��Ƃ����f�mM���ȅ��^����l�U�EhO�-�D�糞q��UhLH�-�VmX@m YP$K4�[�d��E}�kP�2z#�5N���1�&,��t��{���<J�R�$�ψ��U<��x�֫E>\����Ǵ�ٺ(��RԘ��aQ�ݟO��"��-�T�~���r�kx�=[�>A┦�@� y�;Ɯ^
o��U.��/	/ش���[����|*�I�m�E3�(�~���<��{����c:���J���?��+�#͂!M����jP�
�����?�.Ї��9�{:�|&���W�C%;�׆�I��]!b|*^\X�������L�Sw��f�v�3}Q�5^�����A�a��[<�h�)`��Cp��u�y@W0����)l����G��. �!� �Xgڝ�4�h(�A�h*�`l�$��4sO��Y�7�δJ�h8��d�}���j� �tX4��Ȳ��@q���''o���6�4W�q��w_֨ ۨ��t�y%�Bd]$]m�Dd�~�j$��0�t��а���4+5�����_����!㾅$���H��]���F_�)��Y2��)�E_kh��%%^[�-�g23�[��¨�+�lJ����&�!���2C1��np!���b:[�eU�;��Ƹ��x�
yM���:���&6�9 X*9M���gx=�0@�}��pe
�qo�
|�戳=�x��p��ڤ~�?@�ḳ�fê��(���'!l{<�3fK��Gr�����=�!d);����ߛ��|0�}(/4��G��&]�-꽒�)�9誽��.�8?�}F��Cp��2UND&��pU�� R�=��!ə��M��i�E��ɏd�v	]��]��z� ��-�w1(��z�S���?�Ag�B��hVbY,]}ƻJ{��Z�g��*3�*RD�J����f�}�/"�d6�v0}Q����@�Fi�[����||J>��F��A���,ǚFD�[�n51��sRa-���;+��X.}u��2!�,r#g����&e�\SvJ&������AC��*i
��Pz�}�^�:��a�Qs�ū����j
��=F���͍�����ͳ�������@�� .���Y�/f|�At\��h�E&:����0@j�W�Z�P���IG*=J�GW�m�-{.fhY�.Qw,0�'	4���1�N�:Wgmw��K_9.~���c�_�kS)i�P�I��.�'_�Ǒ�B�t�Nrc�" =p4S�8��T2�af4[��@I�w�Z�d�K�o�������ŃJ\РڙG��L�l�	�����x*	��|�R�ͩ����-��;*8���a������T�_���N�+B�i��[	='�Dȭ�|S~�bʳM�"�X�����`�������e�ɥY�v�J6Ӣ͖��T�����q�9�_DY4ʶ�b���]���v����f�55Z�n�0i��y�6��p��p�wZX��~;�;���z����l�F�R8=�>�X��e�yv�5��J%o�6uKؠ�(yo�A Wo[���J0`%�L�� a���`�Q�MGj��\�M���+�l�<~!�%�W,u��.Q��6������I��P|�tX*7��,����ij~d�O�!7DI�a�AI����3Y��P����s���
*7$�"|~l�DK���h���Rf?��(��!Ȼ��oiΝb��ඒ��U�cq�0a�? �a���K��g�f_SU�2��+�j���P�E����X>�!z:h����������&+�8|�8G"��%Gp�W�WDrkJ=Ѓ����;��I?�U�i�����E~T�+/a��.�&�o]k}�~r����V|]�r�.�l|3l;���l��P�Z��ւۘqT����Ș�2%�+�8�}Y��!�῀���l��#�c�a��kô �Iz�� �=X,��S���a��GtY�f�<v�|�;�v"�����<!��;��2�/|�J0x�?����_1�]�����
�͢���P&�c�h��
��5��l�`ǬC&;�Lh~?@���9ot��z�a�#<��m��E2`5ri�/��+���+P���6��O�9g��9��\Q�j�gV�0�Ԯy4�H�zHX�r��<_�?%�.�U+ ��u�rS���p?�A@�-N_䶋SdU��oWgg�9�ԏFh�`w0�2-Y�3X�E`���7\�GcL:�B��SH� a�/���@rJ{n �K�n�������F`��Z�u><�dhFO)Z�;�ʼM�ϣ]�*ͣ�o�ebs��x��/c�yP� QF�!}�ҥ�ħN	�W��hj{+���DI������~��őx��
��#�����p9��+T8�d�O2�������K�bi����W�x%Q��T�-J������} ����b?/�w��n�+���-
�+�����2���<S~9��a�|�2{�~�����_*�X�o� �{�'�n��%�J���iR����Kӿ�y63S�����rx���J0ܼ7�1Ì"�ղ>����L�I>ʌм�{��'E�=y����VS�R�=0��[2�D�t�'J�7�mc���@�ׯn�:62h���Q�C!1,1z�
��/)	"��G�wS��3�p�9�B���qV~�;H�F�}�GH�Du��z`�z�~�]LD�Y��3
5���4��X򚈡m3{}��R2��1e;��A)�]nQz�q�D���?%}��UQ�G��F(ձg�ɾ��6S����>#�n�%W̺x�6D�����ӆK��8S�7ͺ�w�IƘcNУxT�`��j��/�{K�»�c�1����v���vT+� ݻ}�{&ۚV���twT�`�a��4[�b��O�D�䎑�-C"�����n�;� Ƨ�oPM?�8g��9O���Vd��X{���s��ؒH+���9�l:�m�K�a�=I���*;Tfabc����	r|�<�����%�!�r��x�(���a	c��������O�؆N�i@�O�񧦨�ǲFrn��^�~���{J�D�cR/�50�ܖ�H-�ӯM���=��5�ز��k�z9��9�z�M��TÍ�/P��^�[I#g���C�	�e�1�(�S��&�)�[n��7�� �4�w��')�ۡ!�&�=NV��5E�L��K��J�V�~< ���S����+��7�@�"�>�;r:���?Yr�`�#����Z�
j��K�A��gw.�9=�˭*��깳�����j�/���Y�!e����eyLj��u L����v�����!֊��Oi�]���ƕcㆥR�4�p�Ua�	hm�s.-B'�����6�c ��!���+�!zY�/�B���s�4�้��7{2ws63�osaK��|	`�/s1��J9��*!\�(��kR�˫{�5ts.�ί5Z�Q�\j�[ͳ�b�u���U7�+�^���s�1N� |��Fø����r"����B8 �%� �,㋙����%�V��|����$v�Ji/���NzF�2v�e��O-��C߈��%�����C���"A��Ye�am�(�b�F%\��Ǖ`J4�s���_j4�m�J}�!x�����]���5����I�}JA�uF~
x�r]6�\}�JVw͟�裎ñg��1�-����#+��^�3o����86��@|�M��9e���t"�! �����L�C�WH�SG�= �P���/�ZA�kU�t�3�Zk�|"*���`�9q
(HL��x�Mɭ���GB�g�u00�sb�ՄOx�ىj���Ƚ05�n�Ŵ������N�}ޮ�ҲLt�#'�3�+
%=t�?B�j�-�!1�tTi�3#V
^ X�j�wC&�'|�ڐ���ݘd�dX�'�!.2cU���; R��B���g��$N*Ȁ�ްuƷ���vA,�F{�P�k�E���(j}�K�JLK1Q6�<e��ݳ~ı�_Fun��H���j�e~���9���*��{`�0��Q��J�^�	�i��C`|���W�f?Ri{ڀ��s&��͏w����xp�冸7�%G���s�[+�s]��9q��='�Y�	M����On6^��5b��u(6�T�?�N�|����4`X�qPݫf5j?yWH�[�͋��4C��Tj��3��G���6_�rl���5�h�ٔ����9T]|s$�.����*3_��V�2;"�SA�DOz��'�Ub@k�q
��_:��S�����
4�@l�m�2�)�[�G�)��N���T��l��q���1�GYr���4V�g?��+�t�O��y�:o�~����;"|a�߿�`��� ����+S��ZhR
-1"���-�k��^������e�!�)�H�����p��������9���&F��1�:�
۷��r�4h�=���� /Κ,J=wq~�t���w���"���`�m�7�"������t�ݘ7�����M�,��wW�a,��toN�E� 
Ń���Wb�d8���X���s���5ӊc;X�۩A����x8��O3�69��瞹}�c�M\�����wAG�bs�遨GaTE@��s\ؔ4E�_�cFOSQ��p���V[ǃ��ROp�Y�@��"��3aH%��M����5���g�:S鋒�ˍ_�1\����]G fI���&Czcӝ1�x� 3����!c�]M��?1�ַ���JV_�~���t0Y�Yu�o%D█.m��i�ե	���>Z���0��<��4����USk��!R�Yi�X��_:�"���Z�ko��MC��;���I�Iw]55LD㛢��"�&�@����&��M�F��az�����E�K��v��I��C`:�V�P����g���5�.&4�J�H~˲"� �����������!��rY�sF�颻c������f�@>���G'%���,O�3L�:I��ґoW.��}�L��9���ޑ���㲷�:ߕcTC�|��:��Kㆻ�I�E;.��b�~���ozB��P�Dyb�}��ᾅGl��T��
��Vq�Y(�p}��
�������ٵK�E{�O��j]����*�{�,��^�Ũ�o�Dq����b&P �A!L��q��%鄰\�^�%�r"��FdWEm>�Pe�S�s�KĸU�o�:~'�y�!�,��t�3��݃I+[�_4��q8�I��U��GH��[Sk�؆��u���/GzUj�U:����EH�0�K��j��30B};�$�(����P
�xm�Y��}�\g�w��g���� J�3@"�������T>OM�`~�s|'� ���Y�6гhN����O�D�z��X�{����rf|44ɵ�I�;YD��dn��؞YS�n\���	��y�vL`4KX�`J��k�ܿ�v+��;���}�)U���;�`�t�R�nn��jM
t*E����C�S�Ɣ�g��?EN4��Y�$��wrG2�zph�.��,ѯ� !nң��I0��Da�o �g�I�'L]6�O�O�EfʵR>IR[��4�7=Å;2a���܀�r @
�2��!F�]������ҳ����b>R#1tH��r�	47� �C�sz0?z\��ȒXUr8�Ok9ͱ�"A���S ����e_{�ԯN�x\��)GU
/�*�_�+�!����pV����"���%�N-{�ILT�`�{�܉eP�-��J{�9�N�R1��:5E��q�k��������o��P��D>�On�*"V�~��F�FZ�"��<�(�v�k?\-u`z����薚X����n#�xJ�K�r;2^�`3�V�H�i�����q��ݔ�����$�5[�四I��*}�絛a &�Ӈ�W��\�t�c�a�D���_C�G��5j�Ja��m�.c����Q�������f�{yy�� Xc3�v�<.� �8�Y�ՕO�l��~h̊Dx��W�$��C�����I�̍
3H��ſ(ԇ��Nb/�vJ��Ղu�~ӂ�5&��4N�*R?W?�z�)���9B\�/�,�b�W��kY��[Z��y4Z��_*ȹ�,�I�z|�ޠ��E�ԞT%���AFS1��V�X7� �cW����UO���r��d:�	��?�F_�������\�j�u�x����Z7+V���f�^�]�+���v�j(0�]I�kD�ļ��>&�����y�I�x�Yܸ�
��s5�7{~>5��>X�s���]�����O!.������eP�W�R�_i�'V ���g��O�D߻q�"��K�Y.���؇�7�{��t��椩�;�a��)>�ce�g�/N��n���K�/y�K�F���K
��*���$��&!W�Ld�W����өO�4M���\�ƏZ s�e��W������]���C�_�����0JwM������tq�������5����ym��A��߲~+g^��C��x&��iB!�N�gǭ��q���%D�����_τƛ��֞v���9�����9}���-�+��u'��C�XPX߬��ϖR�0pm�h��̚X�;=�E�8`=S5v�x��k,k���_ی�h�i6� �^�,�o��� �����qc!�hBu[��ײ�p�C�ՠz#�evJe[Ȋ��J��6��27��H'�#�[1��q��>.Y���z,9�_�S=�U�H��mj)0M�=�J�F����=�/�Q�ᐱ)x�(I.A����^��z�!��\ŞL7���� ��vh[Ô{��?�z�M��f�;_��"(ɛ�!�h�丳}>�r�=��P4=�%hs����h��=k���!q,�u�}.:���w�h(�	�+��i��?oЇ>"�_��5,��se�A��G��
+�]��"=5�̬>�up�jv$�1���)�.�k^��J��
���w����ط��/�X�tw���Yb	f��j���6��O��SQxI(v��w�M����<��@�(1��� �5# 8�w&�/E0~��S7ƙ��K�}¶&�p�՛�73̦4��u��~O?�8?0�1�g���;*��:r;��`T�w������3M՘&j�����������ϵ:>����:��������G�kP�]�� s3������ui�4?{��7�FiBO�V�Քu��_t��8:ç�c��8�u}B��v%�q�1?�p��\P嚒 O��s����4�Kk �t)����+~��Z}@`i
����<���M��[$f��P,�%
�Cp2/��V���=>�'zz�+Y똱��XE�:9�*�e�|�ג���DR'���W�5�)r�)�.��.cַS�g�31`(��O5Qi�KN���]ӬI�ѭq�u'U-/��D�����"!�������q��pS�*X�?Bh H�?j�5�,�(�"��%�� *��c5^B3	���W۟�w����u!�RI5,���'��ْ����*p8�g7��-9�^�}���1�~��������kb��N���r�sQ�
>Zs]�� �X����<,-Q%yW�� ��Ow���;���A�9�[7'�tE,^q�r
Z1�uΈI���*�~��5:hW&=kh;*^r�k5�W*'Z��j�G>r�Y�c�EU
��r�����ᱴ�ɺ�n�[��WV�{��<uѱ�'�Mry��-�N�����Lr�5�u�0�
���XSv�=��t�n�ݜS�7gA���ւ�0��+D0��ߐ!��4���/���7N�񀭐�zX">3,v��!@�F���D�9����D6*���W1`b/�"ܟ~��g���E��d9Q��I;E�#�Җ%ѩ?4��x�<��o�X�M�od�'�p Г������8���V(����F�I��@����y:>̽�A�aP�1ᒳ3����ξ^(I��2T���G� ︽�%��v�"��l�zk��Cِ� T� �9���{W�сK���]B����Z|~���é��  ���?���|�"X3�V��ERl2O�c&�չd�gw������h�%���=��*&��v�Q9�3Tt��:\a ���T�F��C�ס=}
b7]�m�5��`5����81����X}�ڼｩ�c��(vW�	_�a�5M���c�P�:� Z�ު̉��Of��e��s��D�>�P�D�OėC8m��w�����F��è�SѳkϞ��	��`�w&��q�	"ơe�^�T�!Hw���(�bI҃�Է��OeD�k����tI��|�g���Z�Z��1�0�W������܁��R�>~��ֹ��^ಉ�"z�&cYۏ�� ��ͭ
`�C����!L�Ss����0;�݈0wB�� ����Mv'wy�Ň���R�O��xa�𭬭k�e��aWIbgHe0���C��J�$a����:,3��߈�{���C�
1yVX|5T����dɏ2,	�����2U�"`��P�P�FVn;l�c%?[\�p���Ɗ}e�?��=��g_������$u�N(���'��o�����(�J�����Ek�E�\Q�'���°�T��G��),B��(VZ���j�9�\�t�|Y&�ax�F�a�,��`.�����>�ͪC�T���:с���mc�R]TvcJ�ق�}�t��d�g��y�,>B9�7�W~�SB?����U�悂	po�va�E!���H��\��n�~˲J$�'�`(z�����z��[��r����Py�Z5�G��������I�����Fn��mT(s�'W�1ɖ�#�{��3�G����P����~�)� �J_�������%I�򈐧c@�ຈ�sQ$�,�ӷ��!��a+&�0�Ea{]��d����K��L"�()�@䈈���K���	��L!�Q�nO9�D�='?�T%j9D���H�V��� ��K�=7��>ص�æd}�O�U�)��8�:��ǐ2$m��T� Ϡ?��/r����͜�<�KkN���G�(hg��R�����T��gzDQ�![�j8��{��4�8Q�'<�D+ЗK��Ӗ����&��f�:!w3��}yXYC	�Y5Ĩj�9+�>
�ў׮��^b�H_�'��������W5C����:�V^z�7Y�_}H�	BLz��6�}S�͌S � �Sì����9H�h{(J����&��q�X��� p~ۮ~g7���\���u��(Y��A8D���*һ�#�����i:5i��m^a5sB�0T��~"m�����P�YRz��E��0��,���'/�T냨�P�u����_�̚�L�Ё��A�r��e��2�֎�wo��?}���b�H���ɬQ�����$�u�_LsWoz�l[�˒��Q۶�������s��.�{�Z�{��j�ǰ��0�M/��WBN�}ù@��śf,��A�e�
��b�Rz����]�e��W���"�<�u%8TmaP���0;/ĥФ�V�@�B�d�a��-1���("]��"�a���! |2�,�gv_D.	UR#��M���>R	���I��;8��Oҙ�Qs��\S���sl���rv���6�F�S;��Hb���R	$�T��1�qeZG;Ѿ35L�ST�����Ĥ1�Y(o���4�v� � �C�)Po�2s��s������
֥/#^����K�U� F������Bڧ��`J���,v4�b~�v÷VNr2/RЁ��D#M�寤����� Â��+_ U��A��ׄ�k�܁p�1"��U�,#�����z�#E>�?&��|�X%�����G��U����=�%n@r����X
ryK�%Y���q�0)�:H͇�`T��)�M����xJW��EbY�y����k���.�e�疔3)�8>�+��b�K+i<y5?����h�
"(D�k�py7w�%/&�\љT9�Ⱥ�����.�v}������xB$�לG{���\�\���_~Ck~i���_v�A:��\�O�v��g��/��`�E�6_��!��l�b�� �6Rcq��sf�/����G�b~��A΢�H���f��+M��l���`}�\1�a�s6�t[�#��!���i~� {��W�!���^�NGV)����KV�|�Z�5v����Ȇ p��#��
.O2��p�	��B��e�$e?a���ꅉ�a��M>���q�R�� LO%��40���s6m�!~
�쉁Tŀ�'��@�kB�$YP�u�5h�"t��A���LMP�w�1)J0b����s�%{\n���B��iu�5�N����ȥW*ʼ�I��b ��,wk[��>n��3���O\1si)�qϙDV� E�w�x���Mk�P���:4�����<�@?(g�^L�钖�52����0��%��ƽ[ �	�Z;�6��?��G{ h�';㠆!�nD�/2'���ɔ�b�wB��C���8v��wS�E1�;qq�Φ�Z�*lXߌ�wE���l��fVvl}ɕ�*���ϟ�;ddt��cw��dDdjZ@c�,N,�(�I�C3������.u��$��.��}��g��LL�͸G>+SC%j(����f'a.S���мn蝏/KO���Y��&y:��G�U��b�W]�)u:lҼ�����=r�^�������f�ROGH��O"n�.���FQ�V�wv@1�Y���e� g��V�.P�~O8JT&�7�7$�U b��E=2�A�"�+����P���t0~��T�ZX�P��t�	g�Ki�_5;��Qzi�u��(��}(@�چr��2߫��2�1~�؄?9���9�Aͤ��r����"��KeV��a�tX�n��3�S��m?���!��[�|^�>��Q;p@�̵�z�w�6�c� �$;�x��šՊ���
# �g7��-B�#��� �\���#݄Q8����5톆hH�Z�7��0�*�G��0�5�7FkYD�x�$d�j�B���_���M�J'EX(�-�i��Zj��zo�b[�@p,�I�D�=��kQ�f�1 {^Ĵ���[�F`��.���@+b(|b�4iF��;���}ʄ+��V�}嬮n�'�8�	��_�Ϭm��ˬv���f4���6V�7~r������ޘ��=N�Khр,2�Bc%a)8?�}��,o���E��K�k&��@U��D/�
H*Xhu(����Y��>����O{4�S��-Kg��d�h����H��T�X䏯�H�jX��W� ��=V˩��
�T�e`�UN��b2G�kV��7rłX���/�?^��u��4S��c�pW������z��+�J-|w���n9�7z	�x�'�]F�Ȃ�Q)/!��:��&ib�������Xs�C�o܈�>-�%qZbB�_*Y���������*�ލ�4�1������a�u��Lc<�[�R�k&{.�����g�FM=�Ђ*v�b�9�b��X�{QB��v�����_%ݵ�χ�s�Wp�l>?I�dOn�� YҊv7_Zn����=F6�����7��Z��;�J�����o*���e��ϯ`Z�
�-+�TuWX(9�(��I�N��b1���|xs��Xqn�c"W��\(�ׅ��{G�|�E2��z$E�!-Mk�UN.�N��o=��Q��a�b���GsX]tS���ո�!2�lVnFPDo���H~��h$x����+X9� |�Bh}g�O��4��(������Q8��r���ϩ�O9,�/A�ck>*K_��Z0˳cSS��M�H>ϗ�'��P�e]�O�_�����(��B�?rEY��w_���N��/�n��{��n�Ѽ	@f%�M������,�#`��H�h|[�ّӵ6	y���U���r�e2hL�+L#��^E�ʬb֛��xl�a���?�^5]N�Z�Խ?�-�X�9�@�@�x�oԺD�+}���|�Tl���-$S��$�|����@*Y~�1�L��<K��ɤ&`�F)\�sk����䔞KMV9W��M%h����h]= ���C���F~�Y��?Il�-�"3��)@�A�cbn��?O����]�;�/�������a���Iո�~T�Xm\�q5�)d��
�Ǧn�I��7��y�ʜ#�;v&������0��I��k�N�{���Р��6��s�JD�䪼�|�o#%	�D*O1��e0<~{��7^�j�����
�]�d"v��c����]E�]V��љT(����hVxg��pa̘����֯z�.+M|k��E߾�F�o�D�L�D"�����Kw<|ҟb�#��T߾o.'�ǎl���N��_1o����K�A��L-��1�
Pa��{,��;Tq�%�m���~���W5"��g��ۿF�+��.��#�b�o�u͍�}�0���OE��s��{Q�����/춎�&�1�;2�����Oۂ���I�����/[�6���5�v��(��O��s�Y�PZ� ��o��w��G�OS���q�����g9zË���nf��-i����0�b�k�nx��S�wjk���[�����i�{:�W�6d9K�������_7I��}�ߠ�I���F��g����~����lM��;�&������J�9@]q0eM��>�{��|��a��1!����D��� <D��I*$k����4��05�8&h!�a2}���F�1��R�N_>���"R[�]�^ L��i���.	�\��A7�E���w�`���^Q���4{��y!{���w��'�mO�f>�'ȍ�,C}����_��#JɆ� ��9���a��7���.c��7&�s
�u�^�{9˃�w�o�9��36��-A.�5�蕙x]� V�	Z��WK!ƞ����W4(�ј1�&wف�r�yM5��.<���1�]2+�~�V�ɻ�X��T�䷓�}�T�A�b)G^J��lN.E�ybd��	��=�����%fq������Mr"y",�bP��T{$� �"z-<�C��ޣ�:�R�@���
�u)��b��l�23x��ӿP
��pш�{_dh`c�7��P
�R SZ�O
�3���yd��q0��z�s�
�l��=n��z��I�����R&-i9U/���ky�(�2Ǳ��Ǳ	;,	����$�·y�P�?}!.0����W3���a�S`EƒA��~�.M��՚�#æ������z�, �`�JД֏h��*�v�#=��g/�>'¯1J�c�1�e�Հ�ث�6p� �����c��{�v�7�ȧ����ŝ�]]��<8������z�`V�)pOR���ߢ��?ի�"8�},�Q��1u�	�Mi���܂X�}�JY+�x�˛���a�Os�zOD��5hn�x�$������.c��#�AS�v
Z�����_�6�x�N�fh�IƇ�\襽��G�7���p�h�22�	0��+����� ���I��OZ�ULջK��R%��u���9%jd���ccchDq�V�ѧ,=�i8w$��Z����o�w�O�f�R�H3,u��wj?����[��\�Y����_7kA��Q���r=�5��4��� 8���EQ��^�=����7�
��Etb@�[���ÆKp{q�� �_����	z�V���СȤص>
��s7����:�: ����h}��nǗ���'� Z���=`
zP�<�Va���w-�>)��I�_�
Aљ'�/��*��
7G�R��+	��ԁ���J�ʄ,����B	�.�
ſp�뷢UxwZ�,�,�R[�f�l#����w���$��)0�;s���Q���ݺC��Bނr��[���'�X��N�u�A�|�q���}�p1|��V��t�8"�B�P&t���^3���H���N��m���$�yє񳓵�p!�,V�2�D+֏��s��2�����#����ȉ}~v�#u��zI U�3�W)�����<R�s������q��$�����!;�hj8�&-�\['f��L�ԗ�̰��C0s�N:���}x�b��͸�(�$@1#��=�|^��Z�?����	����m��v����WJP��ca︞�t�L}������1Lzr�_��������	2�ZE+���~,��@Oq��EQ�"�=��Ӈxs�	)�5� F$�Y�3?��M0��!����B��x�B�ض�Q�T����ۖ^Δ��9D�+�b:Z��(v8v�&dh��\]���s���S�}!��)I��ROR峥0��o�cR�l©�϶)�����Q�y*�P��PC ��g�����+����/za�M�~9�t�#!==bW����ڶC�̜��z��:�poM��CG*�m�Oގ�lLQ�Y"��	�@����'Iq��]n�dpصF�يḫ�e�p���_�n�����0��
×�2,+`)���@�p;X�{4yS��WO�$]A������C��@o���3�m���1��xd�6��7���-����_���U#}?R�<�%�8T��HmL��G��;���
��F�y�|�Ƚy�u�fQ��D�{<����'Q��Ɛ.hX-��r�#LP�L]*��-P	��e��=��{mtt��ݣBW"��v��]Zwԣ�8�K�	�F�^�H�7DF��d��r���v�`J!��	�������2���l�����A���\DG�����Hi��:�]S�^�
%J��VqXڪ�2�a7��CY��	֨�D높V���-T�lNoԥPS����� �z�՟�����B�	����b49���^H����:zA@����C�A�e���k2[�v��u3-��&�h��S�9�@�bm�IS�E{��G_��<@��vB���n�e�R0�~�L������WX\U��Pk���7�0�Rk�!�LJ(�T.�HP���]�4���T��E���.����i��d���b�����(W��4��׎':z���<�.�n˘F�x��UBq4��ӭx�^��Z��R8�舛�9\S�Yo�(z�.t�p�d"۫�I�=r�\~ (W^�b��|c�U$6��g��j月�`�Nɶ!Z�1�Sg���F�lp!��%Q����f�o�'�t�����|��c���O1�d��FU��+҄_�+.��k�}@�X�
'��XW������*����az#dj����q�)+S�"�:�b��[�/J��\��e{�@c�s��t����7K�m���v��"����q�:>bs$�ؚ��S�2f2�i���ZI0	h!�_��}�'p���ק�r��,��$!Ь���<�㨌���qK���ܶ�i d!7�>T���$F�\?v4����I�xε�0��9ny�ў�\��͛p�k&l��e;�#MRץPQ���3hZ��\k����d��C#�f7�1nflZ�<�{��P���a�v5�D�UO��訖�.�^1��t��5rI_�U��1��<��ړ���N��=xT�8�E�+������9��8�Q�0���g,��whs� ��[��8�����������s�QM���y��~�BM��;�ɀ�h��b��J����-v8ӆ0�.�m��iR�R�(b��C�G���^1(���?s"n���]����6AtV�:���Õ槳XӮU�O0f�0�$R�$�7=�!c��D��dr�V�է����{�5�T�µ<��tl6>����JR���;�LPa�Nu��� [;du�Ql{\p
A-ԍ�U�s�׽x������o��g��ѓЋFL�LV���\���N��\�l�2([��JV{���%-���u.~�j&��{�8��dZ�3,�@��v_R�:��/8�x3�`;����?�� ���5�h0r[:=���ά������ut�^�)��oR��c�8�(���&����p��=�юL��xX漞�\|#{Ά�a&���C�K>"O����,��i��W!P�jc:<���;)������x�"�n�-IPYd�27�b�n5E����}����$�;'A �ٸ7Վ����~�����*���{\�v�3G 5P_���?i(̍�Ŏe��-�|Ʉ_)�쮓	/#}F�X�5WrF=ɧ�*g�l��0ލE&�(?6�
;�w�����j��2H�uF�('<N�)C|3(�N�������w���P�b�����ɬ��+�"`���Ph�0gMg��A����wu��M4���o>����úꧩV���B|�W ���]�q�}�#lꨈ�,1��;�"	���[��6�B�ɒ�׳�7�e�(�)p���=��j�����M ���'AF�Ͳ^��Q�O���$O�Y��|�Ή#"?s�qj��}a�UY7������H┆alA��^D�T��Z_p�x6ˉ'z��BL����E>����T�}�����"���I� �p^�.�՟�(2� /]g^q������U��cm�n�� �9�j �H��>G!���5�QP_�}�K<���hM���fÛ����\���t
c!�2ng�[�3�&n��Dd�1�m{�gw�s����G��p�m宝A�='Y	�n�Кėf@���"v�EK��_�����c�vP
3�j`������f�q	8�K��ƴ�'��5X3����e>�4ǭ��lOcE��Ulc�|%"}�<@��m��۳DᲟ��Giv��`��d���>��a8P��C��r���#-����G���T�q��&���ף��cts���աY�� a��3+5%�^@��4�nS/c��H����`\�G�=�i�_t��;���=�yq�\|���]�:�[`qt�/|�b"����׳訇���|h7k�to����F1:u4��vʟ����X�ÿIkӁ�9*P��(��HV�ߌ�,�B�\C/��?Dԉ�ϛ��ޔ�W8����L���~�σ9��2�I�F��6`fS��6�tG7�y�"8����Nz���W��_>����vR��6�8"��P�#I�Aa6ݾ:�V��Yq�a�)�����IM����E�$�_�*����_+�*@�g���Q�z�E�9��蝟����������/������  ���r*��
�^����dB�$�����x'���{Δ6J�����@k�����>Np!��˚�������4�߭�����oh����/*�R�xD�J��Ѵ]V�Ӥ��:D(df,7��jg�ѻ��k�Z�Y=�N�v4QU7�ւY�?�F5B �a7�pS�����&���#����~0^�pi�-\�;QL�.��Q�U��]N��*M��B����7MJ?��?�!FP�?ʕ���u�z�"�Op\�Ą��FćnE�]@h��X�`��Ӵt��/���@f�L9�su�B�~P�O�n��1�lU� �I����֖ph.&޺���(�'t?�y����`
�/0�Ұ2td�#L��~r.�U����Y�����}J<�Cs$N2%�j�՝`��ɃI��߳��L�N��o2�Q�gΉ�V�ټ�[x,l�_7����-_�8Y��?܋�+nt�fH�r�0fk�΀��=!��&�8`�Kn�2��r_�;<[�� $��ܥ�n�+���egS�gmG�'�8�,Є�4s�+��Vf���8[@��.?�o���,c��d��!RV�����g�
����=h�f�!
�Z�G����M
��C,��͊�cy����.R�-��H-}S���A����aY��,� Igf��8���z�2Z���ݣ�0�Y_eڐ9`��_���}�[��+U��.��_֏Ȼ�҈ebTW�yj��(��A�N����NwH���U��hAxi��Ӣ�� K���,�.&���D?�x�x;nU�^����=�QMz�~([�s,?�+������q<�}��UZdS���p�+���|��ǵ�ޞ��I*MZ��F5���0�H�&oN8o��܆p����2A1P�g�f\SNz�xa�
^d�67?�{#ʻ*ad�X����I*�|o ܲn�K���M�� �K���D-����%����4�j�}���k�E�Ax#���@s�D�p4��5�v�Lvc�R8����{)�}��l>��}�d��r�����g趴���GM�A�������	k*zw��E�3��|�C�g�0�ĺ�������������S^�L�Fy���eJ���i�q�2�a�(U��0b�|�賩����4u�����d5{Qd+��tOZ�C\��n�k��I(�U:�Q��Â�I:�d/��1tP�-!-,CP�L#��=�*�7�D6W����kx���p�: <�M`�G%��I����F��NY��aM��ʉɥ� C�."�hCR���t�����Ω��M��"q�5>��ͅ��(��?�f�}V�����bj�'
9%��5l���vh���f�hȕ�ml0;���V:��Y�(S��!��9j��;\ԫ�:��Dy#ܜ�Tಎ���	 a��ş^��I��1��f������P�(�65F#&�!������0�@��cz��$��[r�*����sG����S:����{3��H����9^o�]Y7��eו�=��=h U�7�܎�E��y�,#��Ҭ#չ�D����j�	�'4LDR��fG��z\�4n�8G�������B�@B��vjw��ZP?+,�1���$�����`�z<�P呬 ݶM��?HO+�������p�آea-B{T$Η�<�kdP���R�~��F�^��%�6��7<p�A�x3�x�9�5�Wi�<f*z�8r|�E�[F%���	K��PXeR��B%�ĲP��/\�d�9�J�\x���hU@�o"�����XĤa�!{�IU��'zSLF�ZJwR�x�gt��/�B�>\����治h��}��z�����?�������X���`�EϖCa_��>�@��tb�!&���h|υ)hv4���bt��{�!�>�����e��R�
���QS���{�.�b]&����.gy���]V�*j�/O����]z����I���Mv�-�GD�!�@����e&P��J�������;u�!��p��hg�AH�]�vez��	7�X�Y�&����~�l8����	�IU#i��2�㛙��1L���3�ג|��A�S�w8Χ��R�(���
}X���E�h~ 1u�OK5�[��[���ا�OS�3?�)�my0�zS�������0��$ԾV���^ڙZ�5��XFtdM�ZF�\Z�R���-�O�&�L�폅"U���4 l$X�ː�a���+��7ha���D�vm8�{��'3��(J|�n���{ qE�\Q���	�In��/X�K�:��v��:�\ R�ٳps�4EGU���WY���=��hRz*��ʽ���}���������QQ��Է�N*�hg}3����ƿ63 _��S���`[m�vڼں&;.�~��j�G�~�_�<0�Y��kӟ�1%_�I⒤���@UM��.�\=do=Q-��͚���_���G�ߚ�7��*���o�ԡ�#�!���˲��s�r��#Ҝ��V>��� P'�.%|���,#�R^}��6���D�Z���o)����,ᮜ�� ��;��3*+��)S���~�㥿5Ə	���@@=Z"�����v'#�[r�N����r�mϻ�������(00�G��Ÿ��F_������p܃��n�T���)�#eU����?�0*7�)��R�@�+��]�Ҕ�Gw���4�zQP�8�Q�}9�'�RjV� ��.�թv�z?�O$��d����|P���B!wJ�,��fhg��b�bv��w�Q2a�����6�?x�L���v���7cb@���F����0-��Q�>�2`1"h��	��i���Du_�0y�kz=ǅ̇8�>�α�l��A���u��a6wtͱ	�b���ō���֚9V���;1�V�x(ϝI���'	wm�ezJ�����/��}�X�렿;u;�l�)N�R��/.c?'	m	���\�4QA��x�<�Ae��A�G�K��*�A�+����5y�亻S�&o]�bPn�z�G��<ʂ\��옮م��"Wy1��(s&�wL�	Kň�E�+״���3��J1OG��Bu͜L��Uy;\+�Pn�!b/~����_u�,)��8o��q3b�0��)m=�E�<i�7�ts�і
�����T��/h"n�>'ە��)���roǂX+�2�ʋ�!m<������!%[W��|���c�j(rF�栃_q3a���g����E��T�?��o^gk\̿��9������A�#�}��D���֑���Vk��N���(��5��42p[&�s��|�������*��K ?_����`�á��\%��vY/�׫�/"݀;�򈪸�5Y���~l���F7{��ouq�}?�N}�EK7��/5�m]YdRr�zɟd�l슟B��#�Hfj;�}YںD/D�9d���0�X?l&[@��ȕ
B(����Rǝ��D�5�ĝ�0ވ5�+�n@n��	����>���?����եxH��`��bm9�_3-��4r��y➿��u9z�X�2i[Ĳ[a�;StX��v1��b�&IA4�$�qqA_��h�I��Fa横Q�6!7]�&6����G��L�uG���f�-�=�L2j|KGM,�M�9�ۚ]
nS#�r�M��~������^tOTɊ� ?�>�>>p�@	�;��VmW�Ĉ	"���*�B�"��,���*��춞J�O>K��r���vt8_}ݮ�0�&l��莭�*��,��L��5�;�V��N���oPc�fM���y�b����]��bL�aOg��F	�Qƺ�Lͪ�� `��>��L��o)��T�fdĵ<���d~Xz	�I�ߡ/�TV{��򞺀���?7Q��:�lp��J��*`f�zq�9Q�5(�_�`?�;m��21�t'�
�R�t��!�^K��U�ܸ�#-�3�\�	�e�c���n��Oƛ�q^w��J�O�S��Fo����XV$��ٕH�I��O��`x�}����=X��ۮZ���- �UJ4�X����>ݹ��H���k�;�x֣����u��ġ��"�1�*�k�Yq�c�T&���
qV��"
���.{�bƷ�@rG��2�N������L���_��N�CQof�� �����Ծ"����`ٯ���=�u���U7�u���N|s>�A�}�>��?y��q�ڿ"Lf�-p��.�Ŭ��/�u,f������h�S�8j�F�(w7��(	�s��Ϸ���ͱ�S���Х{���P%1~r�yb���3e7mBJ��D����
\��6���Y��$��]ڰ/Ȩ<A'� �ks��7|����*=V��{e�	<�z�U�X������.G������noX	���QL�����
�)B�<f⺴Ꙣ*c,c]M;�s)e%�TI�*�j����Qѭ�iA��s3��m�V�ǥw�@e��(~�\�&�1�U����`��̞DG�) *ʃ��kw5�<_�?'�B|DO�W��ό �ǤP�>���]��G�`�!p��}:JaY���
�;���%i�k�w�8q����"��!��:)`vZ��or�:*J�{ {93��)��V&'��H�̄�8��b�J%ơ�����}���E^5��9����0��Ӌ��7Y7�P"��KȂ�30�`���A�@���ǃV-v;�Z��͙<�.�*s7���L���Y�Av4mּ�_G$�ut>�po;��A@dy�9	DDu~��0�:z�Y�49+�a9��UÝ~�i������p�NH�_�/U�*��T#C��>0�����CO&��2N�5��]TtzlU���FJZ"�d�#hlo�DZWm���%9Mik���_hJ�b�V���T=1��dm/��p.�W=��� �RD��7� y��<�q��޽�	5q� � �#9Ө�2���ۚ���7-}h�u��m
��J�G�U���A����v�p�
���ن[i����@>��s�.`厌�y(�*\�zY��ـ���tJ� �����<R�r����t5��s� ږ������8���.��w�Q�ZPM�K:r0R|�V�0+�D�~ѭ�������E�~��%]+m���-Uf)hD?n���=���9� ���������B-F=�#0�[:�	!_�Vc(w�D����ƞ�㰲@֨��q�6�ϋ;�-��D��7&qh��$�a*�O���sF�fۦM<ޭ��з��^��;�o�G0�<��En0�&�G� �@d�5�Ղ�%=X�1�FY({��&��,���35�4���Hy�=��_����{O7��Oڌl�c��.l��=$v�ܯXd�z�ΰ��4��0�r���f���r�k���d�.�5g��\����Q6r2[%jr�F6��g��:�,B�z�F�[��E�3��7����8�<�RrBʏ%ɴ6k7������־��x�]k?FJ[�d��|����o����l՚��ns�n�O7�(�����F�HǓH{h:2a��ŷɴ�p���>��`���*���
9�~�6��(ʴT�k�1�?(��f�(���۳k����hz��&��;�!���N4 @� .����z�tX{*r�j9��@e|�G <��LnQ-d��bBxRS�x5�e霿҃���؎WM%ʞ?�Jg�(,U'��I�L��dLQ|s"�>��?!ZxԻC��s�.g�ë��� )��铉�j'4O�qN�z�<Tpz>|�/N�Îٍ�(�/ɐ��G:�U�~p; ���g(d�S���m�'":S�ݓ �eg�Dv�Wh�;��o=�h]��ޗ�Wmi�����Ug�X]8z;8�p�?J'Y��	�t������>��F*hL��!椺0�N���5h������<U>������BDy�/��C"���-2'�x�ݕQc6�=�h�ְ�>&#��g�M�ȟ,y�'gP��+s�e�װ��t����R�Y䈚*�O���нXL_�nN���+Q�?�Z�y������.-d�]O����>[.h����y�;L��oCİ;��i�o5��?g�E�B^�m��KS�ϗZ͙]�鿆B���Z]�%ʢ	(��f������m���ɢ� ����a4N<�`��.>0�yb�=7t&kvޟa˝�*�^8��+���,�x\	�N�?�����J�e�3W׷s�ꮎ�&��x;�ŲW��b���u���6�Z���1�.6����)�م�m�8��j�>�K(B���eU�Ւ��@��{�]~���F7�zwc�?a��a �j�JTJ��
��>}{%��_'��$m�������y���he�Хs�?�.�jޱ��7���a`���t���w`���lIڌr�����'&75I��'��^,��?|y������}w4B��=�D+��b	�������o��?SB_�ZkC;w�U�;��S ��L�K����틒�Z�H�P�K��B5�k�a�9V145?/�+����_j"��|
k��h�
R��&�9������w�u��]�+yo��!���og1�/����+D�.^���X	u������p����E6��������#?ep�f������+��Eϗ��^|���;v��0b�u�c�~��*Da����R��~*����|8�����M4޳��`m䳄���!�@G4��jR֝�i|L[i�Z'e:[K
�F|5�u�>Ts�����V��IwK�5\�X7p+�Z���6Zp���Em~���O��qU��j��j��ƚФ�����kc��Zl����ۊiq3&_��dv���'
�FT����-�e��+C�Ǌ��"�C��M閕�������q�h���݄��GD�嘲�KM���WS����ń�_�Q���2d)ງ�-��sA����y���
�)Z,�d�y�5pJ�
3E�dy]<���}z
���f�F��-�;�����}w� 4u���R�%ۮ��r_43���丣����ۣ����e�X2 B�R�Jϕ3�ﺕ�(Q�Iޅn&�āX�VP��
*��} ���B�W"��=��/҉���zp�����M�{ٝ�A�R���!��)].F�A�\���L��I���W�u)C�I ۱IBP�ϰ���f��Z-W���{<���Q�:��=��VVd��*#D���3�����!W��|��4�Fi`d��i��p�Z����c�5o(���W�|8��Q�w|�Ku(����*؈�m3�*bii�K�*Y
�C����#����~�95ȴ��7����Q��~�(���>t)�n���v�����]\@�6�J$����
b���ͧH��P�b5I�sȾ4IZ$l-u���m��,�6���Dղ�:���'�:@�F�����C��g����6�$�df��� o3���m>q���V�B�3��Gl�í!h�?M-�Jޚjf����T뎃�����?�r�no9zX*]=1�ڂ+�Y56'3O�4gy	V4��+dm[&��s����"*�@-A}�̏*�G&���Ǝ�e�x�Rf�x����s2���x�9�ea v��|���Q
��)�vwѦ�,!� �@5�~5A֡2Wӌ�¿�R<�VD�If1�%0���+��7Ęq��(�4�M�g~�ߦ\���Ё;f��:�(��Q�}5 ������e�>-�G��E�+�ͭP��k$qoA�B�۞��m����~��t3h�7z�VB��c1��p�^�+f1�٪�������2`��n�SpwW����8��3����ƕb�(Ƶ&G�7f��K�Y<̠�R�0�D������#z��k�d�L�xel0*�m6�}[p��/��ŵ:F��~
��k��:�n�����d�#�8wE"{N�H�s�j��M�B6cUӓ�b^_ؙ��<I�y���wb�P�-s�����x�=���ϫ]��ݬ�TS�j��^�XJ�\J_�]|#)Ȉ:]��}̍X'��@���
���%U���,]��Q�/B��_}�@�k5q׃���xy1/_��W!nm4B�x�����,���f�;��(͐sz	�S:�o�@�Ÿմ 0e~M�1".;�U�^0��� �tkvN����?E�6U�V0���bR*R�1j��< hu�#�G�F{��� ���2�8�<�/ᶣQk��f�a!;,�O������4��&��]���	��n����`�r��o��k?F&� +</��ñ��vU_�:�e,X��c���|���^���f�f�y�V�V�F�<O�U�+N�۸�C����=vYq� ���֦��N��j	�@����<U�U/e�_����2|ϼ{�7���h�F f�ۈ�z��Ih'M�� �X.���?���=>��vq?��O��+�Q��>+>��87�P�U����Y/��>����u: -bJ��{��4^ĝ��������3�g�v�)>��B�����A��������Z��Uc-�r���R�ݰ�:�fK�� ~ќF���z0d1|$����uyx%����]�N��d�bw2������i�`9Kw�kB�����do� P�����{f���*��O�
o1��-	�Z���Y	�ˎӭ.��jFI�YI��Rh����[t��>�H�����!�T�L<��Ǎ��X��x�B�3A��(C=yq��
�(�$�L�L3F�	խ�[r.H�X���l�I$0<!��l3'e�}�O���[�z5���v7:Ң<��4i5�"U�"���m�sWqO\�����q���;(��q�.����?��
�p6�I˽c6� ��gW��;u�r@S[��m����I�([�h����)c�������\���P�N���K.�1^��]��mFߕ��0����&$�~��I�q*��T�k�c��=�P��+d�t+�k�!�֣eN�Uz��ޏ��%�����L�9�/":2�;ov=q��ycW���±Z$�V��&��o�L�s������ݹ�2!Q��>���lV��;Ybf%�3�xh�ę��:�M��F�����2.�5���]�V��BU��JA�8q�w|��6P��/�t��G�k0g���Rc x�J�)��c�v���n.��k�K&�������p��>'�76��ǚ	FB;܋�b���ko�&?=��$�"�/�B -S�jj�!-A���G�k�ԅ>O�H�ڇ��Ƙ��y�v��:Ŭ�4\�\�B=��8�j4"e���x�1���552vw��e;��j)��|b;�ra7���I6V�Y�x3�0�X\v�~�E�Csa�5�^\L��z�Ư|c�Nl\�qE_�_�
~+�Nk�_�E�%�^������C��w���4��3��O+؎� .H��BdG]_��F��!�h|5�\�<����пҒW���?�1(;0k�`�2r��#�l�6��*;a�,(`�zXޖ���=�U>|��E��·H�t�MI.�HЪ�v�
�tnW	aA������aE�����Y�?�GR� ��ࠉ��rh	�C�^e���T�b�cf�Y�*�w�ħ[��ȞQ!RU�~)�l�B��hM�5�u�
ԃl
}����t��:*@m8'/���l�`�x4�$���K� ����N���"�%����BT'���� mw�XMP�~����n0%KY#ߴ��
��jH岿,�@Ct�u�׌�qJ�CFx�DJ���
��r ��?���7���ӏv�4l�^�/�����*�n;��.����Rͻ���4��Nk`������Uu��� �ͥ�u{dW�lx���7Ý��n�X-іs�WGh��G���~B�6�
.x~��	�kk�mYY��~�?��֗��3M�b�W	O�6�c�r���s��[y�']�X0��ɇ�oMNLW����!����P֪�KP;e��I�L0�7��!	�5�R������&� �'������ ?�o�$T�O)������}W{����nŠ1�g���<���6�4E��l����F�����j�Z�+?�'������!�]^M�}����P �)g�J��-ҥ�c���Բ�:ͦ��m��;3R�����s�*�_��ի ��!��hE}���Od����O���8f�gǵ�$2�5l	~�W5SıD�V�#5��ˎ1��DH)x�\�zr/��޽����]����#s"�B��%&�t����A�e�Y����&3���_��݂��+���S�:���)��+��>�T���{�<\�@��c��uO�KؔXi��>Rl[H(f��^��&D$�f�s�J��+�w��+� �9<��.���� �0wz�H�ǫ'���N�]TPZ���U���_��{^���*��~�-���>kI� &pɲd���☃�;����\�d|�h�5�=[j��?Xb
��]Ftܶ�B�)ݪ|�k���N7z���}+&&��[�I�)����wJ��rs�����x���4�R)�i[�D��0�G�*#Q�1	��OD�m_�C�/��v~,����u��KԞúS\TY�K_�h����x�J|��}Ԙ�>f}�J$� C[�5l��Ʀ�1 �(��F�g�lK�~��<95�Y��-fHW�"�8�'��݄�M�#S��nlj&�tI�":HܠFZTy��-�<�&�י��:��n�/������{�Kk���U�� ��wu5�vk����r����EĔmT����h����Ⱦ�^��9� �F2� 2X�)�Ԝ���]��M;��{7�~��o_��]�k�ц��xODsY@i%�J��W�#��Q��R@�W��K��Gu�[���[���W�����1�:#��\�x��d����A[�_��]d������(��ɍ��*$*�:�C˓vָv�_PS��,�nbw@�[��~�j������p6.\�H���k�$B%��>?]V8Z/��28~^ �U�X���(�o�����"Ck�Q�l��������ݫ�
T��NW��)�i
M�q����]No����ؼ��zV����V�ڕ�y&=��N�c����{��Dx˷��m0ģ��ܱ1:�B.=/�f+ך�v��Q�c�(F�]0VOCx�I�f{vq�z��]kw�&�`	��a�#�g@lW�c!I���#�f,}�ذOx�|���A(���}*3�����{{�|��b�26 B|NN�7�b8�Õ���A�-��V+�P�j��T߳�x4o�ަ]���"5׮y���RB1
O�~��	ڛ���Mk���m���سɩ�������Bxð��-�=��i�:I��u��^u�7�1��0R_`�N˞;���n�w��Y!�M�ٸ˅���򗶧t�V�/L����q�H3�VM�	
��Q���z?��D��� ����&qZދ>����'v��P�*����V�ƌGJ�?�t�[(�\I�s�۰'I�ɢ=�;��Q���"�v6-�Yz�V���_Q����W��-��A�Wʟ�t��0r]<#�%���{�VV{�O9�jw�%}!t�+{v'����7n����?1e�^���}d0R�zǢ���^zvF/�T�JY��и*��q5.�:�cy������U���BtSO�p�{��R���U�Y��A�������:r�Ym
7F�
Z�E�(�2:���~|Es�	�V�/U�8m�'�`رL,J�
�r�Gv��di���'�2�&�
���ß�hk�d��`�!5#7�s%��<��	��	j\|�l���כ�r������@�t -n�V�X^�,�����7�j`�6E�Y�+�;?���Ϊ��W_\v�I�!�uB�<�v�g_Q�U�5*U9Tʫר{Y�mv�"�����w�ae��.�ʢ"��S���T@nu��80�j�P��~�|�)���4*�t_�T6������%�[o �'�f�Ύ\x����5,9���[]�OY�ma^n�#r���-���<�My��8�����a����T)�<z/��F��(��,SX8���_�W"�s�6��r���mq<�f��鸱�������\����]�e-�\8i5$s+�� ˸Oګ�!f�7��p�s��������Ψ5`'�AT)�o(,�S��?#�r��@�P)xn9^�9f��V���S�i~��&�,t��#R�pi�c�#�cHj�ʋ�ݟH2��ʦ�ุ���O��-�7��t_��/�|�.�<�K�N�5�?�Qz#s}��ٳ�\Cd�ۃ+���!�qPg)������r��t'�AT�f�Kܸ'
ʹ�PZ7% Q�u4mą���E��i��冣�W�ܖR ��X��̃j��8�,����y+ɘ�Ծ)%Ԁ|
>���qM��Ҿ�d��cκ��3�ZK��rk�ݽ���?5{��v�/&;�i���kr�Mq	E���aI����R+z������5'C�>Υ�������F�u/7���d�bn�_�-�� ��Q�;0�Y+����e���տ8%���k�[���r���";V�;��!&� 4��ȷ�ꇺɷ�0a���*�,ɞ�F��ۓ#C����ǉ�ֻ���l��*VӃ�.�A�@j��^=i�ף����+��KN��ϋ�P�{X����􀣰�rt<*�r�+뼉�Q���/�ȈȤu�<Ϝ��Ҳ�	�f��Fi���b�q��ƣ�8�?��2��ix�V�:�yym��]ҽ��%G��M��X��̙���j�j)3z k�D+0�����q����qXE�:SƳg>l_�֠V���KpT9�3`�&���c-^�����o���e��92�\�9~r�4��-�ǖ`B�#�B�Nv'I�@&Θ���?�eV����HB/Q�n����ٴ�l;T�)|���w�+�V��tB�y�>9�f�>�Q!�p���غ�OX+��Y�4#dq�"���#��g).��5p�e�J�/�W����@�C����V��,�`^�'h�Y�ƈ�3�p���5��gؒ^�(Bm:��^܎��h"��m�b`&��,� ��y.xM{ch��`� ����z����u�,<� �h�oY�O����Sip�u�~ ��lX�"0�h(� vf�o�2D�P'�G����iz�r��[+T*��W4q9غ�)8z�J;s���ՙ���
�7�z���հ`{^��#`80|nJО�vW���̈$R���NK�e�N���՚�2�"��nR/��b���o�(�~���c�iOb%�>G�L Sd�@������C�b��K�����̫���Y\�a ��2�ݾAZ.^�'y���`R��$�iW�3��S��(�ꐫ\E�$�8��Ѕ�/����z2�Ϧu����k"�	Az�B���D���ū˪���_�S�������Hi2w��2�i�֛C����7�~2�}R�~�ο�c�*���!�sa��E<���[��%��#��]�,|�rH�~ŋ��f�xA��pM�y�t�
��u����
{R&qa�ɠ�+�sc����_b����%KĶ����|�؏��l�R^�� ��Tv �y4�0��[z�z��? ��:KW��3]Dkdj�����+.{���>�@�����ۊ�d�B�`��))���)F��k���+â?Z@����QEF�&���I����'�(�ӝ��[�y�����lk�@�rH��i�[��8����6z(��2�b}��!�/8lȪ��8�T��u�G��n�u��x$_!�&�8�ʚ�F���V*OR�IF+ƚ57#��t�'�D8�6�\����2E��ʴSie���;���λB�Y0�χ�z���@5����2��G������8P��.�3S�};�n������K�g�Я��o�o����/S��J��n�/���G�z��h;g��9p����j���/�%���J�x��*��g*7�K���C}���)���׋��	N�ΘG�(� g=E�(&���MĆf{3d��҅ɡe\4�0T%J�� \�F�tcg�b��:������ ַc��������"uȇ���\Y�Ei'G4^�Nf���"ְt�8���A�ց����;�|Mڥ]G�eu��%e�C��EϚ01��DͶ��3ː_��}iМ�I�9������E��m�����~�#�Zm���I�.P���MW(�
�l���EH(Ǫh�-�bo��# �3kH�::!���q����g�%'m9h'��PĊ����-�\5��ͪ��9�zsG��5{"�)V�a�iE�*!�d�{*�M�S��/�����b�r�Hj��,��ld�[,��n�9s��8�:��!CyH�B�e�F�f�&�� ڝY\�y/9��
�-�m��I�z�ha� ^�x�ҽ�k�0�Md�]�Z<��>�.��o�4��OH�>,�# �W�޸[8��N=M�E-6��&�>�}	4�ANf�I�u��sٓ��D#��1kI��RJ�Fx�x� \�m��ۦdE�f%D��X#���ț���n~7�9�4|V�:(��x����<3�.�G}r��Ov�]����?@�P�~��AF��pg��FÚ�����'d���c�}�W� :�_��qI�A���LS�ၜ�:}_�"��p��k
1t
��OkHrk����v��]<�}bp����� �����6�27�L��0"cP20��?��*�$0�L:���7k�� �q�����3��s����LR\��8|snj�4$I�B�����]ZZ�(��o������ �֒|��Xwo�9�L�� 7dF�c��ry�C��T1��OP�/��r&�o�&2Xd9͇;0!/ͼ��%2-r3ٸ�sp%�>:`}>������ہf3	�o3?���a�#��dޯrW���E-�� ��-�d{9�r�
�'����`A�������
������_y7�g�Z�l�]Ar����sI�\8^�Ŋ��?]m�� ~��324i�}z����Q��nH] v�T{��^gRη���ޟ�Ϟ~!�d���f,��|�Z�ј�a�E.4�4\�cjS
@ݖ�@���TH��^��״�����D'�$��ȡ�u�{}/�r�_y�ՄC�������+Ʌ��*�;�rK�H�����{�f\{���J���? @&w��fV�װ��BNr��b�+1\q����)���K��3	�T�[���0bX3IF7��j��"��j6Q���;�JQ�n�����g��xZ�/���M�m$5H�.C��~�F��2�x�i�F�1rP���(�[i&���+_�0���z��e'P�����6b��s's��o���_�3�A;ʟ�Xy��*هmAw��Vͣnڙ��m��� *רH�<dx� ��Xq���d���l�ޙ)Z���"���b���z��a���[� �u��4o	D���CJ^��R��R=��`���JDg���v����5MJ�7�O[�&1^}�J�3��O-�\Z���8�I�LK����g��ϚQ�
��#��?�	�N��k�> kÊ�.�zw�'�{	y3i�.�9�y��J�ɫ캪�G�?�6)�WJL�W�T��?��6���c��Ϣ\�S��4�K�����+p;G��x�2v��z��3���G�w	�=dK��L^�>��g�-�E�]�Ҝ�i;���a"�"@���~f�H�U�Ñ#�.:���w<޳gwc�s��=@��5�����p��ΒHZ)T_��g�X(qU���&mKD1��An���%��5"�	v���䌠�"��)CYsKT�)��1�|�!k��:�c��k>y��6�C*����}�8�Cn�0� ���3i�x������>�����Cj����0ߊ�.��<���L�;yE!�QHT�t��i�1s*���a�>ř�h��pa�jkC��OVo��Wi���7Ț��3v��\S��T2B���F��W�7
$e������ݬʨ��i^�5������c>��u�cla�|D�P��`���*��[L�	K��U�O|�aU�a$���R�[q@�"��'t���T�x��:Ӳ�G{� "[�鳒����!7	����.i�8<eެ
�FL���$���K���1��2D�����#�k[Zմ.h�=��e�2�\�����जf������["q��Hg�e'=�R]<{���B失��|�db
$Iq �3�K0�XU�u
%�ڊėfX��KQ�tLք��.Ѵ�QS����A�Z�߳�����������$c)�����Z��G]�+L���d�cĢ�x�ڦV�#Mp՘|װ���:�⭠V� (��t\��u�p�>c�}�5�9�v�=��ʮ��_�>1u__���2��R���6�#)�5��� �㦋mQ|.�<i!�g����b!�qZ�7��}��S�5��GQD�	˒��W%�Ar����6���%OG����O{5����#�A��[�~J�:=�����;�=>!m�CЕ��ڴ��ɟ��$/�j������,�:a2�3oy��$�Ǣ[��ŵ���p��=���ͼ���e2)���ر�����g�1�]�;Ə��5�:n�O�Z�H�)]���Z'R���	p�����o�-�q�W�R!0;Q]��P��� B��t�\�)���+����n��&U���Լ�?��"�
6,�U9�TZ�;Pt���E���8�vI���6h�Jn~�;V� �u�H��d�4���P��m�
v�S�f�1R'r�]q�3u3�f3sw��cϞ��g���<EB�<`�:b��i[���E��� &e){;6��z��Awo:bTTb񶝡G.xoro�[@-_�K�[�.0T�c����E$�4^U1N>����?�	��.���~���׮�����J�>��ք
�ʶ�(�m�4^���J!��O����,̦ a�]�h��EF�`P�Ŋ|�I�8��>��xƊ���t����Y�ĝ��`Txݜ����<����%�	!�?�g�4���](V�K�ᅗ�Io������@q��0�-�P	�޵M�����`N��w�:������{�G*�:�Hsd�tٲJ�F,�scS���1��O���w� 	����/���j��g���H�_.�r$�QO� pr4N�^�p@�V�#/7��5�F�b�Оw�Ӹ�L?�x��㦀oKO�\�߄P�Ja��|~�=-�B��\Q�p�$���>����M�{v���R�Ɉj���ü{��[�>3��ҟ�Ӗ��c�N��)�D"�Sx�CS��+5�愕��i�s������ �(p�qEՑ֘Ca�f-�E�SW�K�Y"���V��U�+n�rGT��I�FZ5e�$��ݠ�D�#��b�:1�Ζ��.��9��ž��\`��\qM$�ܙ�H֘�%�}Ԑ�mac�!f���w���w���ݒ�j#��3��Bv��(,%Q7�(�~'�i}p��L�&Hĵq���-A�[]?4K�Y�>��8��x�� S��{ ���9�y�=�]��;rzq��1M����R&|��aot�m,[�:Ti�l/z�ǭ�
�e��;��6�bH]�N�l 3�La�j��I�"cSM]�bR}�B�'���T �A5��t��]�BU��^&T#�v:�6����u)���n�[�/q���ڼ+Ce����}��jj
A���vO2��J�@���F|��G����i���d����\ �Z�C��Jt�{oms���Y������F��}0���.!�yt�Wɡ���+����[F+N��ϟV'��-��W��񪔼u���~_�|C'74��M$��e1����Q��U�u(��^t'���
`�9�����⌭&s�~�U'�u�9�����F���h�A�����5�"��?<�hn��4�\���o��$���Rk?�?/PI�`��5�Ȏq�����f(�tM�U�V��T��;���@{-?��}�L�])������}��A����OA�'���z@�@K!�t�"�~�+V���6%@��ܴ�U~6j���9�N������'��uvQ�~<�6�D�RWv�y^*5�,m�/U�V6R����{H�Fhp�\��q �X>����XL�6�-�\�(<��_(�QWAe�G��E9=�?��9.�x"��׍G�Ȧ��� ��H䔮��f)�6WL4w�h&z��e��^�� ���n��$��J�����z��q� ����g����/�����s�h(��4z�#��G����k���/��'�=��d�	Y�׏�����/�����i=@}}e�0 ]\�V	���շ��MJVN�:�H��U"�vÊ�#H��U���I�B�P9J<�T��Z�Z���	��2U�@ˋ��#E:,ns����IO/�[�'ʮt�ap@I;��O���Ts���|xR�b��K��&�V�e��%߁g݅��:|=bI��Ѣ���
��7B��@5��R�q�V�j�������+��s5#��e��7A�5���%�-��AA)p�	��f�I,���j���w67�Ǟ��B4��<�H����BT`�}B��/�
��yG�юo��{IHicoz���kz|O��{<�O��v�M*{\����>��I�*�`X��|S_���=���g.�Ыt�4y}~Ie!֞+��>����a��l@���5�h���6FP%��������P"�~���Wj�PND+$%�:�F}�T����F�E�q*�	@�ٕ0]�VЛ�Yk>RT�y̓�Ã5lV�4�]X~Y\]J{|@�,p�6�X�tSb�FuS�B��N�3}��-M�k�mI��	�o�cD����R���_�wq�g�d��/�����8�k^D��!%aJ�)���M����H�|@�9�?���-�eb��ϭ>Y8Ё�2�]�"	�?P��	`[���V�bQL*��1��}r��ց��&r]3;��sp C�!㻬{yCG�cY���y�|�mI{�!�|+��! �8ss�]����J֧�押%�am��^�b�\�g���]�%��S{K&isC��QO�OCV��}�M/���9 p(�;֮��Sk ��Ŝ�P�����c���T�f�z�g��p�?L;Y��_w�f[e�����ƀ�Y����!tvϜ�<:������'�a'a�2[Ѐ�I}�{��я�|è#�|�u�!�c1X��O&!s/ �>:���'�+�Ā��R� 6��1���Z�<6��U�В�s{��rGkrZ�[v����<�o��/�{5�n<Ou�g�f��5{j�T�l/GV1�PK~���説��|s���ְ!I0ۨ�@�J��
q���A`nMp(^���H*_���  b�&�FD_&W�g��J%p�$���6���Vt�K��y׉�*�fE)Y~�|��O@��X�Ѥ���]�'�lW}��:�&�н���(��=�3�QB��T�\��)]5��,��á�a�t��h�-j�����o
3PyGut(9�U]�!pk}
$Q�h6B�Z�v�k����`��0Z(����[��w�%�%�|�Q��y�Q?�Ma8r��]�x�!��n�W�-ΰ��C��np��.�����#�E�A��-��r\H�D�z�f��[��5�f�x�΍<W�4��垓w�W��b�}��|�y����]ߌ�x��I�e�+����Kx+�`�5u�G9b�{k� �ۗ(�F�V��4��,�
2kC��X����b�xEV��������������TS�Rx��d���6��6寲����c�x�+C���/sd�T8�0��TPݦ�
�!ke6����g�U�фRXz-uE�PA�=Ye*�G����(���F����N65Qz.h�S�X�ڦ�@uV�u+X)�3g��n���i��,��+C7�ݾ���e\|�#���~�,�=��5��P��QP�mz}N�Ř(�Ԋ�R��n��=�IQѮ�� �L6���vʘ��������P��0���Y�r�=V���?�ު/�~;bزjB�y��sB�֝ �~M]�����Y_$�y��M��)e[�)J��I��F��㱢��pg��%M��D��|���\l���c��g)�>T�!>BͰ�x���t<�+�=�I�����x>��0��Ƿt��z��b
R����.��,�Ue6<Fɂm̨!�M)�EO��rA㊷�v���O��v*����Ե�9� �v��85���#R�KL�Ҹ���5�����ClQ���rO���)�
5	�&{��_Q`���<;Z��F�kx;W��Ѣ��u�շ���)J�����b~��>�%-��d��^}O3��+�y�]�H�`Q�ry�؞��0�}����8�w����5Ә-��צ��%Gn��7 �\�ɛ�!��V��oùa� ��737��nP3��+r��C����Ό���]��:r�j4SEo�Ȫf#��!�x_�ic=:{�!UV������2��>h}F�0��gj�30��s�PN�K3�����y��x��gV�:D�>��.���*K��ʃw̜kR��HY���l�~!4��]%�q����<�W٣X�(��g�������5�+��<5G)�k*惱̱}�!��i���&��3x��C3Z!���4Cn�,.�J��s)%��Z/&�R�0Z�.|F��
�[O��uíy���v�^ȡ���R':^b7=�3f�ƿ[͋�v�>���˟#���N�l%+\�Ȯ�n]4HUs��&�w�&�Ϡ�"�tϬ���{�:�<-���F*�y�D{�
F�˧�Դ�n mq��b3������9�ąw=ޜ�Z�zo��Y�}-&OU��xk��b����x��J�@���?%�������*P� l���bG��/�X]С4�b�U�2$�K�o#���T:J��t�9�쉤2�P�s�k.�k����ڟ��Hzܖ8#s��'@��Պ6��h7Hbl�q�/���Y�K��)�������_)�V�a!�@�7'�o[����Pŷ�czmf��W�C�nU�|�[\?�.�y8�~
��HL�<�*�y��mV]#�����ʾ��]J��Nt��YWU����������O��xU�u1hg~0�70�GY�mɶ�H��fh;^�A�Nc�'��>(;p�W��[�B�qB�k�Z|P.t!\?2	�������I؇=�p��k��oC��f*E��^5��O��f� �ϧ������^��~rGfXә}z��wOs�R�
T��D�
����}X��(�&<�@��v����I�� 6xt���r���a�w�{w0Z���i���V�XxG��"x�Y�Nz��6�[�L�������lsm�,UH�@�15~�"�������5�;	��oi�z��aA�;�	>��8:��ð7/���5�(�U���K�^Z�� �H�=|��O��gZiz�2]#ԙ����F��=)6A5 ��=i�I_J��$8���zR�xX�����R�1K�`m}l�U�Jd�x�b߅ir����	�tu.I�LT@I��`���C��{�7��"�c]�W���;��H�ZK�}��L��ֶ�K� m�Z�}�hH�C]\C6��`.�!@k��(�1���|X�˔z�~ �k�#�+ΣO_�s`b'��x���	f�I�/�g���$y�4�˓���s�z)��}��^�jC!��c���F�=���O�݌��� �xl��4�ko����CK]�u�����W��3�������n�+l~�]n����J�1
p�=�hXq�O���8Oe�Vw��EJrL���"?��[��A�����X(,{�mA8�=S�Ţ���Un��8Vn������޶7�Ai��$Q99����4�,��k��!�M���0���g�P���(�\�=ju�(���l�f����_&�'��n���+k����Ӑ�)�0`�\��X�Z�}�=v��]Y�G{`�3˖�5]�(�Rt�>�6���տ�u%������Ii!�=Z$��{F�u���?/��b(_�ʎ��N���\�J�����{Q�UT�djt���%ita6��8%���������"�4EtM豈"�	�#�`V�[�UDƋ((������d�7�H�_d��pb��U7Nܑl��ܺk<S�D�i�g�`ӧ����P��}���,ҵv�@����;o81�	���ȑr(q�9r�n�fA�����s�nJ�Aq2��'Ie���rkz���Y���׃6��9q�(�0��>uB(���~+0�#ٽ.[��>�Bc�{k,�<�X0O��M�i}�?��7�@̱��F���]?8&���%��!�w�˞��o�Oo�%���z�� šWٞ�OZZvE�pa��A��g����M�_�zQ5���HGH��Th�.c�kn����X�V"1��%� ��}���>6�g��'��a�-�)h������h+��C�>xZ��S��F_�"p&��j�t��_���|��ܥr
q�����������F�A/�/@a]��Ye�@3�?\^+��%��/v�����0����7��oZ�`��Lƶn�W���(J�@hP��Uv]�u�1>Z � �`oQ��]���q�������s��F4�$���(�:�YG���vpHp�JQ�1��@6��:�Q��b�&ؘ���md�W�&T{�f�N�<�C�����)QOw��`,�n
T�:c?���l���3��=����Qͅ+r���na ��U\7t�LFI� \�{j?��8򦣜"�~�����Q�51!Eg�8L�l� `#����75�9����*a�����$��2������TU���)�⑬���n�X(��Vί��}��E�i�v� �A��'��
�d�Zc%�����%�;gA�������Z���g�ua4��{D%�~V�ǃ���ܻ�[ۅ�SֈBC�D��X��+�r�Vr���� `�x��KA�n��řҸ]��_8�C�(3������� ���0	*g��HZmZ�o�L�|&I�a��������4[ȘF5�ŇS8���dcn���L�pU��O�s���s���&�G1Juey��Z9��������%g�zoj�1��(bN;�~���	�&-��0ru�����^1�U� �9��p�}{w�_���a�w{n� ��'d_�Xt�C�mɎҫ��(Df�:�FC����PtX���u�6�y�Q�f7��N ��PD�������<X9>ڒ!o���$������(yM�&G�%�ww]L�R/��CGi�����QŘ�kU[J�m�!>��a��3�.��_�! iF�N�8;�y�Bb�a�G�u=�a��?��-�'�V5Ϧȝ&B��)%���tA[�/h�X�(��Ƹ� ����� ��ھ��r,�LZ��A�H���?���Q����:U�ۣ�]U�ÞŲ
Cʉ�b���3���4�RL['{LlwF���r1�ď{�}�CF>����j�4W�GWS��¾)�>�j��]��OTޒ�l��P���cT"�M�5Y�ʍ(�4��sL!r*��lz��	��2:��v�G�=p���bw��C��d�F�mN��� %6%wR:h���Tw�2�H���j���v ���(Q��Q�K;���_ҿ���Ft��}ƃ)8�漢��uԑ�/��Z�,�{���=c��U,e�s��N��`�Y��v����n�@��!s���˱i���L��>��W i�ƥ�w������z��w
�y$�2�X�q��S��'��Ou���$V-#&�&�IT�rƤ�'ȇ�Br��f	~
�&��#H���e���[؆���`���\B~��G|���X_����oayg�̼�
��pS3��0_��%�
B���bN�U���k��"�6?-o���|/�Y�&-YP�0��g�R���G2	<_k<4F�¬3èjU$tx�^��@-@Ԭ��	�,L���*"D��F��������T��ܪ�P���Li���C��>D�FC3�Z"��*R��W�U���� �X]�zy\��ɽ̞=��G1-�c�m��RO%��g���Ьo�<�r�,nAݬɨ��=�	�m�J��T��qn�����#�^Mc|��Z��֎��Po��:�rg�ɇ����It V�����
�jW`�o�Շw�Ƅn����CXW�{�m�Oۚ���y3Xil��9�}o���ˠ�H�@/�tM�Z��W��7x,���v0�_��}�xY�I@��?�U�e}��E�݄ؗOaPO�i|�p�r*Q��B��|��Um�*��:����D�t]�Pg�i.n��?�{	�OS�6���B�P]��4u �����PUe�����3;��;��D�a�F�;���S�Z��+�PR�JB���J����pxn�B������f��ԉ�'�:LM��q��U�ӣ�o�4�D��Uvy�nޱ�d�|�C�.Uj	�@+h7����ī�_	P��S�J� Lv�G_���*������j�ݳ�%���څ\�E.l_|���l�C������ؠKAw�;�}�h��%���9�n\\NJSn���@R��pұ"���y{(}����1C�[�L���TQ:�6�Yc���ٿeo���U��]���.��\�����E^W�xM9������MLj�F_��r����P����z!L?RvUd��f5��%$��:6o���=ü��R~�ư8N�Y�oV\��0l��T�n�.۴�LBc�	�=K�|"L�:�X��C�2(����Uʬ0\e�=ۙ�a+�JL�������+��	�O��1��7���5�S{�p)����Dq��e���I �?�>���L>eVsc���9n�h�����w��ų��Bih��#%HHR��;���u���Ε��8� ��(9T���\
��D����d��ħ�b�C���6�Bjb&��xQf�j�'�|�䜿	҅IM,�5��|9g���\&�Y ��4�:�g$L����=A�rG7��I�.��Щ)�C������硛t> �Z$g�H�V���p���O�~�L����oM�²xr27������� ���	�Ր�gM���YA�j��n-��
��~a��5.��5j���ڗ Xp��Y�S��-�q�w�P/�?�^C�����l�\��ל�>�K� �����E���CBAR��a�f�X7��ȅ��<2M� �`;�5u�#M�z'6�������@��j��*�WU�$��dC)^�F�����K��j�;+�49^�'�Y5I~і(_�y]�0�n�O�6H�$����|M<�k4Y���#$��a��v�=�����z6�I4:��|��3�9�҅-���g�^�b�>C��ηe��	N�����gk`�����VI���������(��~����Pxe��n$Rf��JSFU7�,n���&����k5�@:إv�^�p��<�%D{)4j��"�P]��E�f�X�l�����'%����O
���Ej��9�%�m_��4����b��F�]����Pf��Z����=�ZA��8Y萍`��7�6{4�lZ�2W }6�N�ۃ,Zd�Q���sh0�vU��C0�&�_,�we�/T0Q�����}z�qJ�����R�fI_�gQ��?Z~21[����fT����j�����A��X�\F�HM֩����J�7<��zUl���ޖ�|�����\���h"�&��T�_o�|eR��c���;P���"�Pw_J��x�m�%���xۏ3���$�vNg�x�&�ȉ���ƛUcy�%~�Oو��{�����{ Di
�n��s| .��y��R�  }
�gV�]`O�=ύ��5��"�2���!�1fmذ>d+��$�����;���t����u��3����u7x��G#�A��b{��]�/��l�U3R�|̺�ng��S�
_��g���n�?���ؾ�X·�
��Μ��m��ej���yT���k�ĘC��q�;�j�c*����x����,�Z� �Om`�)ͧbq�Ǥ:_��� ��������R�G��7���z�Y|oXFe�#KZs�I'*��8�������^��\�]~������71P�!6d�&�_!���t�9�ݍ�+��uӘ��U'%��.���k,U��Ɇ���B���"Sfq��o�S�!�1FI�d�/�}�����ws��,�|���4���Z�"7����~^�GY���#��{�F^�;���x{`�� �'	 E�|K�v!0���1}�t�<f�ٚsi�ʯ�e{�P�A��5��������Y�$�|6���]�G���P�9?F���zh�;��\����A�-.�8U���X	B�ɡ����,���m�.Z%�ȟ��:�~�Ӷ�-7�(�����U��8R�R�Ĥ���g�����b٭�?T�-�Ml�.y�Gk���m�Y,�I"���p�;l?�/�I�r����5����Gǚ��=6�궧��u�����'�o���,xbN�|�G��.n�\���㑣\�{��$�Çe$z�t ,Ք;N��E�4Z�O"^��|VK�]a,��ڽ�f�ʫ��,)��6��`�e��E^ghܢ˾	ט6mbj�oE�;K	f_��ɍ���(b�q��[7�6[b�X��.B�J%�����5�Ar�$z�C�XWC�w:��
8n���o
n��}88��{�m(Fg���4��Ռ��?�މB[�}�]'�E���䇰{��g�"OkN�2�������ݞ[��qR��B�x$&|��5 �F~��}��bd�w�|`#P����nT�&��a�F���f�����~sz�vxqK��ĦSaɅV$�5H�P��"�:��?� ,��h�����]�i�O����T�ޓ���c �=�����5grO���xc]�%.�1g��z潅�������	���z�}�C {艩�M���R���I��O�O��w�Gׄe�@^~9C�,F���,u�V���b.Kg�������x��T�<�ݖ#臎*�XC\����Ȓ�O����Y	�dw�/��GOȘ
Y�<k�aq�"Ò96��Z�3�;!>8��R��<dx�)�Y^��<��𯝿8�G�ŕ��`�D��蘊�8q娸A��폪g���F��Ѡ�z�MKW�΂��`d�9��d;8�6���1�=������@ߜ��
�g�2���\�>Iv�4gjyZ��:���7KM�`r�E�O������?µ�r�����Ӳ�>�i�����Mn��nS�ᩓ{"�v�|�驲EA�l�[I�ߣ�x,=	h�����}��?�$bzr�L�ش1I;T�~�gp�
ky���T��H�w�@��1���%�u2��XH��5�=�T�S	�ΟJ_&@�<��VS�m��4`>��؇:���s;����mb
}=���5������I��C����ٓ|���&n][*b~�����AHCt�b��
��ɥ�����Y:�&��8ښ�^��#�=j+7�����D/�\l:UN����vI�9���Rϸ��|��8�jV��-�Z��ܺZ����uW�gW���2}w���G�������o�\[�,U��S��ti�rBj~Lj�z�?z����;8�+TH>/{8ߙ}8t4��
E�h����@N����0tv��d��!��,�	Z�C��m�d�@�x1���TS�ֻZ�`� 6{JK��zD��;;x㘵��_�n`�8򫏰T��F�c�X�v���sL~�ϯN54�h�)=���\eq���p@$;$'@槇z�����s�E��;T+k��N<G`�(@j���m�D�5-a(��p{��o,��#��{�՚@��K����|���f�+i�����j�ü�q� �(���i�zk�푺<�.�p����Xo;c����/\}{9Xl�Z�g��YI�M������rt�}��"���k��5�ȝ�SNU�2���Ρ���������q�5:@k~���d��4�m������S.?_ﱔI��	v��=L��T���Qq%i@P �<�H�4���=�g�V�q�H���6��w�3�����%ż��;BSj�l�+��a�Y~���%(6���B}{��I��E.�#E�ʗV�F����2�T	�LXd:	���<��\�t����ZB�x"h��r%�VG�3ʲ���]t�Ϟ������R�-0$��3[f�+ ���MP),\�O����Pm�nɁIGm�Q�,T��}�����7+*D��5�O�*h�d�5[	0��� (^�^�y~�Zg쥓��ع��o��e�T1��:����,iЩ���̿\TNQ��[�yc��z�+.����vGT�p�1&�;�����?���l��C��f��������s��m�� ��*��O�D3�R,�j��o+GW�O�`}QY�ǻ؈�L^�D���k�轔
Ӄ�o������/���^�����\K�T��"o5�,4.e�G�i�А�al�C��y��
D4v�� ��sJ�d�E��O��_:�ˣ_������n�j2z���Qm7�Z���x	j�i��-\KEa2�H�9� |���b����eCb��U���k��r�v@��U�9��,?C!r�ǌ�2��D��X���y� ��n�\��M�G^.f3�[:7�0�����澑57A�Q�}�¨�(����9D���_+�5T(�x��O�m:�oz�0a�j!�<�+U���jB�`����NOL� ��I>�������%�Y*�bY6����+��L����
J��]��xM�Q�����E'b���j6;��)�< ��>���x|n�,�{ԊI��'H�_�˥#Jb���J,�KK{�ܳ�f�kQD۲��+�kB�~&t�W�N�d�I�փ��V����攢ä�*{kq�
����c�f�c��((}$�S��@J��� �زK�}����&(;����R;x��o�9�Ê7���N�i��iH6m��7Z��N8�of-��K?i]KMR���J���Q�\��2S6>�!�O( (����op�nZ?���`���,%�_R��J��q�R��sE������	MK}�Ew��s��ҩ�f��D��;��;Lo~�_<��>	W&}��_�&|�Rٗ�G���y=״�.
�K��}���:���h̪���*�X.��|�{/kb��p:���[�bvQ*i�_��z����Ƥ;�ü���ͦQ%O�!��+���]�%g�m�P�C�M���r_�!O�:@s�*�<�d!u.C�)�ĳ1_`[x�v��d2�W��¬RG��@��h�ӄ��U�%5���:�b��Ȋ!��l��uh��˖OЌ�]��#��)�d?B��/���M&��`���yq`~���_�J��],73���a|���)�Zg<����>���?g���n����s�����G�[��`\HvVUIQ�#
��ʩ���	��A�iUE�l��Aa@�S���M��g���Wl�g��"��x�����q�� b��)6ͧF�B�q�h�9��_�o�勠%�!���AD�T�r��X��Y�C��Oa������4�%a*D�~��jW�9y/�-7:�mS'��멈;k�~i� ���7��[ZB�GV��/���O���I�Ζ��7�d5t��WSB:�����	E`"R�e�5r�iE������&�M�|�r2D����f��츉�0:jP��+���
����zS%��a"�%��ȃ"�9�G]���f���&���`��|^�hd����Ko�P��z��Зl|��+cAꁰ]�'�E���QPL�F�/R �0Z����A�?�I���|�lG��QCnhA���}�pt�w���-�.�5w0
f���LM
�=�p!6��2d`OhQ��>��x��80]f�y9V9R��϶e`�X�^D&��B�V�n>y ��U=y�f��B��H �v��i.LR�$t�Tp�/�%,fk���M2���@B��B������ �[OR,.��
�mM9�Dn�ƒxI��Q�ER�
�/$�~�ߪ�L�d*���!_ߗ�������Pg���XG���4�0�v�w�������*;z���{�Q:L�Z[��@6�[��۞���JfJG-���ǉ\ ����~^���Qn��~3YX�A�Z/��%~��A:-�h�`�����Yhec�6�f��;I���H(Z~~,��U����+�ȿn:S҉̓<Mw��ъL�u%��W�r�4gB�Q��]����U�0�7�5�P�I��B�^�/r��=��{\����^q
�D,�t���G(��.��SE[�RT͛
�/�0`�1��w�dY'��N��@��3ی^R�#٭����O����mG�u5wSz�sl�����y�i��p���G�!gٝ_�8G�ύg�̬F��q7)��dU{�5�Yo_ɢ�i��MR�h����[R��	d�uM)����fuPQO�cK��ၗ(�)x�Zd�J���xธ�YE���S<b�@3}��㮽ɫ�n߳H��D���)���V��+��^�����I%�3�"G��3�J�&��Z(k��Lq��/�g8Ee)����)B�����8T��Cg�$d��7��#��8��_�ׯ�C�ӥMgǧtL=�2���:�>-i�S�n�I��1�d���,9�K��)?
�����ō�,qE�Z�}GX���s�P�fN|�B}�xw���7t 0��|T�}$�]
0 ?�9_�̒�,�!�+w���E������x�8�*���0�GES�C���w�cԍf�m�_���×������L91(Ge��`0�4�S�������!뚔tਨc�R�B�.y�Z�j��߉zN��u��	+3�FB)��A:x8�pbʈ	��M��֔�I�)����<���k��$�O�Ҷ�˽C�� ����P喾8օHj*.G�0H��tAy1Q�a��q�2�~�įX���8X�OQѨ}b~%� ���,r%L�9l��WZ��~�����H�od�Iaٯ�C�I�0�6���k��jY�\S�2���}��ڛ�{y��ᆑ$_}Q]�h�}g'U9��H7��ܬ���O��O&a����Wr����
(Aw?~:���ϻ���V���D)\�ud��È�Y0_��-]�>z?b����){��ҖL�i�� p�(�^�g����/�0#�e}➠���~� ]!�?�̠�y	F�HE��5ʼ���.��A�ҕi$�0��,J�Kj[8Uz{�1�_W�_7���o;XU��TB:j�A \WH�h���+ܩv��{�l�b���R���s=�G��S��h"g�(��e�!Z����dɳ���pͲ�Y�����3���_?�6��@v^�_�)���2J,Ŝil�\%�	��&�ΡwѮ�!�ޔi�0���13�1V��^Kd(�� �M��K($f�:�q�.�0O�6�~8���l�u)U�B5L���Ja]��;��P�6	=�㣃H�J��h5���#�j��/���D;t��P������ldTU�� E��*�[
��E+�|���"�/<ŕr\�EB�� �����%��$��9��	�*VX������6[ v�d��"(:�Pm�ɷ��?	��K��|��YH~ƞ�3�P�+�n���*{f�L��pT3]�>ޑ0ӳ��E!p��l�i�#�jH�}z5RX��w��� S��7M��H�c1I̊e�%"�	�����!l.�N4#�z�m�7
]v<��\=?�8-����m�4}�z]g3i$5/t����O���^�H|] ��{��E#=>{|��z��`Y��/�{*���f>"�,�&QY�#��u���f�gF�q� .(�B����j����r��� 1����B��h"[Ɠ����vA�w)P�H�Òq�c�GU�(Y���aH]�K^jn�'CũFң�F�&3��%�g�Qן�*����+6��Ċ��
�ֽ\��ś���}�{)�����'�=?z��<*Y���1����J�`� ���@�5
�U�?�T�	)��V��Lu��W�H���aћ�$���eZ�m`��B����Gھ��'�R��]^QQ$�׳��r�4�[
�z��8�A!���~���ҝ-�Bxزr��huym��z�B"��,�yPʛɐ���>C���K~(�^F���ݦ���3Ch�御�7�����5���]��ާ�ge��_"��MM�ۭ����g�#�V%�+�f��R���J l�CJ�P����,?Z�7�Ȥ��m�D"����J:�Yt�����}��n�`T����C�k�1E���JN�V6ΔB%%�� �)��YB�9�������0Xa޿�WϤ��v� �fB8�S�|�4'!8��Ç�M������!T`��<o�+��H�CU��!��s�*`%3	&�R�3�-r;Bs���&u����q&��J��;�~M�y_�*#Dn���v��r�O/W�U<�4X/��&[$��^�1���Zj2��]��4��K�]��p���r��?�8ص>��^��>��?m�Y�%�����UZ�yK�ȳ�IlG��z,�6^� H��S�0}�[R	̐�I�1�i�����p*�U���2���fˌ�k-�|�՗�z=g�(F����A�o�v7��e�1���׋K���T8Qv�����K�� B�������7%1���2 6���l��=��"Α�� ��J`��b!���rzLT�1���c油��9�d�.�S���f�OO���>{>�m�{��4!s{��Ig��P� }�&�#�[�y�"���>�We��7��A���l3o �?X�LaH���7��}ّ�#��*�:�U:�q��C8��g���	��7gP��a�p���c��QZ������?NCS����>�b���їI��sNB1W�.�[�U��±T�J#�]ͧ��ǫ@����<���JW���a`�x�މc[��D/d�ĕ�&���d��ֺ%���D*7���^�dʩt���'�K=���s\��S�[KYI���T�w��dE3z�e�!o�����D�-~!�� �؛��KM������翶~
�qAu�=.<��:��R��jL˴SS��A����{r��p���T�X��U���C�E���E�4מ���6d	����?T�5�w*\�y�����Ϳ���ˤ�Ca^A#����N0r�y!��1��&�z��ۑ)�Z�)ߔ��*�˖}N썒����K"0<D�	M��ϜbZ|c�dC�j���T�_���J�s��t/�|*��C��LtC?+y\�5�Y��@�O-�X�b����J�I�/��P��~5/��7�?�l%�+p����oZޔ tԈ�Ŷ�X#L-ⲣ���{Ѳ���Y��/᭕P�i<*�Ղ2z������8��Ɵ�l<��W�#{/��ަ�u@�|�}��W���JdՆ\�d�� ��������0ǯtE�+Y۷�ru͜
�i�b.�����+#��� 5�\���eu�u�a���~\O��	jg�{zl9-*��<�s#���J1Y�
�nƣ�&T'�IIf]}��X�s̉j�F�GD�	���_pO@UP���I���K�Rl�w�����8�x��Z3&Y��q����W��-tG5�P'E��L+'ԝg����b��m0D�}<)70(��7�#7�Y:V���Zy|�l��%�v�9�;��[O�Wd�A
<8p�lHBI7���5�b6=��X�o|��g��<ܣpO�	���~�V�1����^!�Wg��q�a��:!a��Q	��,��v%�m�H��k���K�"܎�68ś���K8ֺ�{�����1}h���<e��A�n��&�ֈ�a����u��ñ�U��ҷF�2P1�Ȁ��.���A��ǎ�><����-vU���������;�q[j�'O��)�������|�Q�:�[3r�P�m���[X�Ȱ48���O�S%S�)��{J�:r�w/Gn�j���3J�V� �T�q"i]2�g��0W�}me�s�gnS���/�cJC�Ͱ`�d���fB��E-iT,
 ?'��A!+���x/��bF�&q���>�-  �`cE��Ҭ��:X��]t������8���ɽ�1\�����k@fS�Fm{��so*�ks�"v�δ{Ab3����t� �m���R㚝�KOs�S� �3&#09gk W���g 4R���]����]��v�e��o /��Tb�Ui7�lSk��"��Z��~Y����q�Dd�yN:�w�$z :*���߼����,y��DЃa��W�7���|N
e�A��Ţ�.
M��L6����2�����u���x4�� �6�"뷵rI�'�\��왇dŦ.�ۏ�՗*ճ���
���e|$�
��A�R�I^x�w����
�o��t�(���Q��i���F��Ў;�"��ѣ��[��cl�3�' ��=o&4�5��d�}2I Nu��(��]U��>[��WLG���۝�T3� �#���/W�G8��M�"Pf�[���]ߏ��4u��!ؾ\��7�z��c���;ͩ����̠�E(�W'NQ�Q��#zRYV^Ͽɭ�'�F_���D�a2�y�@'[��}b��p�F�"������~Pɚ��?�G�W ���Rl�;���*:�|�Yy9.�(1�e�e <�PL�E����{w�g!0,��>�7lMT�<�-}�zo�E
�����>�n���(-�UҔ7ߢ�cn�rzY�"%@��Hґ�1/���0�A�#�\'kG=���;Xr�>�#�Q\�'�8�~��L�"��'�����ͧ�꼐�~�`�r"?OF~k���$�?��4��h��8�������&��t��giV���������o��ﶄr����VY(Ϩ7-�Q��l)�ry��K��'���l�f����;��3�I��qF�;��!{�/)6iV��@ϡ�07������\�ƂN.�����n�)pאַ���PG\[*�@��w���=��!��Pԙ��L6{�[/-!o����?�۹f�M���f�I�]$rwVH�'��Bv�G��'�T�<�W�T,���>��S�-�iZ��Q�B�B����!�Y��e(��8�W������S(�]��؛)͏����A)�Fߨ�����������-P��"�O��m�[y��^�+�Ѷix?����(�ܠ�U^ZK/ַ ��2����o�j#��f��ԙR���jf�Q����0���}L�����,ó��{�?~��C�߱H��H`O��#~u��~PW���\~�#�1��W`���p�%��Ev{�М�'�	�����|���i��7����Q��z�� ��f��ml���ȼ��iZ�t�7cn�őh1�Ha�1�dp'�-eyP�Ѽ��F����%�.L�f����4 F�
��f���N�/�KN��2�s>ofa.(��H�_5Ҭ<	�bK��w�3�P�+������j�Ϊ"S��F#�U��ضL��w���r$j;9�bC@l�+���C��m��R�(m�+���|�7�V�@�B�/'^O�{�bd\�w�Է�����up�y��!?���H����:mPq��ơ�x�]�n��)��6�g���t�������OE���6h��?�e����O�i�W���7.����Y;_�����rM�S=l�֎}Nq�jV��tz���t�峿����de_h�`�
�l�Ne��el �ʊI�����Q���C�j�+�wc+u����Wb�+��T�*C���!������o�;'ioX����F[k�4B�v6�.��l$�F+����`z�iA�u���GW⚠��^Ἒ����,��Бw�~&���E.L�h?̹KE�	�\lB����m�:��e��dO�Z(�")�Y4x"T�!�~�E��O?�ζ�+V� m��Y�
p6����g&Y�B� �y
^�j酿q
t*a7�=6�����y|�^���G�����Li����� 20���7�L�L�/�y�%��_٫[��ʯŕ�ؓ^�g9��X���N��
Q<�f��B����e]�k��$�<u$�
�a���fi)ME'Sv�T�ج����#��b"���ʫP���sH22���1`��x�YF��a���睇�C��6���V[�P������eT4�����<_���l#|���_�������{�[4Z��>��޸O�@�� �|ծq��Jg��ԟ�v�Fg3/p�7vG\p���h�Vv�����(,@~��ZM�=<?Z�%Afok9�p�Z^��
Q�z�%]�yCq��T:'��V_�G�5!|6���s�f���q�f' �)3ؾ����}3��z��� =y�g�sY8H�a�G��|�#��l��d��|c�6��O��D�/c��z�:+�伄b����V�`*:7K�-m6�kj���\�[���b���ʻ���@�����s.޵���ݦ��Ѕ����,�X�TaJG��_�\E��=����oA�9�
�-?���'��v��6����c�`Ҽ	P ��9L�z9�g���CW�.3x9�x��Ј?�3	�\Ɛ�k[y��p�����s���INh�PH�+�0�C7)���Ju�j��_��y-�Qe��	�<�����ב�^ۭwDk��������o��˞;8Q�����^��7~)�����X�����C�s��/�sY��x�S�'�t�ǖ��T����M���J�n�S�Mr#q�D�[s#@����x���4��Ѕ�K<�Zw�"4�]�S�olK� [�⨑_r3�=k��4�؀`�4��`N��@�)~���z�[U3���
�D�iHge8s8�ޝ��_$&��c��8Ȓ!L{��JW����D ��l�7FI�c��m�p��������;j:U|:U]l��Ȧ�Q�pk-j�Z��_��}�?�R�edV�%��;���f�Ӱ� � #=� ��{�u�0�T�S�#	4��OF XE�FlYq�$��L\��#��s�y��I�I����Um)p�I�_H�K��W��{�L��q2�V�u��� �תm|�$y��au��[!��'o-t-.��g
�tAA��=�/��,yr9d &�_����ZZ�(d맀�-Y����a��8S��5%�(W�k�E��2!��6�$q��g���УH�	 �mKk,	QzN$cB��ů.��wd�����@5�CNd�:Y���N*�B�V���Ԋ��3��]��&�M!/(��	q�;c1�v5v�lwӗ/�� 6�ݱv��4�Ksb��#�����T_������W�y���C�� nF����A�G��y��8]і�=��+���c�r<ch��x� �[t�X~+y���
�@;�i�r���ɓ`�۫'��ܳˇB�����׭@�$�S�]��~Y��UX�Ĩt��L��\�������r��(OӦo9mkCs��/F��޳�U��1���N�cJl��R�!��ɗ�x�t��!�,�W�I#�T��l}+���BĄ�o�;�����{tyR�뢬��h>�>�0=�,N�+��lҪ�^� ���ux��2X�<v��C-q(%f��#�t���$K��JĿ�EM�+'���E�CS�).�n8D	P�oD�QAsf�i�NN^��u���<Z���wJ�;=�0�F$��>U�\6��/Y�\�O�yߩ�VW~j�reS�iB�� �6��6IdpPZ�%�I����Df~�k��?]j�<Q,B�iQ�`���(0�
�H>q�3^k��q<\���5�7�i�б�v8Pz0Y㙑�~^Ȩ+.8!p��n�db|6��q[T�A�LGs[�(���=�4��ݙ��47$�`���!f6������+�~���]0�$/"�#��P`����K�xDEΧ#}��!�����$'��x�{��(sf����{[�����L���+G͈�'�M�մT�W3�5��2t�*��W&�ɪ�0VWe s������*�ݔH�h��2G,)�A��Ӝ�v��%x�E¶���}�N�Z��S ��3� b1OsQj���{_|��������Q���z����+�����I�
�=�I��f_��i�FUt�iY%���1��K:������H�~[�a�e�X֔��"�^�wx&F��*���IY�b�I2߯-�������!ߗ뎖Uj��|Cal�^T�R�^��h��%�'a����Id,ep��]��!Ln��`}7.�]�u+����qY������afLȄր�1ZdTM(iE��z4B\z�A�!"�~Ud���Ǧ'�2�-�b�s��%ZNQ��p��o����'���y1+��z��/]� ����L�7�O����uh�[�r����wk	 ��U� �k��"�H*��37q��?�N^�t�aqq�O��j\C� ��I����@D���
��7�2l��EG8���q`��NV~���]H�)L�閸^4�Q|���o�w�=��3�w�B'���e�;>�����6N��u��^#��rm:{����f=�̐�s�h8Z�A��[��c��#D�Ä7�	R�U]:�<RO�Z���V|X1iv������r(�n� 5P�(����U��c�H�$��Ҥ�(k)ʤ�Y�~Nי�Į���/���mV����q��K���A��/h�U�yG�ŋ��P|��6TH��M��dff�!������v��ЫE�T҉�`�>��t�B~ހ�2�y��6+{L���tִ�J��q����-��m�N�Mv�:Bl������gL*�/i���dE�#����U��w�����ܯ].}�I��@.%�A��4�J�q�e2x��]k�����g����Aąi�$M=Z������|�g���h;��V��p*bY�E�/�G���b<�`����5��m47%�.s�g����:W6?ٌv
 �^/�A.ҕ����d 0ˇ8YA�N
�)7M@,tf��4F����V���e�Uhr*��������Q��IIb��z*�E�5%p��g
����Փk���*�l1�9��I����$������Ujx[��<⫯&}nY_l�)�C���,z�D��i��T[8��߈��'S=io��'�I5�b{_4�����P��-d�8#%���!`��$11m�s"b��I7�`��t��h�W$�g�����Iz$,���wqM$G`Gz�ϳ1�Mi��E8�E�Ki�KI��"�a�Ϫ߂md�kD�zL�]{�,�^����W��XG�Gf�
�`�A=����&-k$A��G��.)F�k메���9=�F�����W�h�q����?��CgJ�d}4.Ȋ��˷�fZoM��;;�?N�s�u�Ʀaq!������?����+���)&m2E�:I���O���Sv*���:.ƺN��j��Җ�?�^u�����Ʉ�9����ge����>J�^������[/�S�ښ�2Y�ͧ�Y�p�t�m�b�t�WUK����*>)VTB@x	��/t����b���é7�#���;¡�j�VD�:)��y��������^���\7e1D����l��������ik���
㗛i����&��5�J��EF�%�EhQ�l�2��N�0�{�h���}3-)N˄��$����;��D�v�ߙ�����$�&l�aGٵp�V&�FwR������_]G��h@��/;�S�.dܖԦ��_��oSɎT��78v��pΑ����Hl����|-��(˨7�n�if�څ`d��i�Z�!�*%F�,�n�Q)�LM:Ei�m�{��l�ѯ-a�L�-e���W������5�&�0C̴��*B<΄�a���c���I<�l��=%b.65����r_3���?�7���-���G�ݔƈ��P�b/��^y��?ahm��B�"�B����D�9rL��H=�x`�������P���r�,L\�����f�nk������e�H�O�/�&��RM���ykr����n!��@��� ���Ѕ{�Ec��Cv���o�<��u݉���4h7ޔ���Tod�$z3��y�`�`?�&�
mʁ/�P�6寮B��L��8�������>�8��J�W_��/g�{�f�xU�g3�MeX��z�ǝ�s�����T�a�L��7��tsi�Rf������5��ԓ
n�ޮU雇�ބݥ�5���X�;��ݸL�1�/�4�r0�C,��џ�)%�2l$��mQ�ŷ������o>�d�v�f��Ί$Z@/�C�����U�/�i���zus_����	8���?j���o�wݶB}%=��n6.��;M��v�!�2a�����^9�"�)�|Bf���y�0�+�gơZ5up�V�s��,k��ۯ�,�N޹X-�%*IQfT��6�5�l����	#�˗���Ghj��m��o�@���D�z� ���{���}��u	(`s��N-�Ө�R���X�� *���|bA*{2��`�mr�g�{>y����$��5���^[�̛��F�$�k�,A��_��}�@�S�)��f˒n)w,zDU���E(q�x��)���j����T�7�������Ik���B�}e6,�U� =OW"�{J��wS�)�2�������Iկ�
�W�l��Kn���_+�K�k6z��و'1�U`,  ��c_�b�\�����]:;��xA����v�vk�d�]I�3�4J�A��W�H�)�`΂�9�r������;�_z�gӓ�G����Ɡ��&fA��i���5j;��UfN��P���s�ήS�Mۇq0�� �l4jc�]��=��S�}��nȚ�^ZZ٩f:�~V7���]	��Hy�Q�w����Ceh�<kx��9Og��X�	��@�DڸQb]� :6+n�����w°N�pd
�P�q����?q�q"��I�"���A6�O�����4��k�>d]Lb���0�8@Qfi��oĐ�h�&ȥ��*�m���*L�V�h'm�CL"F̤�FZ��}H�b�������G㌡p�.X���{+F��nا{���� ���;td�!�>o�������Q;�,��?B3�M�Wwÿg%���NX>:t���}�GS0�����������gZ9^�8�V���e~@���9�6v�;t;�xf�Pu���I�,�ʀ��t%$�Ċ�Y*]�!��f7V�\IE��=}��;��R$Ũ��;�"`�%�ҙ~�>;�t�tE������ۣP$�z)�+�g�����U".* ���n��\A�'ꭞ9�\�ꊔZ���y�l��D��M��j]=��qS�G�풽�-�>X@�g�Pp��<0�J����U}WQ�����:O�^�s_���������%`> �E���e��Eȷv�� �Wդ,?�����)l���1w��@�^v�k�o7nDE�~�G`���t^��ˣ�]��7OK�^��i��b��Z�|to8y
��5 ������m3�|��^�xu�a��n�k�Cs���e�5��������MZ�x'�������F=��@|^�T��Ō��ǀ�h$ZᲙ��ƒ�cW{�FA�R=���L�q�:�}�\����,^�܉�;g����Dt�4n�\tx\.��4�k�?�>���^�ѓ��,7ҋ��֯��ґ2�4�����-��G��!X��khgT,�v�Q��w��%��·�>���-7О�z��o(44������t��J�������b&h�ы���S��w�b#�D��*���b���q����q��N��B~��q4�}�P
��K����z�N���m)�P\7��b��
�aV�������k_��u�%�U2T�m�aR�L|c��s�����f3ܳF���i���}�+J_�+Rn��@*��遜��b���FK��P��q�D�_�0,�P��� T��Ԩ7Q13�	��֌/@��]�P9f�d��G.�����Y���q��?�蝏�,�߷�!��IBbW��߄rB(��b�״,�#Y$�wyo4��[�D=�Ѻ��e2k�_+�3/����DŶK1�Js��w7����{��(n]�,�eWl� ��l[Z��c�[7��sL�"�������H��'��Cd��Lp���h��'����p�$,�P��!2�IWF�_9�x�>�[}�Q�+�����1A'k���~+R�r�Д�}*�o�������*]d '�[��F�e>�$�'p�W&�f���M�X�<7B��vd�O���U�c�#����5��{y[�&�\r-gS=m9:�3;\_3�)�]��/j�;n�;��=R�Vu��u�ҢWg�<+���;�W`��>�p�Ng�6a��]�]a��l�9�	�R�S���eӊ�q�8՘<����VW�?�e�;�"B����"g9s;����=@
�t���Nm����8�<���(���W�Q6�e�r�l�L���kY[�+2wv�g{����A���u7@�em˥~<JѻtT��1q���Ll��xZ9������F�w��	$@kY��2m{@�\� z�6��i�Z�(G�iTaC����5�&��3��~�+@��G�vԣ���,y��f:�iB�z~Y�����jLX=;�vc���"��4���EtSٲ:�>�xF���
��q?��ɧx3,*n�2�Y��roM�hm7�^�CI%�-3
mi����x�-��@G�1�V5t^�2&�NRƭ����b��;��;Y�T�*�!_Y�B"=�;�+/�ó'�A��e,��F�̯E��Y5�. ��xb$��.�M$
���T�ojN�U��W��34snZO*�2p-�t����yF�L$1rF�����K���i/�&�Q
S�\��3j��(U�<��ěA��S����9���^�ZG֟�s+ov�m�ҼV&�<	S�|���V�>}��+P�I����F�(*~�� ��˅�\#	�W&n��4'�@`\Үh �ۀ����|C!�Hy���*�i<d��#9�E^Jq�4°���^R�#��Rf�"��B	�k?�Hq/o�����|�;<kn���MG0YJ�q�N4��b�3�������+n�#���r#<�������+�$,Ki��CB�1
שӠMC� �ٙ� 1�olA��Y|�^d,~����M9(����$�T�2mPd��@�XE���'��O�V�>ĳ��2+���#d
��S�n9��$�BZ�nl�D��B����� ����Lri:�V\�h2�I�zȸ�����镋 ��
��*����qTD�|�������NrK1�wp*��l�y>L����S>�]���@KF�L��У�^�x�;���-�2�rB�3����\��� ��'����+����x1q>�#c��Mξ,g9�Ś7G�9�@�M����e���)�i��Nc������q�O�%�X���:�,u1��E�\Pe���r�<�um�i��(}g�i6R팝2H�d� :��w?*O1A�H���o�c���%]V8�}JB� �����V����6��+I1���"F��t��k�Zx�^rc��oٳB4�wŕ���I&�t��ς��&��1�GI �!R]"�C���e/��T苂�H^h, �Ҙ �_P�K��<F�����s��WF�l!a;f��;[�]7e$��:���9�@qz�� �v�m�U�#���1:U�ϯL%����L��d��Ym�����Tr)eƚm�P������`B4B�;0�D�j��R������V��.Ǝ)~����ݸ��H�`��y�ޘ��e�H�aꡣK�S��C-k�F~q�s�}�U*쮷� y*�$7�<;�WϤ�2;9N]	���� �ŜO���b�����^��*�oI�)��~�ýx���Nm�nқc�w���~�#T-׮���)g�|_{����p߳+$�x�7���&��%�e�xկ۱��M�/]=l���B��_n%t2����ĳh�C�Uz/�DE�U���R G4��e����C9��*��9��UxO�Xmx��oI�������A����e9���}��1��'��@�^W��2�T�5�:��\��!��GS_f9�n\r����-��GX�s�Pt�+R-�l"~w���hk5`~�:5�{��f[�;U9䈨a����Vty��V�"�{9E�;�ʀ��ؑ�%J{�2�):�b[D85j�Y���EvZ�B/3��B��K��5��o`T43��̕#d(vky�n�{R�v��i�.vr�]�\�o��[ a
f���c-<BŜ���"�#)�������ً�"���wBeB;��7A���)ǉ���_0ek�ԾF$)*�4z�#��L�"��	�Hh�m|#��9sХ�I�Y�öM+�A����)�����0�E�C�ja��K؉���2'x1�����ߚ�-:��s��B0B��ӭ����qo�,����%w�33�A��������i�o��3
�����fR�_���n��}7qt�`0à0>Vx�4!]n]��J�I�+�kCL@�w���B��^V5�ݷ	@>�-�:��zc�u3�zO��x��r%;Ӫ>r0x](\�2��UΡz1C�i�!��u��Q�zD��l8���R�[�����]���ʟr�0�mC��v��NuHM�"/���פ�t��a�!	�(��EpOs�6����e� S�H����#S��}���^����T'[F]hn�<(�m��:�g�+�^v��e#�b�M7U���
�V��G��d��%V�~0�>��@cE�R@�ޗy��U�����n@m���q�G:$���cYP��5�ᠰ�em
��Zm�=q�����6�&�O?�m�5�zš�	h����W��S�}�G�OK�F*K���W��`,3�}@mG7b�)(,����y�nV��,��� U��B���\Й��Ҹ�4[X�e�	P��$,X���~��`��R��(	��,&+f�a��&J_6��/�?C@eN�an��Ԇ^�=��d�*�f�H�Lй �g���Yz�np�g'�R�O�V��ӈ�.��Qf�5�ǒ�I%�<w�S��tmmǇq��hd�@D!�I�V���Sv�����xׯu��_��-�v��������baO�U��ΪB5Sa�4�>��r!7�-��Y%y��i�1�C�J����j%OD.��ڴ0X�D��d�++��$I�0pZ6���+]
�kf��1�5��t�O�I�7�֓c �+Wŧ�v���βI�j��i�����~
Bk5bYI�nci:Yz���T���
�1�F����^1��,�&4���Ȳ����%�v�y�����C0�����.���}JJ�������uw?i#=Tܪ�e	��Qo;��z��/h�	c]����<�pd��b�b]]���~u��(�X)�B�,��DA+�~9������3��Zs��t�Lr�4�{ڍ���O���
g��>�=�S�z·u����C�����4�T%J23�ƯjEwk�#��L����]��E;�aݾ��e�D��
��S{�� /i1�tOԬ}=%s�qé��fi���S�� s�:�f��:G��'����W=韁&��7��A����]h�
m�)T3����%�A��"%�H$;j쾝bH�x���lBL�a^~o=��7KEYw8?-g�} �1&��,SG#��Ǚ�|n��F�V�-K.��?�3�=��^�i�C�C���d�����uh�&'�\���Z�_�
QW8U`%��*��A��c����gj�q��t@���:�]_�K�o��4\ë\=��/?B�)�s�r�?��cC���6Qo)hk`���ԏ8��mdtC�D�jOtŜ��6��@=g 1�p�s%�cE{���%�>����Z\4��}�Ƈtt`_ d$:����s�����bd�R�N�#Ӂ���������(,͙=l>[�L=#���@��+@�,���߀�D��J����I�A��+��VYSm�I"��b�ढ�m�
'�ɢ�����bk^��<P������k�]w����"�B	�p��*�ُ��)�AT��(�G���3��n(���a9�ړו�_��f�J�����mX&�/��+ �~z?�������v'�(���s�_��g����f�h�S�zP`�,�\?�j
O"���C��5���#�㢺�<�C���A��s>�aHAa�ɞ�-�$�=�14i$*񟛒��7�ʾ�2
ݵ�mxB=�,U�a���� Y�ᖪ6꜎��BX���**/�f��"9)3{>lY+�8A�7e��n6��Y��!�U�;^fK.☽��ň��vj��	r~'��1-�����Zl?�5Up�Љ�I�D�V����ƽ,����-N�A-m(�>xЀ�U�.R�?F�[nҋ�&��>�e���T�G#HK���E������. �MLp����bD�H��{���N�Y���/�7a�"�&��oB.��7O�5Ϲ�4�Ā-^�p���M��g ��d_�f$�&��(7����O��H��-��D/Ηr����h�l�Em��`����92(^>j�t��w��<l��7����f8�C�-9p9L�d�Gф���Q�[��.����Qe
aUQP�5��a��P$\g��5��*ŵ�1õi`,�2�q�[���<��Pi#d�MF���^�����z� l�f�闯M(��?�LL4�+|p��]_9�a=��%�Dq�VSH�<R���L���`����\>#�����!���Y0
8��S��ai�`�$�UgU�����Jg����ߠ@�♉�u&N�r�'�E��>��W�o�kM��8�@+�؉d���, oN��!�U#���;� �I��9o�wB@��dٻ>�mɗ;~�Zm�I����'P�I����b�H��^�5���F/Ft��& �����`gM�I�̚h�Ճ,����S'�N��c�7�����u ���K؂\=���	f�59��9�tϼ�`���o���{|������״�e61�>aȟ�^?m�K�S�Y�AaNִ�ƶ85Z�cӽ|L���*ߓ.񳧱�*PT�+	Χ��VD��n��<��;�FB���_{
��
1����SK	����,}�#�z"�_���"-��6}�H����v�>e���l�$��@�q~P�V�ڶ���je:@9o�jȗR������%��PO��P�rP�b�ja����:^��T��G�I~��鿅ߗxG���Gc�E~�Z��=����'��z|9�b3(-ܪ��0\��-�<UU��Qh����n�������rϳ	>s�%�@��`�����\��`Q�*������/zɈ����Q�X�fXm"nr ���Ÿ\�k5������7t� ��/�/��m��0��=���љ
�%�P����~��db���G��e�HRa�����`%����='�0�|��-lAq��^«^C��8�(�~�X��8�t�����q���W��8{��U�*� I��Z�<ZiK$yS�[�̐ _��]?�ﺠ5��jo9͚�a�����s�ZD����lQ-�xƇ[ƈ'�����t��~䍾�z�6�}N+�d��u8�ǹ�����9��A2�3�)�u�/&Y�ޝc�L(ӷF�A{HT"2tN��d
��\и
�(�����v X���,�,�Ph�#z�뛍�Vܛ�m�����AmW�A�A�F��=��X�&�X�
��*L�D&���F�5��ydF�yR�`���x�u~�x]��$r�� ��o�5�F�^��Ɯl���G�#�ۺ6�	�}��e`^��I�3�AO��#���:�����r8���4��,�<���N��N����Bs�7�:kҋ���\)�zB��{C��D`�WL[_�4����C��8�r��.��9hJ�+0$�H�#W��UH(���7��� �߀r7�q�ȑ('�q6Z(W߹��S�� HB�&|�/�a_jk�? B��� SNc�	?�>Dlj�� �9<38��a�l�n�=�GF�kb�b����ɠ�y�!�e�F�e�R�OO�)���s�LV�[����%�!��'qF��JV(Im�Q."~X>]�a�~T�k���^���p{φ\^qim]��š� 2��E�!#c����$���8�a�G�R&x�>{�9Ml&�=�r����QTź������7�q��+�T ��i�gj����Y���ޝ��'X�V�ѹZ> �����p׮R�z���sw���n2rV,	�Wlך͙���(�u�wď�+�|^���:c��@��|
����u��Y.;�<�T1{u
�����#\���3S1�'d&�r�.I��qXEw��W�,mA�ݔ��Ǘ��Ώ�1�y�K(�m�$�4�^�q}�|�wl~�e(BbIu���/������"1n�V��?r|�K#;�+��`�͔�J�����皴|�z��[Y�߲��L���Z�7d� �1q�W�_��š�B)Y�H��^�B�����c�ۭ)�~��V�t������8��e�b �U��qz��e|��굶��s*���znh<�l�
QUQ����cҐJ�4,�ai���B����9��p^}�W!>�K;5l�.}1�	�>/����Ǣ��1�d�@V]�Ae����
�.��x�K��,�W*ǁ�.���ס���jl��6��|��/��&7�
'�v��m[��⠜��70u���Մ��2��J�E�d��~i�P�W�������jず" I����P>���2�kew̷j��w:!��s��A�9���|��Y<`�d���Y��ϙ��5v?�Y�_=���u�Z�W���'�*D�`s�Y���]](�K�!~�*�ߑwh�Ƹ#�u�{�_�=�(�k�СF�4�?Mc����=F�Xzݩ;ʣu"��"����
�n:_��c���a"~�o��!���f���<����������"���jPB7���{�YQu�x��=W�l^�� eIgh�mPlX� ��t�ͽ��?cQ�vc�v���������8{`Z\9*L$@[
G�A�щU��ZXfK�.b�ؽ�t�l�y��e��q���휃�#����sUCu�4v��z�����`h��賞eSL5�R��N���~�s��;�����+*����M�̼M�U���m\�n��Ms���MR
/��ҩ�k?��d64;����/��cZ
���Q�^N@���tt��o�@�����E��yz��]��$W�쟤c�;�w@�r��fT�œY[��ςg�������g[2���?�0���(&�|X�r�n���4K�����$w�;��� ^���ǾO����i1N��G.;���/Q;�P���Ud���ɻ����rФ�a�7^�,��Fk��HݭA�QCi"ظ��\��T�8P�Ե�K��ok�|��sܠ�b���!���Z�
�8�Xr�:�7��SY \b�t0��<N�۳aS0W9�u��A��n/�Nky�9��Z�\����jn缃Qb�(���9�7p�`��:"�ܼ���ك�J_9��9�TSh��$�+8�h��/���K�R��]4qh�G�y#� �D�C�k���/���s�'׼�I�)�m��B%�"ܖ*3>�oN�PLV��.�"g�9X�j�����^�6(�L�ڭ��~�`�0T��N����c���i�h��/��}K�6��Xo8rԳ�V�3�whV�S3�z�;��q� 3g�@��24�pWdh�����r�/��sp��Jk�(~p#KC���3��7�Wk*�7���fZ9�!��Og�P����Ո�i\�낤�o	\j#�K�}#��RV7����}>J,#(����v�A��[T8���i���l���\V���!0�^�s��:G	kׁ����#
�E�.չSv�k����@R�h������3��V��j��̺ns,��I���W�5?��' ,�;��4y�˴Ѣp�Pɲ���&����K�u.����:�_E��U�G�5�R�����
�C� X�ݽ�	ۙ�K�?c�{�<ɶ
��d���1s��gy�@�GD���"EE����/�7*��6Z��t�"��BĂ%��\|��[�H�����,Y0佷L�K{_�{S��Gb�9f�˺�V�'�ʃ���2�$N1���\�:���e��s\6�>gu4k�E9�ئ�?�%�1�4'���P��HC����h��O�хg-L?l[Q
k>�Z���PR��lȦ6K'��Į:�$�.)A�l9]�}R����������75؋��l.30�z��*���	@ܱOl�:�<2V�_�lQg~��e�J�=��N����S�&�W�t�\��n����X;	G���9,SCs����]�ǆ��[�)�>[��u��"��.h�aH�*�rԈ�L�
ܭ30�O��=��]T�/&�K�C"�j�zJ����}|����O^��D��J�_�$���W�Ny���?؅����إ��t����n-QV$<	k�{s���R�<���Vp�d�[]����
�x��O��,b�\��f������
0㆘�F�>�鋣p�,*H+�l�B3����c���X�����bOM���\�V�ܚ�m��-n�d�/t�l�fi�;��|��$�E'O�f�������E�Q��15[��W2&�=�ͦEIl,}L#5ɭWw��Z�,�d�w�����d���)��Ճv�ds/�Lv}_�+Yyw< int�g�m!L��A�ƷML*H����^��:k��#��aOC��N��S�A��)Z*g(`݄�W�NB#4ŘP�[����nr���㇊��W�%�ᑃ�QՈ.��xA�L�K�r�h��Ň?���xlN�)�vn�$���>b��x� ,����0���aQp�\��**��"�ر]�|����@�e��,P�H}����]bp���E	A�-������U�Υ����ކϫثh���9g��t6�h�:�TV�:�Τ�;i[�Y�2�A�S�ho���@�5b��Wn)~����A�Jn�̱�=Q�P��LX�������P�����΍2	�zHa3��T>b{c�
xH�pG�TՌW��f*/�Y��E�wY<q��,.�r�I`f�tD��oUz}f�RFI�F�����]3�Ե}�A��Ah�WY�,�F�=����:ɓ��^�+� ��j�z�\�g1C�
ح��귑3}yu�9�z+f��r��xX0jö0��$F�%?�x��m�|xhE����z-���ei�r�R����vq�nx�77��������ZC��f��\�	����j &�l,1��-<ŮS���25Mr|_Y�Q��C�e1T�� ���j�e�����ň�3��,^#v��:ük�A ��<��?-u���v��h�U�����"�^Z$��`�]��8�Ic˵��=�uS��J��YcO�3x��b��Mϧ�0j��7s�AM3P
�<��F���B�2���3���~��C��ɔ=�ͥ�}����EZU�r�^�/]w��-{	�f�zk�O����	�aʘ����IT�L+V���e�\;���z+Xα+�ga?d�@Y4)�V��*X�d��p@�2�2�v1�bu�7���s�0���փ�c.�.5���ݴ �*�Ԣ��ILx��:�SUSm`TX dv>�?}����Gv��R��o
M�3��Ys��?FV��|��-2�z�-J��aG�I�xW���6 o�Rd�]{'��nxA��g�O���x�:�=(߉7ۦ9�m�(���$�%�6@JuQ��I�ƃ�w�����!���V�������Z��a�<��AZ��t,����_^�iD=�<�a�r=H��0��Z�K/�7��+6i��{����j�{�mz�;��c!�ƍKa���M瞎׀u|�3RX@�%4�瞥j�"fA�;�lG�#����#6à��z��t�$��Տ	�^UO�B� 20�x�N�&��v���p�;�(ͩ�ט{5�i�e��T�����zu��űz�^�vaېY )�a�����\��}��ekỵ$5��l�� 9�̳�S����CW<O"K�|�I���$�can��z�8D�T�6��A���D#�O�jG���?��0x+}�<?���{�ϔ����t����qM��N��]�8aW.�-:����v��k��0�{�Z���l�)/����x2��,qQ>�(w���ս��K=.����7}	4�U t�l�H�>�q<;�m�tq���!�j����h)���b��bş� O�h� Bz�M��S�B�O�>&�mu��78��z��i7�~��A���D��OM�*�T����4���Ϧ�ڑ8�	 ���ּ�. Y8�~�t"(Q���53�8:�(�݅�c��������6'ͽξVUT�X��Y����?|��z�}a�i��[}c�F(��6ֳ�����[���}��h�|5�*��|��x.9B<k4��c/�Xpt2J�^�����L�V��WZ�뙪�C��|`�/�f���<���}g�R�;r�������=�����t:��lm�A{�\�	Gfd3{-&E�9���+_���©O�96�8�ۥ����g��~1�Ն�t���T���Y
d�0X`�&$�)	�ÓU䲝FO]0���ǖݺ�ph��M����S�-&B�]FsKd�ڪ��^�rS�b��0>���>�����ǻ�S�3iGFs�S�HD�鲫ql��}�Px�N��e��e%AGV-Y�7�0�~�a�r�F��V�'JHv�0d�k#Ond?�Q|���z �-)d$�E������/<�]�	qGy F$��J�g469$�%u;�Եh#��
��a���J�X�ض`�qr�d"��KuA�����]&O�D���F�
���ms���҉^�S�ז��TP}a?���t� B1��)W�\�S��������Ww}�Ś%��F���foK���#|�c���ɝ>�b+x�o� ���g�tjy�n"ZL-��q��� "4�ǒ��#֞�:�z<�J���Ϯ�A<p?��+ht�5����v���ũ.���w�QV���r�_����@�-1k�n�K�������
�TiG�
'�9�k��h��5#׀��5f�e,���?���)WnGB����E@��}���"}Mm#)�Ҟg�K�:ڭ����=�^��7����ԞQ�����7�چӓ��3�]��Ս���!�_4��������u5�PJ��q�����#L��j@B�.��d]0�!�Zsk��/�3�7�(.�1��rzfEY�����=��GA�'eY�t+�h/Z�VT�0JM����(�7��qF2߿S�j5�N��}h��z�>�7����3��szH�tY���$����j}��!	��2*k2נ��R���}H=8�?|��[����YKVGrD6o��vфە��@0�G����&Z�,G����\�G���cO��V�����,������OGD���UɈH���8�a�B!�ϐdJF�'.d����<�È��`� %ժ��hQ�%�=�#���Ȃr���ar�����T�hōS1�B��G��+	4�n�1"#��d?��hC���(��I	�h���LO�OG@�AJ7��5HeaPb��v_8��{R����{YB4XH�Mɛ<ׁ@�"IN��L���Yb�\���JĔ�d���b&r���6�@ �m�1���xp�,���F�JD,����;4�b]O�5)�ejn��k��mr����òl�4�B�*I �}B�I~p�s��Ҝ̦f~r�*"(�e)���~OX��ݦ� 
��u��m�@LfH*��}�	[	2���Ik��r�tl�_4,�I�k��0o���?N	s>�W�I�`�ޫ��9��D�\�AwۤԸ���J������X��{�JE�j��!,(�@F,D:�+�������Q�N�HSա��+�7��
�C3x��N+X��I��N�����[���"Аfa������B��+��Gg�<��-��h� 4j'j�S�#�ؽ�6;kݟ�J��^�7���I�Ƙ�_ePS�ل41�,��l��̌�G︼�ng���=v�r|�Z}�C(�7��\I�h}ab��.Y/�Sr�?c�m������^��ɮ�%�2�{�x�qջ�ȱ���}Lʰ�s�n���$�jU�X�&Ѝ{������C���r)��-;���(\�%-9���9�Ԣ�V�({	�DSe;O�e:���Z�_7ݧ��KO3�V��7����E���OԄ�h#H>��l"$�X�v��ȍ��4x�Qs!7�H<J��E�5�[7bO��|����s#Xa����r��[ӽp��1l;d]P�'��'��N9d��ѵ���CqV�r:ѯ��-vC�<$,���%�q�`$���gE��{�%d���ZKA�r�:XKꗘ՞����p���H)�7��I��J�X�7`�}�	�:fF�p�.᱕k-0� ���3�$�qÐ�BsO�A[v;��&�ˏ]g���.Qư�_H�I��ݢCuk�O�!Z�����=n�l$�h^`��PP@����DѴ�*��]J�F�0�]�P���桚��!�Tnj�l6aN�rD�ْ �c2��[6�*Wݲp}�;&�E3Δ3��5���k��P+>_G�M�ȡ���U�D�5���hx9+	f�,iV�n��zl.���Vθ����a�lo�<9�O
��g妐�ZNF�Q����0 x7�h2s����������9s�ƕV<���8V ��1�KÈme����O��6M�;��|;j�A[R���b�����%&�3�F=A�S�X^?Bo}�%�ё���#��x`pu��7��[-�	Ly�ݾp<����%��
+�����6��9g�M𖦇>�d�/�h#4�H)J3|\"������2��~���z3�J���א�J������d��'�+�r�a)ɤ=�i�d��o��o�y�r�,F���}�}�����' R�a��r��VNH6}4]�|�r!ġ�d����c&�[A��'��y���X˴�UW���q�rM�J�F�Î)� b ���!��\�d۪���˂��7��h�ݣ���.*��W�9����6g��Tk*_,�.�'p	%�>0푲VG��*g�y�7�����Kg��Z��5bcI��g�}������V`�9 %�[J���=Jޝ�[�l��s=���i:����m|�/��Lc��h5B����K����G[Y�xOSր�:GH��=�����?oo�	��þd�Ҥ5�h�}?pY��r���D� �����TF�t$�rh��'�o{����&߅������d{�cT/�2���`=�-5�f�!b5pk�nuf�*%��uXӧ��[F�]��z��R�\F�����y?����a�V"�uHNpWS:w��@��(�~L�^ZY��~���6����x��+}z����F��綫�1���K���$���= ���R�]:����B��' t1�L%�����c�5�5(��k��ۏi�(XB�r��z��A�Z8`p4�%3�"��R�I���񥇩 ��J���6y�ɱ�=v�A���z�M~��9������f��$�Og�ў�?�G{��Ҙar�'�Q`��dWǨr31%$�\��Ú�6!���
%��~i�:k��n���&[�)�^琐|r ٻ�s^��	��Jܔ��X3�IV�錦Z_.K+�aʱb���A9�G��_�AV 6��EV����Ak��@K�C}�"�g�	XZ����$8�e�%ڸ����^q���1��F����u}nҠ�5��l�T���L����i��5�}������uliiSS��l�?�:�FѠi��[j:�Fp�T���b�6Ğ�S�~y,�X@��ySI߀��Z�G>�ң}I&����1uA|`c<��.������!5"���=�3��]�r�GD
h�	(D�e��7�5�$�65����y7�]"��晬��������&{1�J4l������ەV�����|P�}R'���dWc��Vջ��p��lf���Nh��@��`;�w����Q!���7�@1�X��]>�԰�I�eh���x�V��ᒃ��m�4�_v��b1�xG������p�V�H�K$
��=��]�P5�k�bo��ʯ������Dг���=7�k&��u��i4^��J�����r�%������� ��|�m7W��kX�':�ˣHV�T����M{�0T�g#2�W�Vܴ����Ń�fwI��E32P��&Ufмڋ��"��LZ������<dfr��X�ᓓ��k�.�ɾcvO�B���>�j����Q���]�Й�v����?U'q�<՝ͷ�Q+�0�9?sS�H��w=KF�h\�"�m^��ޑ��LD]l�	]ee
՚8d�nC����\��������b
kl�uB�/�����d��21hk����3+�2x����W8������^�m�wo+\���e�e�8���|q;�0��^B�):�W��m�15�K\�u&<X��~�)a�7
�qqȪ��鴧 ����*5]��,)�=��=�Eo��g^�l�V�g� �
��m��+U�- �;��'�Zu�
-����N�8s��F����C��]�K���O2S���f����I��Ŷ� K�#��nK2�.}5��JgD��Q7��{	#$�a����,M:m��kaĉ42��C���kj���]̵\kHB�?�(�{6�]���S�/#M0+-�$W����&sN����n�A�����s�K��fy.�!]��,y����7n+L�n*�,�Q���ӗ�կܼ7�j|�jY0��:1_��eˢ<&��P��G���r�D]����A�� �����7.<份���R}X�ɤ����,���V���Ŝ��x��t�
������{�"ɐ0��zl۬[�u7`O�)�`�hC�*�ڣJ��d��ӏI 5c��c��/�vUhI��^��γ������8ӷ*�́����2�~�4�y�|����c^��2Fm<+^%%Ue����ho��	K�H�Ht�àd�Ln����uX����M-"�5���ݟm������yH�I4���dLc\�E�~DKؠn��w\��733��j��67ȴ���������if&���j�u/�����k�T�e��O\�Y�R�[�~�������	
L�w�A�s7�Z�z`Fd}�"L�ǆ�B��+�-S�/�mxg�G�o�$���m(��}|���Y��'%�}sF���UI\0T���E�KWG�&Z�%�Ym(%/���}�eq�Q�]�d��$��p�	5<iZ�	���ߙU�wA��������T[�Ĳ�;�u��Q��nۤ���z����������,m�|d_7�D�����uX��46���Y��YD���d����-���t,-29��*mn�>����E٧�[�����Ϻ�%Mn3�7�y����}Y�x"��v���=���&�À��]\��B�����2ޝ�t�_!S����d��N�u$�-��
�`(�3X��O���QxA���l�P]�lX0�R�����ck�U��Y"\,g}�U�Ɓ�u��ج����u�����-�nlW���I�< Y��P~$�ռ���S B����u���lkG�w%������bL[Lt_�{ B�Ɔ�Z��-����Sm{PR �tRA���L8 ѳnR��9�`Cܔ�g�^�d}��]
�yB���&`�N��=�j��	P@���|2��C�O)�������NQ�Ε�N�3�Z6��	����8�/��M*���5��b��m�I���oX�Z�+�>�z����Y�e�˿�V�d�CC��A���	�EdE5��D}9+��h�SC;\�{rT��Yo��s��DV�%��7�C��0׌>r�G��Nl���ѩf1�R�J߆�Ѯe/bK-[���
lmN�]�3]d�ܧ�����x*�,{�B�@ƣ_K��x~D[Qe�}Q� 3 ���~;0�T��u���#o�ye�ׇ���ʷ�w�?��K�Z"�㰗�sT��Y2B��U?�)t���&�O����}C�D��<J��|Y.��j�TN�U&��.����}�A���%��F	��?٪U`~��]��@G:�@/ʧ�)���z�6%�^ݕ���Q����S8�K�EoJ���X��~�Х֨�X	�Uܓ|?�8��ì��䑭�9���ET?0�K��S���q��Hz'���+�i��;���Em$�$%�B���v*�R�9/X��e0ۀ���J1 \TJN�X�:�l@B� ��� �Z��V�8�K����!�گ(��(��]�4w6	��D`3�)��^.{���ɖ��#"��E�k�BP��.���<4b�u�~l�q)�o؇.[?�fv�=Sb����T��o"=d8�3����6 n,����%/n��2��2�!��g5[ Ib-�����Xp>�ፘ7����$
��U~�{l�u���z�?m��s�����qu$��/�3!i9�� c��!{�:3.oˣ4Ki��?^Y�|yv�Q*�
���97]?L8�XA�x���j@�o6�h>Q�wG8��6�øA���\8����,�C�Y�p���VB�2�$�QY��
������W$ʫ�i2�j��_���H�}���#H�Kޜ��z��Sq�V��TR�Q!���o��}�rquj�fO�uR�X�ap�Vw����]f��mSm�x�h�2i���5��el���zՑ���@�#�D"V;���q	SH:#��F��>U�ŷ��o�����Y�s2����3���V��^���u:f�R��$V|�H ���n��������,(��wFOy���B���5���BE2@�ʰ�{��6TJ��	bݳ�|l%n��`]�O��qZsX�����[�+����z�Gr�v�|���Ӳ_E�Q�~˾_�'�JG��Y�~�
dN�� �4�L�,����0��>,��ZKLD�W�3�,����������\��EYtY.�[��1R�P�z�7��ܩwMPD��sя�^���z�0�h�"�+���3l�a�I2����.n3O�d,G� �&g�aS��S�+ԙD,ņdU�m��Ka�H��{I�,y��3S��䩵{���d�,5����ᵒ���?+��[X6�������/NS���:n��aXH�B%��磇SF�{���)��fjԤ�\�Ι�[��.s�fqE�<����-a}Y.
�!�Ʉ���P��˔�}���i�].u��
!p����XF�Y�k�8޷�s��8)d��T5Ӭ�V@�M U>�����o�=����%��#W�N�Zzh���N���T@��LnP�@G�v�j ��n�)9�D��@i[�ҼD��h���5�2njt��w�uJ8(jٛ�'�� �؎������Q�6ղѳf�ǙYl�{�lI�6���c۪�j����9�`q�7���DK�JV�I��-}K\���_��[�F:�x��q��8c�$��¬t[۬���C�ʣ��d��g��+��&2��[�K�x�v��I��Y2�6��"�UZV����?�V�A�VZ�-O&�5�Q���7�E5��;j"f��PbN�Ӏ9��jV����) $�[�2�e�;;�
}��'����Dα���@�^���&���� �ĚP�*,H[^���%������:�Ub��`K�{|�㧎R����|�Q���Bv �����I���89R����zVL��ݷ�̘�o�����[��dn��`�3�=Е��߿��{��O�;�$v�J�Ά�lz��R���o������Pw_��5�8�t�������R���w�~���OH�u�?mG�ǚ��8�	��2,��V���� �7�Q�_Np��5)/e�O��,d�΄���c�PT�~���-���dk=6@v!tʺ �C����䜌��,�~9�}�tcp|˽��}z9Ew� 	<�'i'?l������UMM�����ƀ$m�A ~�e��/n��<~� G�� �a��R�Yr���f��r.�� C�����%E����O����`�F�ڵ+�̖|q��r��`���c��#>F�{�����e�t����P�e�>������t�,P;�o�Z䨢G?]5�q.d�%�9`�r^�)@c)�^M\���D��㰙�����,��]��N�{���)#� ����%&ӹ	Y�d���}��=9���|e� ��@�Jû��f-���>O1/�RA�C�7��s�j_�j՝�>ґ�7�Aҋc(�3���p��m@?cw/���/$��K�>'�F廩˚�"Br�Uf�a>f�I��t�`	.���z��9^���ߟœ7�v�g�y$�w�0*�iK�:��K0÷+�J�G�R �-�V�fo؝��M�^�S�h���iY�Ѝ����� Rb�Ԡ!��;,/���%�a�ѳ��yL*"$�2��Y@*x�^&���߁�G`C�J�2�>y�N����V�}�@SL�Һ�4��GH�H"�־W��2����<c^ns�$���i�|鋞�J�OE�0|��� ���@(���"�d��E1���b+x���tb��F�z{�?\��Ъ�W�_����U��2[4rf��RW�f"OT5�8Ǵ�'�F��ywAJF���އ�Xь�D��T r	�=t̔nA�.|��4b �a��G�_J�:����h���l@9h���������t����R-��-X�ʉd�R��
�>����r��x|Q�)E�rUJ��Y`��W1�j�S�J]�ߜ"Ig�HΌ�7(W>ȼP�^��^{8(��a�")��|�;"����t��S=�Q�Z�bԏ��z���Đ�e+��JrK�S}�ܽv�t2s�_RQ�%Ǽ[AJ��@J�W��Q�������d-Q�)�nT%�.w%"��� �d���<Y�b�p�83�T� !�lh��A�'��%�<g��������S� �q���Q��1�,ڇ��_���\���	.6د�Wr
Pd�K_=L�CZ�cZ����?�@R	[M��'61�X��3�|�g�0���)���W���kLވ;W��,�d�����df�%�Uo�����a�5ʹ�`����{�$f���:aoޞ칼{(�l�G�mAd�n�p��� us��.��/4�����*�*�d��Ƀԍ
��IQ6���5\�a����N���/g!IRCC���JW�6��vjW�w��������&_`D�d�m��z�,r|	��k�2o=s:C��#�]G�L����_�&㊘��K��*c<�EɌ��扠������	H�>�|�M$�y�~��WH��ک������o%p��}	�7����4C�$u�08�cW�X�K�=��$��ԫ�,���P��Gp����\��mYh�ȩ	�i��xY��Ɉ>]�/Ul[��]c2c{p	����$�Ĥ˹$ժ��mb�Z�C�ܑm8�K2T�ɋ�Z�����y��!qTwh7��=ʘ�_���_��l�E�>�}sL���q�G�F5���xz��}��5��
��Y��Ԭ���C?6ϲ䃁�U��B�/Pә驌l]Hg��g��G&��$,��1���C�?��pz�+��$񁬢ۯ��>����K0�\�(��h4��5�	 �O��Z^p�F��I҉�a�L<; �[!����/9e��h�}_ұ��f�m^�˃��f�"O�y������O���E�h֓�P���[���2�\#���iz��s!��'�ehI
�I{<�6fy2B��%I0eglI[9�<pվ(o�I��\_�9�q"W��T3b��/�����r�%P{^1k����������i䁒�j�[Z�7����z�8Q�'%��Z�@s�k��ܰ&�K���X����Y�K�_�]���>��]�:3[��;�pa��a͌�]���cn�'��A����DkԽ�]��:
g��k[Ʉ?�y2>:�E��g;v���X��(�x�M��,BGI�qƽ�ę�jj��6 1��J��l��*Ꚁ���)>�-��"�,�{L>8��[����t������4�n o)R*���\��Ҧ��RX�Dhjo#?��{���"k�ǀÍ�v�TN,oN���DdQ�o����٣��iE���ˬ��ӫ��Ԫ�.X��՗9�h�
;g�_(�V%�yAGBWMT�X�IURa�8�J0�i���A�[։}.WXW����$hI]]�Iu�4={��T��=�������J�Eo8�L�rV�%v�>�9$����� ��=Pi]���3�:���_����~�e�o�3 /%���Q�Кf�S��@[P/�H�)Z���J��Z�<7�E�%\֞���gj^Av�i2��W-��1Ym�I���S
��Ћ��s-汑�j��6��>Q�t̖F]��KK:�rG��wП��+K(���F�[��(�7��G�����&�4�HϬpY�r�tU3Ɩ���~k�靖鮸�ڼ	3��<�Ӡ�����#���w����x�U_^����_ic��э���b��<>B�u�x_�ڐ~�:����A1&�x��ı��Ecu�1�d���ȹh�J�B���o]֣l���>�;�{S�-g! tdU�"��kK�d	�1��M�a4�L9�6E�h��B�+4��(hdxUy6�'�5�z��M�2�4���V�
ؔ��#���C����:�3^p��Jt�q{8st��xH����$w���$n%��޾�"A{�3�p813�F �o����i?0_BW!�:_A@���!3��=�\�ۢN���+-!:�N�S�8����Swm���P#'i~A�{���n�5���S+|ʉ~
�� s�|���U�垳�5��e땲y8pz�����P�ks��OO�4-��p���+��Qp��[��~(�3b�,������N-Q�FZS�Z"�o�l ��0B&��x}�n����,aG��#jpˌr�j��0�O�&sC�{��E�G�x�hUZ���y_���0<��q�#�q���e{_;9р�!�uxy�Sf��e����\�k��5�7y�i.�.m(˺���������*����������~�HF����]���ojv�P��� 23�5� ���RG���le+��nI2���k��uPR;�'���J7W.�N�g�L����)��W�lF�^�P@w 
�~�&j�')j��V���=���I�@��D��e��"��z87�*A��W�$���2��x)�4���6�~.�v/��)�^��o)��,%�t�N�����%�KI�Wf��¡���bl���Un��ON-�u>�_rݝ�= �����dX�{&L���?>�d�N�W�5 Ԙ�Ў��GG���#��;�ܞ�t��q��FR�l-� ]j���s�ה,(�[~��:�`�-qk�5q7	,`�1�U���L�����sW�c��/S�I'����5r��i&����G�p�����S����}�C�����7&��Ȏʃp_������ɨO:F�3f��E��4+���j��sD{��_S��.8l�O2��<�M�7±:S���g�T�E���L�������&`%o�+�+�-iʾ�RQ��p�	=���mo"��)�a7Q� <[z�W��x�a^:0�ٜ������4��JA`Ƭ���*	���.� b��z�ےZ񉺷W�[V������GÖt�L���%�Iz�\������Е���uJ"dW	!��yZ��ߍ�����x�s�4��`��)�8�aF�֘)b*ͤ��]n%n���4<�*�Z���y�Q�`d&�]��v��@?�
 ����s���1�N�ñX?��z�l�P��Q6�^���sΟ�(�	@0���YH?Q�ϒ4X�q�;�~�.G��L'��v>$v����h�K�f<xU���u����E�����7&_:�bd�h\GL��OI��E٠z�?��:���_��?��${���"��
��l6�����[�P��ڲ�x��@�Hp:V��Ena��T�(��$~|Hߒ��T(F��r�Iͺ�ۮ���Տ�g��g8�����Μ���EأN���qCw��X)g�' �U�&�Q�z�]钄�|��1߼q��O��7�A�t�����誇��B�I縩 ŗ&��>]�k��K �s������/)?����?��"Xx�f\�*�x���<H�m���82s�wT@ڡ���kZ9l�B�[�P��e��rع�@��(Z��AQ[z,o�{���ef��y:47��"�Bb�c�s
6ɤ7���8
`$Z��f���m�5ߺQ(",�&���� ʏѭ����u���"�19Ӂ�h~؝���_86���#�),��rspBx��ڱf�-s�I�>sCM�s���$i߼�
��g1��(.�Mgo-lO���P&f�?W��j7p�)�9�L�O�<{mG=��x��ps�ߓ���E�Ԧ�I��� t>�4��SN�2�����l�S� �`�WS%`���(n��I�,���2��[�,�y
�zgO,C?h�Y�DF��Vrڜr}/+!��ǚ��� �P�'j<)s�R���Dƙ�+�pZ�w�
�S���.�n+��a|���ps�����`�;&�a_P���N)��1>�/�^��8ʟ �����1A�l�vDۍ�k��)zB��WK��g��=*֡�L���r�i[�fX^�P}�!
Y[��G~�Oll��w�7��{�9)~�hY�'!�Z�qOm�a�������e��Ev��t�(ݏ��?�bV��F�T�t�z�B��?�S?��@Mw��&��CT!�s;��&}�,س����刦�*nW�{�4z�	e�IBVd]��/~8��������Pao���v.R~��_����x=��,�S]f1w.���NF``åd�>g�3 �;�3<�`��w�����"�0�n.^�t�j�U!3��>�h���Og�IY_@"�`�cVs7���������@C+	��=���ŻT\�z�n�3v�'4�lD��6M}�7Rr��m��#�W��6���-���N��d(�p����`�1�3`��Q������)��?2?
�7�7��'C2��[TH4v�����g� �A���'j?�u`$��@�D��,@�8��`,�t����V(���a��\�n�c<��*���r�1��gɰD�x�c����o�~�ˣ�G��g��1\�Ռ]Ec%U��&�mp�s�U�
��y�6H��.�j����☆@g��uqWl�Ż\����~B0��5	>n��8s���ױ�h��#���"I����#ek�d��˒a�dnH����X��c��"5ƎRG�q$4;� ��.�i<	��н��~h��4�K�Z
��c������mu-��a�-���O��}��ĵf���A0Wr�c #oi�O�/�1qv���_F��z�3�*����d��7��n�^%"��3������ק�u5E��=$����$"��n��w��Ϲ���se[�lubk�?6���l�����d�����!���)�fB���5H�X��M���1�t2�k'BqL��|'�AD��D��2� ��U������̳ ���{@J��y�2�χse����:+���_�^?P��t�����$�-�A��F6��on���'��Tb�u�9΍�eDS�� �i�Ǭ�m���(���ܢ������f��#a�|<#@+��sm��0X-�Em&�	�����1�h(�byҴ
� ϕ�������?SMA�"c�9O�qs�%�MɊ�Ɵ���E=���OӲv�� �R�����x���b����a�/_#��:���l�	\��&=r����u�V\�%�u\F*�(����8YW#GS��E���.�U�KE���%g/b#����l��x1`��o���s@��`'�צ4*��MV�I^ui(X��
#�����%f�6��J �5a�y��	
<�JD���d��[R)����HZ��y�}1���jH���pz�!fts��t��=����
El����^�P���G�h5���R[-kyӝb �)��=�dNǵ��5L��P��ECnn��:�xF4*qpϘ���z9Q��䠹{7�#"�(��>m�F�)kHHg�B��S<q K �/Y*�XYd��l)3甡��΍��FHtGc0#����!ݩ��on�t�}�k5�G�mQpc�jT�E��-�G�jӵ<d]U9�!>��0�t��H��W���4L�����Z���4b9pIN�`�ej��w�9@c��������N�bBU�,er��4��������^�%x�*�q�j�����C���O�ܞW=�{�=����o�?;�E9D�Y]U�_���}��_?�Ǻ���`�y��΀S@+�f5 �\�N�v�E?^>[��phν��{��IFѹ��J���؍ꨢKP��
��d�-]ܡ_S��2	PQiL�B��y���p��+V�齕�cM�;FT�5��ܲ��`I�_�W�+i�wo�(��?Qlʼ����\�s����ڟ�(��¥9���u�cOx�VN�@1Z���r� ��L��D�"ε�ùhjl<rQ�@C��(�8Q�v��#�� ��i��G6t�Ė�D���Obץ.��c&���m�>�4�ͲV�h�U>�oP�`h�e��1�kt�¡%\��؋O�'$`Sq�b#�,�G���:�h
���r�h����{:��{��O�{�d0y9���!��06�hΚ2{�vL���s3'�5g�n��׼�9��s�z��4��L���0�����������H^3�� �m�X�`x�4j=�+��KB]����KɪA�����$�y���Br4�����:)Jj�Ċ�:����Q�Jg*�A!�e�~�l�����]�c�#5B��*�W��j��}��?���>��F��4啢�@�m�����Av��B!�f����|^�?��:�:5!��2�V����{�|���R�V�D_�a� Ve
H8�0�AH-\�oƜ���I��A��)#�xm��d���!�ƿ_nƣ�<�h9�qrb���v��!(���L'�ށ0�d�4H�g�XG4�v�$����؛�v��f���l7�xˈӂ�q/1��~6۹��M�m�&�i�v��v������Q$��1Fct�$rۍ��j��4J[�z���i�M��(,�=f}����A���q<���@��e������~�5��ͭf�(77��c��~��za�G�jX���(b���D���>pD/O�"U��4�f��J�ٺPo��ssM�1Rp)N��"�6G�r���-���yB�0B�4���,�[��ء�M?�i1(�S
�e(}SC�Q�=g�ѕ��CZ��z���ޠȤ��;uQ�Ӿn�nvv*?M��l����p8��W�'�͋�ר��h����-F�V��a�إ�{�s$��o:m�$i	��Y���t4/�I�b������� x5[&�9�~��͕�t����;2M�(�4���[a��ߍO��������g��cť�D~�zB������0Ō��W<?���9�a�3���Y�V�`4������v����VG���.�1�X;�R���e�*N��$G����B���g�(Cz�Yj1���N�\�'�@����Ź�e1�u�k�{,XgE��ʈPY��;ʊ��� [S�C�aBqي�&�g�o�o?�s�HG�$��C?i�_�/�����#*�)p5�Mֽ���z`��0�>���F�Aw���D�{��Giq.��+�(��={~���^p�y�$�xl׾�߉���|*�0�J���H�d\��C���=�a��Z�#��qf�j�/�P��x��FǊ�#a���&�¥~����rG�G/�`!�t�+�H�ȅ3�!z�Vj�m��_�Q
ο	�)e*z�Hu�A+繧dr�i�Pe����j[�^g"�-�t�N[/�TV���F�-���-��D���N���k/���׈��Y�m<�1������*�%�� �?�On��6G��<�e�,��{���ѯz�
����|�yjG���F���ߛ)�����Β='���'���C�0t�d�#�ڊ�M]��	����vBcZkJO1m��$�`��w��1�I�'��=M�F�0n��82ܻ���@��|�U���*�������M�� /xJ���I�:	������.̆YW�I�i�=��*�JH駐�w��U�#����)����}p��5�uE�����)�龑��t�o}�a!pU��%�/�lzX{ �ZÓ�w`,�k�E�A��f��M*�N1'[$ۛ�*1�y��s�%`�ȑx�뙢@qAx�,�Ɔ��Jy+�@����ʻ�s��1S~ ���8��:���R�Z<t����^	/������]tI5]��K�Csd'v���<��v�Svw��t^v�r��`��ʤ���@C%�W�§�F���MJ#k�?{���uc�)��?X}�?�?8�os�em>��0�!{P�=��|}d ������#�뜨M#��@�󹑌_mi������8��H"�Fe(IXG��`���9\p�3J��v�>q�N^c�A��1��Ґm�	�l��'.���T� R%f��.��Z	E�����z��CP��-,�/W� �iL��O��Y��u���v�ו���N2���b� �W�(��ݐ����s3!�D_�FO7|kZAȒ��$![��G.s����`5��B�,��$��CWج���'2Kx������Jr
r�"������ۦ��[�׮�X�[�Tw�MIރ��=@��A��N��k�&����(25��	� {m��sr�������x{�2e�!� �G~$&�����2lrt��hL�[�y���B���zǛ�����G�%~�w��ѳ�b�j$�6���-B83�Vkl��f�P ��e��|!s�*I��5wc�r>��jE�L�ޤ��v�u�e/�+7�q.U,� ¦�d������b��܊2��f{Ao?����C�<k }F�E�^j�"�{`sd�S0K���|X�~����e	�~��iy)�'�2��c쾊����X�|��h ��_��z&.�s��ը����G��<͊����� �z���+�JȡA���Vɀ��s+*� ��8��O��V�Z��*Pְ5�&�ъ�ƴ��}N�*�Dxbd�,��g��osDUGT'�b;�{��T�|�L� L9)�Rv�5i����Jv���r9�L��v�`���w)��l�o�^1�������[��vT]�Q����ł�B��-#�������<Ro���~8d�N��隁���q��_#��a?��Ͽ�Е#��vPpB���A��^Hl�{��S�{���T|-xp1Y:~BM���P� N�L��7+���f��KQ�-�%LG#����:�����SD�Z(��'��E�W�m��C��p( ��['4��dgb^�0?�B��&[�գ?Ӿ��֘҈���¿��u��+�圻�<�"�"D%,gW�����Hy�Y���S�e�&�'��ےK��ī&d�;�_��'a��4�������r���b�qem�<����*��_>�q�����.��[�`�r�.�7��T���v��6�Ą�M�R��TjWS:R�3lW���\;��%.("����I>zCdM0mM�]��arB,�T*3@���s0]%V��q9ym񵘾.��!l�\�E�yt�S~7�_5Y����І���i���;i!��^�gpU�I2�4�y4��՗���ּॄ@�ӟ��ꚠx6.{���;(Z`'�H��SUV��E%�zp�Т4&ӝ1#��ȕ��\����vF�����}��(E|���	V�'$����YmRЯTM����4�.�ޙ�_[@Ye��LooF�k!�"��I����k׼s�G�d��M\��V
;���Q��ơgYd�%c> 2�$`Vs&��3�>iyk�R
�s�!ѦN`�|�-{ ��Jɠ��M ���\�$�G�S�򅟷���q�'�T�z����}��gS���~��S</D#s�|��N��s��n��LK�{[~�tKZ� ;��_Yx��%��H}����#�0��7n3���j��w�Q����%U�氰m��d]�ڊ{�_��3�C��4<���]	6Z=W��"�+�c��5U���M�&�$<�JhEz7�=��F�"��@\9��u�\D��?���E�v����]p��d�����'�a��vTƑޯ?GJ�G�Ps�h�l��B� �V0�I�i���e�Id��S�R�*@H2��6ۯ�5��b�E���*a�p��y�4Փ��/����X��G1�f�e]�ͮhMA|����6�f�t��&v�̯��w,��"l�B�J�B�#�8u�o{Өk�m5F#�xs�
����џ��?��~G�to��h�`�_�ة�D��ζ_&Sh)��3J�Iy�vel�������G�M�M��������?���F��*�c�i�lt�b3��Y6��l�m(X����"%Uia��UQ��f6���S���"�)c^�n�{w�ؖ�P�Wqd�.*��1�S`>ʹ�����x��^ `Lr�Ѿ�f�5��J6���L��%�Y��g��st)X����h�s��n4�5��� I.�p��G��e�$�f�޴�q��G�&7�u@�4$�[�ZS�I�M�%ʣ�m]�(���_�6�@Z㞎Do��4�
k���b�Я�D������~`�#h�~`��4w?7���w6h�bl� ��n�f��8.�d�)pXy]�4�V��鏘ah4��Ȳ'�i1����P�D����	�'��hG�|�NS��K���c�ߓ/���jC#'�2K���Y/����d>4\7+̄#�sަP����A����&�1��S��~��Y�3e�v�h�8�_0DϟӇ;����{�F�PR���X�o��e��~n�}g�8��n��
�����Ձ�}6.�W�N����<�w��n�ԛ���@����gv!��
T�l�4�n���T���I�R$o4ͬA�K���oW���p�ץ 4�x��yTTA�n�-�؉h�&<�o	U�
�څ��q(�	�2��4(n�ϖr��i�=M�pr�'6�dcLad�	l����e����ᙂ,;r���k ����%͇�@�����ZX�s���>�'}�J�#�U�2��§W�4:��*�h��6�[q+�W@xmE��:����L~��xh�<���g���`�]��?4w#�>)F5x�^�Oit���w�Kj�+ߙ'Ɋ�M�F���.�Q���Hr�M�Q��iHzA�v����(�.�, 9���SJ7�d�"R'�oW�5%"�-��ET�R1*׺0�}=���E�64r(���x�<�[/lѷ_��o��Pl~Ia�Z�u.��7<t]
���������G��}�Iצ�?YG�����	�ʉ����j�z�_v��nR��[�����41��H���K"}9�(p�ge38��J"�;���[���+8Ҭ�Ղ����Q3����P���2j��Qb �& ��j����%I��}�r����p�"��_�<����=!< ����M<4Z�j���~H�����jM�x5?��С�(���qн:e�wVcB:�4�<-飕E��.�U�41��LK���c�-2Bz	���Gj'��NCyr%u��i[	��GL�2��x(��X�]�K�KN=�Pᡵgͧ�v��m}+,D�8S&i�y�e�!�)I`����l���o����t�U��I� ����k"J�ƽ
%�@xW�mX�:�@M�Mbt �,&`8�$3>�<߼?���{�w���rU�6����r|����D�l3<��z�8�Ġ�o�)wx-�~6�e�����cM�����\}�fZ̝B3~*�3�"��M"��
�F���b�<|;S����{qHs�05//' VG���ށ�ki�lcN����N�4"'U��>�|)s�c���-���J���X�������vwT�=�B����+����f��]&vȓK�6�\�'Ks��T���]~^��2v��$�썪S@bp\�A����r^���	ɉA�*�Sï��9"�p�qۊE+��B+ǩX*`�5o�{�ŋ14�ُC�v+zG�G~�7^"�k�Z���Α��kw�g[w9qq��ݝuز�4q+t�҂t�{uz-��[��i���4�dC�$��ʳp@�f��DE~��	����Z�Æz�Bg�ە_�fB/m����7����<Rʃ�KW��t�Uek��8h;8����kdv��G���d��B�2H��X����F*��(;>��DdY@�n/�Ꮴ��m��{��/ܴo2���������8��-C9�;�cł�B
��W⣚
Af4����������x�������CB��-��Ł
�� ϕ�Oױyz�	B��d�J�e�'�Hy��\ıu���o�8s�j�������N�	��p��w�ڽ/.����$����r�o��n�����pm[?�B^~�ȇ���Hj7� �����)��y/S�8���SK�Q���śO*�[^�7`'�S� K`�>��T(Y�lru�j���?��1/�a���ٹv��<����P]��擽�'��I�^��7{�!�;m�=�������]��'c��5#�S�[�9P���ϋY�'[-��������`88tI�T��oNwvhٝ��V��_HI�S��"Ճ��)"���D�����0���g�#�o=�F籵��O'�����Y��Q�{Bt'Y�!���S���Oc�8������B�V�휻�dN���AC#���-A�i�ƀ�S��[������ ��-%.�xl6a?An'�[���!T�X��"�9œި����m]�6�I��dD����b1�o�W7�sҨ�%�7t�z�FXAk�嗉]���
o��Tv�&�=�B+�=#����H/��x�7W\{�b�18R�A�λ&Nld���`=uVKo�G}"&0X� U����$g�W�"up]����|��u/�/�7�㡌0Vk6�ia��z��nqp�7��{�S5�4�PÅ�ʴS�5�0���9XIg!P�Uˎ�	1����)��j�N�6�Ɯ@g����07��i�c��CR�n�ԻE:jV�g/��XS��1^�Ц1c�6�0�i��>�B�G������B��:p�	M �a8�%fkN�4�o����)~%�x��� w���:�>I���b�tc,x��틪潚UV�T�=E#zr������K��J�����c���$��_�D��t,,eu0����a�z�OW-z̭�uHQE�p�\�CS�|�`�팲me�oXL�7m���p$5 9ח��`>��3w�==�z���{����T�#�`�va3}j�f� ���w&@qF���&��,+i�9�|�r!�-Ȋ���r3�5t,�~r���L�r�����*
Pw����S�F��q$�Cf��",�����:q�V�[k��M�-๸�ltY�@��\����\���e ��#��q�bS���^�%���Z�b�&�@ �K�D������ئ�*��Zmh�#���f�9�G�m�9{�m��G��d�� �Kh)X�J)��( >1�C�6 ��nϕ>%���G��t4��1t�ޒ�<��7�B��Z
M���bk(�<���Y�߫�a���D9��9ldF)'�ŅK�27�7WS�F�3SC/����;�N���ۼ�V�@c�e��3Xk��ixص����!�J��,��E9+��?D눽jx��c7c>)F6�g��i�7� ��kV�CN"3?�蛄��P1��k\c���w:h7!�5BɎ'��	^�s/٪Q�#[���/��-s˹������y_�����<��F���{:���N��|�� ���j�?����a��|�=��f�79y��8l_��@���R'���M&�6�嗀��I��1��Vw��9����Ap[)�:��ad��������c���֏�i�����W@*ww{�Y���8�\q$������b��+��(͏eWUM롫�5�%��tdu�C��۲^���R�l�7׮˝.�:`¥w����P�C7�3(���j�{��s��Ш�Y��"{ȳ����=��'6|۱|1��9�ŢS2`*�<�y�w!��c
�1U��';D��8������7*�@�2E�<��d����ɼN��Gߡ�Ϳ�f,�:����9e���'�2� �J��H���r�j~�j+<�ܭ�N�Pj������@��p5�'H_A��¯�L����Kp֔4��[��(*��	�<��b��22A�(���7��d�[Y(쐊�}ȳ���|�.lA��=>�G"����C�2o�M�Q
E�R�$j�z��s���/.h���:�v����r�wzm��FͲ�e����o�P��z�hm�HsT ���):���dK�<Z�AGm}'���S���dv��g�S�B�T��;���(J��j�øݖ�w���9�/z}65{^i#� �NL�a�
� @�調j��]�b5߿�m�Cr��-(�k�����A�Q����r9��uY��qL�F^ڨi=���WΡe�	�8C����P�����V��+��O9p�8L<�j�u�;Lɡ���ƃ�V��|�����D���cbՇ1��ւ)�����	:�j�t�@��+˝��╧奘����@K~t��@�jj��ob)ǿ7��7h�7��&u���d�"n�

#p�ϯ�V����@������j.���$��4c�^1^�����~��GU�Y��'�@F^'n���T�l%I�K4J���T�%WL�^��ct3��(U�Q$F���Ƀmpg�U2�>^��ɝ9���JA��b&�_�.��q��4��N Coӵ��.9e�K���fd�R�v�ah�fr  �e�;v��+�ŝ�3y׊�V�{|OD�z����KT����U�F �p�YT�1���r>%Y효Szkg��\�y�w�+8��2'9ȳ| > ���1p��a�-���kg�VW?v�P��q&0C��g4��,O�0Y�')e�l{4fqdO 8�3KfR)��:-V�\WBb&Tw���h�4��Y��AV�����n��3Z�}�(#֔�]�U\��+,��ȣ<S"xBiB~���Q�~�٦p�o�û����~_o�T��)o�S��s�SE�P�}r	9�e�����{+��4݀Gţ�y)���fW���UՏ��F�JW ��b�Ӏ�gFI������Ba%-˝�&�R�$'���)ɋ��y�V�؟ ��a��q���?"����J�����4ʟq��h�:�жӏd�ðY�������s�u�����"b�54�`��cb�M��r(�����&:�)��)��]`Ƚ�9@���Q�|�a�U�ޅԅ����]0�Y�(�/L�9���	H��l8ӽ�X�f�VV�y�T=�:��(� K��F��v��C��h�za0AW�,@K󥝑����Te�Z^bZ��=O�Z69v�����5����V�)܃58��H��<3�zPu���t�X��e�Wѫo ��i�]MGF�!_%\���T�1aó����q(NTk>�����ܷ�vu����k�CG��5�?ER�uW���&x��܍�M��(�G�Ń쾖��n� �X6lI��ӪA��ý4J�L��
	!Y�o5�d��>ص$��h�,�WQ�u���"Q/��Ł�A��:ʄ�/�@ŴHNw�siV�(��p�yif��.��a J�a��^���|Ǔ�7�VD	�F/n�P�tp\T��P��8��R2���z�.�N|�s�ݬ�=�j�t&F@6���%
�[GZa�5�!Q�ML�xyXe5��_�֗<q�V�~:*=���rZ��eGMX�P����R���ź>���PG�Ҧ;�6��gq[圝�	�"'|����j�dGF���T-X�j!�%�Z�Ƿ�\�`��d�æ�1)����u *~O�qV�XC����|-)a�E �d)�,˧�w�Kڢ����fc���A���󜛑o���U�ǉd�c�G�ՄwU}�4h����w��Ļ�˓���K�IW��lB�$��)Y{�3Ө�UC�Y_ΨY�,Z@���~�� .#`��^�����^�O�j���^��NE����� 	���[�P@M��2V������7~D.�X
�W�(f	���aʍ��&�e�� ���{��G��:���	��ȳ�7n�}�f�g���dnTϢ桎���Jw�4���>��ttc�-��=�r$���{ԙ��!�,�	�N���s+��'��'���]Ԇ/��۰�ha!�$˭
�:��&��M����D�n���ıo�>�����2?Ll?�#�¾��e0G�%5��~���E���-����K 7�Ur�H!n��u�h�~b�/S��s�ʰ'�/Ys&/�����ԡd�|�]�i�0me�X0쳣K��f��]�a�;�9)76~<��{�Q�%�"m.%�����E7��wTi����ֈ�g�Z�/�LjǵoT��y�t'Ɲ 3��;�	���j�GJ[�F�9���F*,�b���>��Kl�'_��	-u�ici:لW�.K�-\�V*�Z���IVN����ǻ�E��Sm��YͰ��A�e���p�S�{T����<�Jp���� p��FS�@y=��˿��lO�8����x"�F'V,ʄ[��,��8TB��X����}'��KV����I5;�7��۞���$��@-��j��[���X��9@,O�����.JM�h���}�,�`M#:
�B�6Ρ��s��a`m�˚�@6��tJ�LS=Z��oft�9�o�E9@T��k��k�@	�4(�m�wJ}ڠd�00\�,�`;H�8�'?�����	�ĩ7���S�����N�=��;�h�/���@���"�0� ��s0h��*�� �_�!����rB?ї.ض�E��g��˱���EV��Eo�8�!��c��ͤiw\ஔ
F���'���x�5�jpϴ|v�K��w��.���g������d����U��#[<�O�9B.4�4eu*�~�U?Z��S����K�c������/���q�E�gH������	֮�T�Ԫ�'��慛s�O۫ϘX���CKt�Ziz����><`-KQK�q����P���E?�?�F��蕣t���N��4���4N�ïU���2���qk�
z� \�!N��W�����;[��;k�*ͤ"�s��l)������%�%z���0����#�4����;�UMd!�rpuw�G�	F"N�3b���v�g�� ��6��Q?�����6��:��)M��l�N(���æ ���ȢC%�ї�l�Zx���5wK���l)�h�.F����T�1S5�W��~���������D�"��.�����yؗ���v.�Q/V�ר�,&��Z�O)��U��F);��2OQ�Ǫ��t��Y�/�s��w��_6�T�T�㗼��n��n���A�S� ���&z��|iϖ�<�Y�H�ö�~��ť
����7��1 M���@�)LJ�nWb�n�}1%@�[�Jdh��֓�ɿ�c���˯��E���D͈�;���čo@��J���s	�n�Q X���R����xk�ޛ�	S�뺗�<nY��M�����.~Z"�>�����FmΘ^�<,#�� H�����G��1'Q-��	[k&؊����P�o�*jܽT�mMFm�&�D��-b��k0.R�%)K:�^ޙ��lD{	�i��+��AÚ��F�n��O�O�d#��txC'��Tf�x6��9M��l���u�sZ�֨w�}���L�%�H/����(�����p�g%�����^�w�Qf���\)ɏ�8�R�5��E��C�U~̌�_�<u���2��N;Ua!�;��z�UR�m�ڻ��_t>[�4���-���;,օ���T����� U��?���D�H"[��?Q�X�ܶ��6ޗ\�3�)�9ؐ��gi)�;���7�`B��Yt��bP��Q�,Xpd��e$�=@��q`�@��`t�\�4/sR\xiA���2	���3.BN��:0#"G�SƯtϖ:�8w�	���լƌ��/�ޔͬ�C(ǡ���~Dn�/~�Zs�O[�cL��I�[֯fVr�.%ߨ�`�#2(ۑ���X���f���T�T1Q�Oh�;�zC�W�_Xk���εT}��	�=]�/����K��Vz�rٞ:H�M>�� ����n(���!5�]߀$�vؕ>�W4@żE���ڮ2���A*R�����y�Zid?Q�sY��!!8�"�>�~R�Y-H*�Aܤ=�g-;�Q%4 �o6���KA���3*r��_�u6
X�g�;XLXvx��U<�/#x �z,��2��<k���]`�F|s#���X�/C�P����ro��5?�>y6v��:3T�ӳT��M#� �3�M#�w�yk�Ž��*�:V9>�6���_CZz�����E�\MpZL�J�u�1k�!t�%�[Ƕ�sqN/��$�A�)��QXӮ�����?� 0vj�����d�e￲�c��y�-_=���OhF�`n���`��ϳ٧`Ƭ�����G��*�����v؟G�tBs޷�1��3��W��bx>����r<��:tp����a��� �@ɲM��+�F��;H4�0`�e�	02%��v���ٵ���'�En�=�	|w�)ee"��O�"%�k���ap�U���d����[Q|��h������'�n ;�J~T����%�Z��IyN!u�@7�#R-,�4�Kή/?K���m'd��;�"��&^�.���[�^eKJ?�(�'�%��K���h��R"TKD=��*�<��
��Sp��Y�,��?G�����?�C���r�ռ��њ��{��`~6�D���˜P3��]�)�T�4��t��}��5��f��Sa7׶i2��D<�
�㙯����ǷMض�E2�ơ?��)��um�a�_If��Ő�B}s�S�D��<hI��;�f���Q�8]��5��NA�W�|l<����=3j�Fi��<��rZC<8��5�����~&P�:j���o�<��W���2l�K6@�;v�7�|(y;����
	:x2�Y��:�k�AE������`Cd��϶a(�{3n�|sf����r���X��s��\NcA#���b^�� Yp9o����4F�=��m���Pl�s�C�l�޹3i���[�%��"~����!��1�C�r�Y����t˸���chÄ��w��3U�Ⱥ�o��_+��<���)�~/�+"�(�E5F��#��Y��ɤ�{��;1��r�����G��z�rf	QѦnn���/�pCUA��@�a�P;\$;n��u�G�<	G���3��s����T���"!�N��J��HO��=.�e����t���'m˂�`Ga������J�/[���?��ib�f/��B@��1����2�'�B>g ��u������iAJd*:���oy�E�`v�!�V���=�&�M	ٳ;�����VƘr��Z�z�����.piL'd��Zݢ�}���K_|$��v>�P#?Ӟ�w�'׉P��:@�b���ϭy�����g�S�v�j笳���'����(���+�t��},oz6+��TMc���*<-�CxL�Y��n:�
�[V�b#����������Uu�mY��V?̖tRԦa��C����Q:�/,�s@�sT5����Y��%�r��m���Q�Q��3��������:aU�	�F��<�־+�|˃J�)�&����_��Eh!u?_�A�x�����5����u�r�Rim����E��Y=D���l��S��T�}9Zy*�~/<�E+<�P:� ��>�)�����v+�4dx|ڧ�<\Ȯ3 �?��.<S�"�� N{�Խ���Q;5,�����ɉ�Iv-;v O���V��g�p���Z�� >�*��e	o�� ����I�>/�E��J�� t�<	\#W��/]/iY��_|��g�i�lͨ��	��zܭ�����6�5���lwyU��I�G�����&2	��9d���?}�\CA�ֳ>��4!�,�q�b����,%9��	y�L�ir�]K���{E�F(N������L:�D�ڄ�Ç>G\�8ƇZ�F$���lu�����
�c�./+�K`�j�I��j�	�_�,*'F�$3u��<�a��w�%u�6��ƃR�E�mw�Sk�{G��e�K�I��+p1�t_�*�f��g��b�5�tR�x��� =~N`b��-���]0����K�=Ǩ�3HS�B 3�h=�3&�P��:��ҧf�F���_�h^y����|�/SiZ��M�=ck�� ���2��D� ��~�������Z�dg�;>�URS�y�{,k��Tg�It���An�}���pF*#�T%���B���G�̒Vk�?���_���~o|tz=1���߶ʃ�~�NEM���WJE��z�O�$�Μ�	=�˲�zO�>��79��q�U�b��Y��+�gB֝F��[�e�G��Ϻ%�E��΢�V�
i?V�5��+�*��V�=lv��䟍�i��d����嘰Q1�&JH"Zsk־�,�,��DŅJU���y�����.ZW��)�·�H�ŝ �.����L�M����b�ؗ�s7��7�.��[KL��қ�7EͲ"#�m��%�x�MQck]m���W���.���3[ q���P�5�]��mhd���ǅ7I�
�Z�va"_7ځ���D.r(C�aj���^�|��(���Թ`�/&�97׶e%Œ�r<�Ȏ���Nht̮��7�gFJ��E���q��
?^��O�!-���6h��^�����!�^��Ai�E�V��5��(41�},a|ô��<j\M�u������	�UF�Ϻn���WV������K�$���E7�d����\"8fط"�{u�h�ٶy�~]�/wzz~J���c�R.+B2K�Nِ�t�a���n��	�u0�8S6�pi��K�)�M��d,��;A���)UPJ�<Vjm�O���a|V���VJ�,eڨB��3l̽��E��B� ��p����f/4�:-�C��
�D�8S�� �9�lW�J3�%P��XVo�w�U,������S��͛C1$��p�-1��a*��C��ټR�u�]��T�d���D��Ъ^ܓ�[^���n�#��fл�5��A�:Bi2��&1�w_��Wq!V�膨㏽�����?7�o$�&Th���e��\�_����(<c��m��S	|ā�Q�(��]�(�5����(����*�	n1�1���s�ug�lɺ�,��^e�_��-/K3Xdg�!|ko��h7���3yE�-?[�DB��$���ѵ�n�a��/�o��c��J��Z6ͺ�S�`��Y�wjΎ��`Y�>����������e2����ċ�#!�i��1{1����]\��£���Ϗ�F�?+$'Л%�4Ԏp��f�CXޒn�B!��9��g��M���_�>>��n ��9��'�0*V__U"GH^gz�䋛a�p)�&
���b3Z���A{�/�PSy��6��dK�w�}έ��kiT��u���z����*1�}N�:ЎF��V�|<f�Պ���@�y�Rs���]t���fC���h�2>N��cM��(��Rƿ�.�t?E���Ŷ���J�5���ю2��^BW��̼�Z���4�ԲԀ�4R�/$1h&�<p�e�C�[A�X�0W����l�k+����'դ��P�]B���|�|�u�>F�8�t��iN�n��6O~�P�\J�ݲ�B���r�����@<����^r��q��S]ngL��w;S�ױۦ4u|���*��#�[���	.l��J�C!D�4�>n�����}9�"��7��$8�_����}>���1�ȇJs�s���#��N�8�� �G����^,;����� � ��2����}�	)ry8<�_j��8;�s��;���JҒ�P�\�;Y�ﵭ-ⷡ��h�h�-yMt�҅����`%��v����=+��썫U^����n�Ğ'��F,����]���S��Hhw~ݤM
fB�ɞxz���o���!���pgrsW{Z�0���%������_�3���ٳ�8Wt'oӭ�tƴ��Wx��=�{[D�I�~w��l���F��f^N��x͢D�c.���(���B���K�ZMZ2���xUѣOl}�/^�T;#��O�t[7�����l�#����Z�X
Ԭ�k��0�/�6����ܬ���� U�e��o�0��X�����@�XӖ����M��E	�kx߆��}#�&r�ӣ������0/ס�7HS|�`j��%E�C-xIm��X�����QIk�ph�4�k/7�ѽ\�+[K*��&�13ae�0���
�
� �RB8���F�(������}�+�<�������+�����h��e�& :bV&�iW��;��BsP�>+��6�G�لz����n�y3��n/	�
��V���F��mHs���&��N�_ Mn��l�w���k�r�F�O�v-���ia􃛟O �UW�0�Q�?�\�ە��z
ۖ�2�����K���YY&��� ������	�#N�(�S(w#`�����&T,֩��c�Y�)��zs_pB���U<Ԩt
M=�(�\5h�=z���Qj5��9�=|�I��_8�f�Y�6�,Vw�)Q6qak�ǰ=�,H���}U n�̼�៽���$l��b�d�C9p)��PIz:T��:�<�V�=<`����J��l�v=K1�dѡ���X���p�v���L?8�R��˓�B��A=upRV����/h�Kl{ic;�q�Z��"gݏ�$�ڡZ8q��
u#+��#g`�^�,ǔ!Ƕ
��WB�V�Q�e����NTcۦ"go�e`]N�(<�+X�INY����ny�۠�Cd�R�cF?G����������$>��<;s^�xyF`���n����F��+�6��w�9�����c=��#k�b=0A��p��H��f���]۶�f����lԅ��E��������&��ah��s������@��e��z���x5cz���t�-�
3�v�|�\�U��{�m[dfxYp�C�Bɰ���^AՇ@`��;��3�ԏ]����j?�l����f�I_9��Uq��8��Z+��Q��A�K����lj���P �ˁ勶���iy�s��5�NYw8���c×tl%��V�A\�<E o|��%���'�E�֕�{[5h�����_En�jέŇf+�ID��#J�0\_�䱒��d�3�L�$m����mhɄ��naɀ�A�������9r���nt� �vekFv�R5.<�i�|(�"x�U�h�襁Ù�Z�h�����}x��IZq��w�D��j�K:�I�'%�����
�ofƙ#�uZ��� ���+�jW���k�Ǉ7,�c��n��0��r��3FK�V{|��P���L�sCňt�-=��	./V;2c��^��->L��߳<AJ����gaƑ��ח�8�*�_Z�X$��ý�~e��]Q*��t��-�<�d�������:�ϢA�m��
?Ξš�.�:Uoc�n=�	��rf��Z��$�1o�~W��i�O4�h�-�-䭞=#f1�s��0�%iC`h.ɲ����^�h+2�Ķ�\���%���@�'����D���9�J�+�p��b�J�xf�16��ӦN��(��g}W�=TE1�z�4@��� �A�p���L�V�aZA��}��wG��Ȭ�M�~[g(�"-~$�0��V���р�R>�M�&,!��H�CB�d?7�����b�o�=s.q�e��4r�s�J��= r��t�A��*�rt���1��1�$��d<d����L�q��}v��#ˠI[� ������p�!1[]�X}��Ii�H	��@b�Y+�S��l1l$bD\#�@S���")�zS@���|r�{(m>L<�����\ۀQa#��'���^G��S�EQ&\�@VO���$㙕J��������&�w�/��ko%���(�9F-r�������UQ��l�(w�Ӽf?�*�P�Ec'�3:(�A�yb2y_�2���uI5�m�&�%k�_|�����-ya�򏲰���Y����>�VE���Iww�؇	�\�V������C��.D���R��2897,��z�~����e��bhZ�_�4b�4o\��.�%�?k�����rd���1E:��j"���O샔B�ux��jj�d@�S1!X)x֝�X�ρ�%�n�������P�Bg/��^˟�5�(�Cf��%,77���&P�z�5E���[)$��dm��" c �/,`�/����+;c ~� -��~g�F�L�>��f_6˭M'u��Ps|G�Q���h�������x���X�T����;��Gm$׃J�*��Mwݬ��D����\�j�U�����=�"����J@!Ap�a�N"v� .@r�s^���	�X���hzV�j r	\��˄�H�Z�C4�(lu�r����UO��������l��9>�o�����ꦷ|F�ֻoJΟl@�:�I�M�/#	]v�J��Xu��\Ȉ�l�����~�.B���ۗ��r9b�)p4�6v�O_Fm]zi6����	�!7�����0�{�E_ա�$:��0���R^L�=7����Ŕ�����a_[���7��s�8g(e�.>i�/1}c�2�L!��� e�[���y�ҁoo���n}٬�q2��>��	���*�CB�?jJP����mn/xͩ�>PTi�;E�P`�*ӓ/*��1:2T��m�!��'�����֪��$�H�>_�Ud�F�J��̎T�iO��Gi�uܮ���O�x^e��ͦ�yA�*QrL�/v�07���\6��!`����KI����Km�jm�ĒY������UM�ա6��[�l���4�'K��
��ɹ ���LT���ζ�*ny_+^�b7?	���*��D���r�d4�P~��n������K�'T�G��bC|b�E�j48��R 6(��"xTB-�,����.3���5P:�X4/6Z��j�-=?����
��Է�d��o1S�W���[�T(J'����&��s�!3n���g�!��@_�=~������SЬ�����g���#�jg���C��h��*]|+����<���?��\d^�6e�X̸�/�L���KIk��ș��FWڋ��>������l�諛������t-n�:2!���k��T/k���OR���h��[���_��W퐁$Ul���:e#X�l�7�#!T�U��B�%�W���=�(���c�d�ҍ�f݁}C��== ���� ��f!�7���X?u��>3�ST�n��GO�����xʰD�nV��q[��
ۉ)'BLK��Zp}m]��A�E����B;-`zu�}��C�a n'�'u;�2�-�׹��?��:8�9[a<�A��KJC���H�EGETol計�9^��߿�ᔼ-4�A�v!æY9��]fx`k[1ʻ�|�LVM>D�ѿ�a��O?� *@��bN_\�]��@o�hp��@B2� �3&Cc)�إ�1�U��u�g�z�|ơ�9��bq$��љ�����i9ZR�b?�N��iQw	�VƄ�ԳEfύL(���s�y ���T:��)�ƞ��c�p;.<��6�pk�Z�,����Nw <A$ܕ8�J��c��jS -=�9�X� Ň�
M�ÿi)~�BQ���4ޓq��^���g�I�>�?�Xm�E�U�uI�gW� {����)��P���}m�CQ� OP��6� J��ɏ���ɫ��m�����b�����s�� ۖ#�,��R�@0̟�o�0�[tC@d��Վ�ft���]Av�N �}�۔����Kt�	D�O�>�Gqd��٘>�>�LV(��S���@���?F@5r����8
�߽��2=��y��p)�C>� ��!�6;�����H2���ǽbֻSe0��j���	6��վj��U����;��Xn!���-č�����Ǥ�¬��U�ڷ��w|01;N6����F_������knf��A�%���J�88�����U��Jq>¬R������;����>Ⱦ�Xi���̣��`����CLjE4~VF�ʇ�c�_myi`�X��2�%ҳ&��v����#�����-�����rDKa�=rNE�:񮺅`�(S���F���{1?d^��ol�1��׷��T����kaS��]��'�T68^�^����hZm=\>Z��`4���K�	a����$g��Z�g�"����u���xpG���A��7'9t\�r�Rc �ڡj�U2<�
��<�o�:$��}.HԼ4/ʢ��]ӽ+OO]�.�gr$o�M��+��m�F� �:������D�����
�%�D���t����Ѿ�-E�:����;=����U,8�sw��X�H
-e���� �3�M7p�/�5��^_��{�6�nm�O�	ң��Yd6a8#*���|�2�\zX,�ۼE�I̶x��p����L��i����Ek�ߖG	7ξ�a^���)t��V>U���bbW��S��q��|2�-�C��k�Rr�=��<0�f����޼� 1ObAӀ�%� u0N`P��s����pBLP�s|���پ誑?f��1ї��� Z��s(��Z��@8�vmۼYC���;1����ĉZ�i��f�/>�o��wL�R�>���v>$�qۢ'םa���C�xOP����Xj1�0�3�u��Bl����	�i��_G���>�W��"Jn��(���ðA����"ʆ�i�8��oP�S9��;3��3c!N�r<:"���e˰v��������{)Î��	dq�$e]�1��=B�����:3��g ����������Y�?��'Ԧ�X���p>,�h/s�@:Ȃ��fyPH&�+�k�w�=cY��,��6w��d~ԙ��N(�(&�-�x��s�22����n+yhO�*���*؍�k�R���R�(Z�AS�������x��J\��="%�X�_��
I����K��:�b��NT9�%�.��Q�^�R����/��]�{x�V�� �ŞAw(��$���HTt�&L�ʲ"��k�{��f]�(�]�����v�Cٕπ��{�^
BF2%ܣ>�mu���vE�@�Ӟ�л���'<��[��F�΄��~h�u�-�ļ�����3W��&x�������ʏPUyEx 6/AI@�8����5�Y��8$���u��#���1����#�.^o]���M�����Y�?����)<����+��mH��E�u�J�e��z6M��\����7�4���&+��-� ś�$2�̓�;E�Y)����2L��p��d�t���,Vc��9t���)�����Qy)�Y\y�W�+�4Q��:��#OEZE�~0���fi������M���K>�/�֞tg��E�->h����U&��Q�J������T.�o�v2hTO%a�э���͠yg���Q^�u�j�g��R�=^]ݽ�W�U��������-�ŉ����?�����@�
�R����`\�.�B=6�A=���;���q�ZV8{�J���ߦkNV�q��A8*ݹ)�P]q���j�鬗{�����Gi��� +߄N�-gܚ�~���ױ!Hb��%�t���:��~����X"�GV%�:��+5��fu�R�*�h
��Eb�`^�	��>�|C}W�b^?�N"M! 4tR)���8Q+�gF��+-�,fw	u+~�%H���x�Z�1H���Ff4�#kiB��!z�Q���+?q6>g6K�y����1���J`���R��iZ�{�B�9�l��ie�:���T0kXő�LJ�*V��̲�%�:/�	0]}�� <��&to��W�q�4��,�*��q�Q˨���+���lB$� �ǲC]�qDd]���R���5~Q�I��(�I����6P·�p�;\��������0T�$��]�x����򩌏��j[d��� ��ö����GH�����`1Ɲe�5��mEaUf'�^�������M[m*�e�W�� ����z�>USN��iJ��P$A�����೗T?z��
��2
T��^8��;�G��C�ϼ���}��\�"`����0���������I��*���0Op�j�\/'���bV{\��ׯ���TMNtv�P1��a�}�m���V�.��&�s ���].]��G2���#�Ak�9���C�;�z��`\�=_:eqJ�"��CeXOFҽ�� ��TWq5?��Xe�W��D��]{�z3F6>(E	ץ���k�;P4��uԬ��K��'�P[Kh�;zԓ?��>\:{��ft��ꌾ�2;t�MNރ
�=�����oG�rO��"�t@&��?"8�/�3���>�\��5d�-LN`�=FX���0�V��@s.���k
��Æ>󡍳q� h���D�?)Z���f�^X�jq����J�j3ꉭ��}|?)}��N?���Z~��Xv%K{�=R�J��z�껙X������Zm];�ٮ:�Ö��g	���15�����=x��^�ɊM2�^x��a�(k�#�cn� A�������g�I��h�/n�`����%Z4{��Ǣ�'i׈ 65hw%�g����K;J�(;��E��H��6��]�^���A7�$ٲ�[��ť���x$CR�r��\����hOD�I� �}�qԾ�%r?Ç�X~D�V��'�i#E���f�d�M�~��	og�G�/||��m�PM&�<u��F��("v�� ��F��0��m�s��&F��K�	��2�ZW�Km9����lx���:ܳep�D3AZ��sm���I��sF��@���.���U�2��W�>]j�ɳ�$�1|q�f�$���x=������/��@���
lW&���]����C�&�ľ�0z�ڌ��u�~�q������F�l9��ə���WI"!w!�@h�s~�7~�am�!c�׭��rT�ЎbÖ��X6$(il���������`�hC��ͯPo�����Pt����������:h��O���su�gb�?ݴk�[(:)!�e$P��[Ȩ�V��WS�K9��O;,�~ǡ|�!�����zH�c�I�*'S�@s��zs��v.�V�}Ǧ)������%=�o�mb�TK��T_;��5@}�v�^v�D���wt���d��20u�>�<�+�uGm:jF�P�qjjl���>p�=�)�y,�'�'E�1_V1��9�S��q�7Co�k88L3� �gQJ�$���c"��FH�M�p�e�!
�����1��j����1�w� s�N��T	���J� �0�F�M}3ϙ��"n��gP�D�p=>�m�ڐɶH�)��l`y����ܮ{a�"��"�-M=�@.n�r��h>P����9UwO�N.G����(�:E|7 Mȥ��LH`b�D���a��G�sS��v��1fD�����
����}fZ��2��1+��]�S#����d��_��}LI�}��"��x�� �2A\��"F�f��K�U��ha�]N�����bY���F����g������P�-[34��,(%�3S�Ƿ��t:����v�`3��I����+]1�i�^]m�������:�K[02�����'�-�X,�w*����w뗟��)�����H�e�@�*�Y�� �"�A����G.T����73��=�UVeW��� \:�(yϋ����8���tH��+�oA%�n ��=��s�5�����y\��.x+�4;�Ƥ䩎��Z>�)�d��4f$�xF���4���_}�zI�𡢓�Ő2
�Dnf�?O��.��.m~lw���Bik~{���|�^1���
���3���E���,�A�rV?hU�ɍ�d��
�rrY�ņ1� ��[�M=�\ ���Ӓ���e�Q��R&�T��A|�JY�<`�Q S\�p?�	�f��>+����[��F�Y���1������qU�I�>4u�y�ܬ�1��?ƘEZǲfD����I��'!<���TT�� �
a����d6��Zc|���H��
ڐ��
.�i�|�$�mS��w\M�C�2Hx�Og��g�o����i���*U��T�oN��D�*�i���T��Y~&4[���l���8ӳB��#��LMzUaI��i�P������Ш�e�������T�w�d�-��gթ�]�ƣ��x�:���(���`�QD@�rd⠁�g������?�����ٵ�b�HɭT��At��:{�8wN,��7_��]�o�߁`2љ��I�Q�x3ԙ�������F�
�=�mWz>UeZ���G�(J@��A>�S@.���ػ��㺵���0�d6��,o�}0���0R��h�F^�2�蔶mm"�;9�1K=��M��wC	8���i0$y��8�M<��ߝ�9��_:����-��)�������䋄��������Q�}�_}^���#ЂR�F-JN(^J D��%LN#���gԩ�o)H-n:C�$<�j��rP�oiOlю����!�e�d�uw����fW�u�ǻA�Y���GSM��Xx�e����.9���?�1�K,"fs�o�Gk�D�$��l���}i|4�iP1�F��ڊ�b�6�^��"���̈z	x�SR�_��v�>��7F3���+x�La�{>p���X���.!�!���b�����q�3��D ď�
^:,J��>l�w���T\�^\ޓ[%Sb!S��̧�
�Y����B�N�w�Qt�vOǠ�:��Zys8+�"�аo>���=��*7����S��SȠ̈́ �L����(1š�v!�Q���\����bG��WP%dѣ�Wq��b����y*�lZS��r�>��$0���h�R�w�����b�L����#�_�N�nM̱j�(�pl�oD���.�y,+~Gt5�w��$���7cw���L�����`_��?O�ݪ����*m�m��;�S+�si���(���A�p+K���k�|iГ�Kd��rކ�,���W�-R��!�D)�{n�{wO+:�GD��y�Z��^n���3h���=|:kް�+�5��<����o������؝�;��z��R�\����6�җ�`�E��L{rSj�
q��+tI��I���j��	R�g���F7`a��P6S��3�� Oqn�&Q�?P����5>�T���6��6�FHFܱe*B�gp=��}G%�}�㲻�ף�2�Hv���m��A�I��n#�~��ǣ~��2���Qլ2	� 8��&�mmse�C�5�H�#�ވ',=���/.�Pq4w�������gL:Uk&����eH�Qj��uT],�7�~�8*f����m PE���5�ɫ�|� Y��]}��zx~o��eʚ��"3=�o�FS��=Fq ׮��|�=��}T#8>E�b`�/o��H������m���?�ߍ,F��D�яn���%#��xدB�9c섦��N�x��I �F>�[�}$BYfZ*zx��Zd�H�ہ9�ط�^�c����[	u���� �D��M����_@�+p�,�[u)�˭�a�h�@O"
�-�݁,DY�ʬLE�/_4w�5=U��<��]����Cӂ���b�� �?Kgh*_����_In,��`�2d��6�<Q�i��ϩ+�3��c��Yo.�@�:_�U@S�oE���"Hۂ��2���,=�
 �4�'"q���t!�}�Z��	��sҀΖ\���hS,�4身
�}ٽ�,�\֥��.�����\���?��H�$�<h�6�r��x�O�d!�Dq�͡�g������qr�u@��B@Ff��.<6�axEve�����ݼHt��>��Mn�Y�̰ɱA�9>��H��`�{�cV����-�����ޏ7N�o��h!��}��b�'�$����L��ݰ-��zk�����;�3�U^���w���7.S�
e�p`K�����5i�&'��}���[�ˋ����"�s�I��A�̛�gk$��)��?+.l� �"4ˮ��X�J�χ�#��x﹐��[`Ȱwů��J ;���]8�q���Y\�qml�=2�c�J��Y
���Z�1/:�S ���Gk�V�8�"9<޻F_�V��N��c�c�]c, 4��D��#��9m����/g�We�(J�����=Y#���N�D�H���/��!�z�.����O�1�8�^0�o:E��?�%>,��%��#�:��\h3s����|��ł��}����ԃYڎ���)�$��l�Ԯ�A�O�%u��c����JG�צ�O�E:66:���d���%�y�w�Ih��xl�y|a+4�D�=����L�����<o
6O�W|7M�q��R�7�+�ڗ��
��y���_�H��|�Ȁ���&_%	:-ٙ̵:���1��n(��m����n| ��Y�|ڑn���3y�Byz�SFW�M���CPG�s��4����T\��.n�[_�Q���@JQ:������z��,I�,)�@6���oѺU�z��-z2�J�����4�sQ�_G�<*Lʧ��k�L�4\
/:J��
y��h��o�ׄ^9i��5Cm��3�.@��?|�#��
2���6@M`������q��@�6�m܌���Ś>J%��1��R���ԟ0j�z��:k��~m�6s�4�r�P5<���^2��=q��1@<��+J���GQho�sww���bFz=^�}ϰ�'��q�������N��&���@�Y%apQ���g�P�]=�:1@Dϫk����q#4�\�0�o:�)��&�QB�ڹjz�͍is�RK��S�"�ܹ�a��\,b��݀��r�)�4��I{VD�ԡܗ�G&�ON��F��
b��B��6�ό��j$һ������qxD��r	T�Y�Ù1�u䉇�����t�nt;�a���ws[��H���@�y&�������+$lk8<�Է�c��.q�G��K�vc�( j�?��A+�X%��rh��Q�{'Q	��T��z��̿^EP�z�qm�UBT�x�ۨw:\���N�����`HZ�N�	�?�F��X�N����
!J�6d�J�	1$�c�؂=��7�]����91���J b˰Q^0K����y17v;�r�e�
��݃�1�ZV���@)����pzF>�J�u�����)� l(��t��W߼+�P��J3��8�!-�iX�Y�xi�n�C��r�,Le2���H'(�&���y���ݑg����� p��sh��妈Nf
eDl+�݈%�������'j�/�i���er 옛ՠ&�6��?}�d���}ʆ!�����J�di%#��1��'�:�>���8�y��������8���B;�t�wO´��\$�ÅK��K��n^۠d�q�x4P kA����|T i����9����+�����>�h:�W)��3*S�.ڥ8�Q�͌۲9k�s��Gt�4�-l�j��A�΀7�Y�k(�@���p���sTpU�L4.��B7uU���!ztAJ��h)E��8�{��[��X'���骃N'�>�~�|'#�dk4��s��5�J`?T��ݫ]/�ǝ��!o�P�4�OT�%ղ��N�#�AJ=��bO�1�m�O���(�9����Uw�P�MYP��N�7c(=f�� �8�9�(l��*A��紱�G�_�W��TG�-�x�щ�fp�`����I�_��ﮣk�����K�D��L�0Z?��܁���8��!E�b�_r�V{Jҝ�.�mC	�8V��8-�3�Ő�i-N�W�:.�^YdB����'��N	W$��/���,{v	ɻ8}���2�3n��:X�zt'�A�z2������B�3����򊋥�<O�Y�-��Z`l�Ө��z��8 �P���)95�q?*<l  ���;H�i l�VF؜�^���Eygi�߫r#��5>��ͳ�{�����{a�]��"Ř�j�iM�n�I�����M�N����m�V��C�Z�u���ȗ�+E*Lnk/8i;ʐaC�;8���iU�E�+�&��Nq�rA7����2����Qa��`�"��iѨYsG��+��e.<�%9<yK��<���/�g}�%׶U�t!&�
Y�H��Ғ?���>�`�~.�������F�_�!�o�|?�/���v�lK���w��w�X$J��eႱG��H�\�d:7D���9Ki�d��6b5Pm���:/����1ni8w��a�=��:��h���N��Pp0�h�	�֘�gV��	<��]K�o�!�Ŷ��v�T���#���K�&����Y�ȿ�R�!;y)����*>�v��hA(<bP;fU����g#�E������ΑJn����4{A�ȱfF�������N�h��c����y��<-\I'�h4=%hԩtWF5�L�0�����;ԓ���z��6��}�0k��*^]�~'��Cl���'f���,^���׾߽�z>e���:�ܝ�Ό}�2��T>]{�l����iC��9��3j a��ʠ��Q�㿓��?T���o�����簚l'x=�S:�`�u	��/魀���5=�eK�
�_W�#o;^���D ��+��gjRQ���]���F�W�d�,'�l��G�{܀Y�>.e߀ZNq'8>A=�����Vi��G
e���7l ���GBM�N�ؽ�V��4�)������dYc�9�DJ�J�>	fi�ܒ�ί��#�}��X��w�%��\��s ��:��a:����鄼��$�'�=$��ܙu�ޕ�{9�V8g�%])I�B��t�������3��~������խh&/Rl��v����[�����9H@�ЍFn�L ᐌ�Eћ��ĕV_-��e���e�U��ڟ��Q�.�I���!%�e���ʢ�k�D�9E���6c�S�Y�=��=�b�.��*���28<���WWw
����WqgG�a��q\�M���Ȫ��@���á1�b5w����:�ܐA ��LD���u\��j�з��GỬ�
�H�+�A�Wp�t�.��PFW`�h�HB%���O/�*��	�o9�Zz�����o��"��8�0%C-W���'��N�u-���=���U�B �	r��Z�H�h�[�#z�~��`��ڙr�dp�f�En��_�4Y���VM|�;4qU�`%����Gg���@α<�i�Q��PK��g��F�lx������(md�@�{�D�޿��I����!��p�2���!�n�ΰ�����!Z��찯����0gi-U��
�\�(�L�19I��A�����3�ߏi��&O���ֿۄP\�~.�g�qQ;����Y
ά���x��אn���pA�y�y?�3P�������n⯓~ |��n��0��	>�����yF�<s�b�u�eA�"�)DC���t1�	u��ɷ���|�W3
��O����9�'�$T(��j�
��t5�7�(���+�?�3�Z��ڇ��S�,��[� ������+����'�n����M��0��tǽ���C�{Iz���ɗd��a�>$7O۩7�a6� �N����f�[���sR�9z³�|�^1��"� Kx����_Z�$҇��H����!Z�����Tfm!�h�q%Sq���a0��`G�+��g]VR�?d�?D(8�c裒Jd!X-�D��Q9'��A�@��_�<��B�fT���
���̸[��}�[VD9��c�l��'�#�5b�E�l�A��`��}�Z���_����k$��R��A�����Y��~�&
Vª�(܉�����@��t�6:��7�z%�r��c�7�����W��R���>oT>�wn���TZ�#v���?oL)��8��5n�W�-W��|{�	p4��G��u��9�Wi�×U.d�Z\Y�痆�Z^ο<��� �_׊s��Ѵ<�x����r���G���/���	�8q���j]�»KM·�-��8#�� �/�*���T�%���!��|�!���<�b�i� *!�,ԋ�~a�L���s�O�EU*�B�X+ߕ�x|g���.3�N!Z��T���$d��=�&�7�,��C4n�C�A��k�G�ȗ����{)��$%��4Y���!OX����oႯ�&<�%_m��ôՋȎ�|��wr�y�#�/h�g�d5e�,l,T����$OI��m��:9��-f�O�~R,�!H�8g�b�{ΎUCb��m��
u%�y�����8#�z�tG���𹍾��<[�U�=��R��D0Ĳ�
5_�3� ��j��6�ѭ�V���ͫatg%��O"��v�+t��O�g@�M�W #g�kV�W��r��-/�^/�-eQ�j�X�k]�Ӊ&��`~�&��C"��oj� �x`S�ݻ����/H�20����V}v�7�Mo�[jY�5T��HN氬��5_e�G�Ӳ��K��2�ߘ�|���C?�j?����}d1M��$����{��&�XjN5+�R�G�8E�%@G��) Hh�ӻCBض���g�S[����;~�Ձ�i-��T��FP����>��@�� �WCf��כ�MM4�_��5Z'粒3y-^�Dr%�1���x�%�_GӑҘ�h|˩x��5�&q��=߰��D��Vs)t_��
��Z1OpG�(<� ���\��{==_��#0�im�v	�]�x�e|�WA&ĩ!��N���(k�C}�l�Xr�d�*����4���엛/�l6�����i9&�;8� �" /g�p��ޜ$���C뎡����$�c��P)ޕ�wa������A���mOD�t;���涋5�����.�F/6��^i��`^CfCC$��L��Q��'�K ����))�Ҭ��.`��shL1�A
���u���r[��=�%�ic�?����ֵ�'�`n/�Z*;q��Q��#�ֳO��nb,D��艚�	B9�tW�O~����V�w ����(%����A<�Y�X��؟�'�������,�y/�T��0��@�:�N��DE��F!̋sC�b����ݎ?�RJh����Ô	g�p����+�'��.}��Q[i��a'��		��*땙�;��͘�;8!�����Ż6:%�+٨���׸�6'��+IQ���!�R6Xn����#A�8�/��e�@K���9}���jx����>)
�x��CxXƺ���y���O��M	�g���캀����h%ۺp��q�|��6'V�8}�P�o�@�5�d;��%A�'����9��Q������YrD�+�;����h&�56�}��I�M#�KK?�
$@g���Q�z�*�⑌(�GȌ�=��J�_�Ѹ�� �`Z$L���҇b�P�2�)ƫ�)��6t
������m��g;�#�D���@!�crh�u{��~��A$�n�7̰Ɖ^qC�_c`w���*��_9�)Q�j�i��W����E���QC�%�����T9��Q���u��S��,������R�n3:��Y��*�9����·��)��،O̊��7���1s�@b�︍x�2]�F�KhVD32���4cc�'}i��Y�
n��B���ԏ���3}=��u�q�yܧ���1i�G�z^�^��Ev�t��I�y޸�u��C�B.u4�&��v���.		��_H~u��p����y�b�_��Z
&���I�β@}�l$�A�<�5L��Bc5ޥK��CU�!V���C����;�G{N�:p�2� �݈F~�FPXs]�n˶n��}���B����=�N��JB.Ԥ��#��ߎ�!��3dd�i�x�&�~�>���H��Ģd���PJ�7����@�N����<���-Z;�q�P8��߄���J���-�����A8M�Z�^ڈɼe�ҋv�3������Q�ޕ�5��O'��a�H��jC�+&���B�w��;���Jd��pb�<�<�g�5��p���ݘT��v�E�� ���Fu�9�gǠ7��W�r�@��k��TsGWٜ�lu��X�a��6�TH"���ivLAz���|@ ��bG���Ni�����~����]�$W�� ?�8=�2���Qx��V�@%��\��L踘R�9����nWbG�FrH1���h����"�`�>�0ȴ�{����s)NL���\$S�˷��,���:�.���~v���,��	�݁'-�����=O��ɪ��P:h#��P8�FS�J�A�����:]<�b��,�#�?S�a|f�o�l���8�Ki^Ӛʗ�3f�����Bx��`��oGa�Y�|�2cΙu�\����]$��=k��u�fJ�bխ��B�3m̩jq,�$�W�!�Df]L�a��y�0��H�kiJ��!hm�P e��dY�V�
����������B1�jp6
��6]J�D�"�+�X���O7�z�v;����'C�Xhyǽ>{��7��7���H��v9�VȫL�_G�?�������	��_�BU� �,�SSݜ�@әȍ:0���)�B.�>�Qܻ���FCs5��Q��K�N��ST|.3���X���;�o ݅6_��_,���1��˞:��2=BF|<7?�B-sb�*�V�@}0�H9������ �����0�Nd������q #���5#���G��J���f�� �"P
{�w�@�y�%/t�$��r6(y_�`����yJ��MA{�=vW�����G����B��վ��G�sJi��O���A�KF�Z��e�#�H>�_�ueZ0DN�k.���hK���i��+�1Y��`�v��GO������	��(�'A���^��;��ݮ{Q'y��?Y�G�^ݞG���2V���Q����
�T.7��!�CAv��A_�>]�Uq$ރms�l)pJ�g*-m�Sg�b�3{+nP�~����]i����$�tq=k2Y`=���������6B���C��@�~���S���,��{�ި�#O<�k����~�1���e
ǤV+�1���s�i YQ��B��ȅCg��I%��%�Fô��^kwV��]paӏ��myv�7u9��,��(ⱳ���u�V��������v��%J͌U6��4��Q��y�pw�㛫@��g�H��J5w��;/^�X��r��{�R~�.-ط��6�4�W�\���~^����O�yl�@�5lG	�9��v������w��g��78^�s�iMz�O~����ZɰI��ދR�o�ޮj.<6��n��#�<�1�vRg�R翋�.��wpʮrH���{%d�#��D�\R'�c㌠����z �tz� |{��Ȭ�������H�SM:��	.��$t�n�(���3�	�J�����~���6jR��� rS���hG�<B6!���0~�5a�t�k�FKU
P���@��2?`�~cɧ$~�����'$A�M� +�D#�Ny�>r�!�� �OB�O��Acpr��fɆ)�<�JmX��{�S����SX�0Z}�w�W��ISkێ�������mk{2��/GyBh��>��u�bb�y��.&��=SwvWв�&�5F�I`�2D}��g֊�c=�`13�i��C��3Bk�[����.o���c�U�k9�L��-V�E�cKLB��)
(9\1�<Q�)=���_s�?a�&K5`,�xyT��\�$�v�ffw��`��tP���OL�#{�ez\���_������˾�R�wǦ�e��-/�;l���x؍I�m���+�W@��ޮ���SȾ�)QJ֚��r��H�����M��y&�`�yX�s���e�ϸ�V��F�+5��݃�Ȣf؃u�v��<R,��#,M���5I�jć�F�O�􈂂ݬ���������]^�X�O۰���S����z4�08�}�#�����h��j�b|�X���**�Gd����}B�g����lMy��d���ˏP�pq.d��{)[6iOSW�E{k��D�����,������!B�����ܔ+5W�Nr�kD�O͚k�hb�C.�i��x�o�o���U���k��x'}�\�,a%3`�(A�T�g�J^���d����J:�/����'�Ю΀F�9c�}MτQ��2FOf����W�ݞ?$K��jD{�,�'�~����2���zjW��y�����If�ݢƱ�U畻E��瘽1E2f�	�p����px\Yxs���mF,�z�+E�Wī-3����-����ue�^z��,�3J� �X��y_H�U��K�Xb��:�����2�b�>oe]���A��ܚ��k�2��9426��j�p��D��[�aj���cY-_Rc����B=���T�ȥ��c�oݚS�6^�g��$*�(�	y���`.���K���őC4��I.Z�J�߭�m��� ��ix��B�q��P��nP�m�Y'���|o#��$וX蠟�ZW�Ho��h��\6QS��"lW��ɤ�'}�2��3I�Eg������z����#���!D�F]�G	�?ej���� �1�A	�o{�@|cl=E�o1����:<�-5F����(f`���.�ȡCj�dg����^%e��?8����G�]g|�t7)�ׄ�Caq�=,jT�8aF�~D��A���@d�'�w�%���@%�S�����'��}.,@�4�x�!�Ȯ�U<�5�p�]�ȝ��J��(w<�5���k��~�A�{�7�Q�X�IN�g�]٭�4j!���۞[���M4t�[�'�sObϡje�p/J<�}�˅�X46���b���j�%�.�l�q�+�ʆ��9r�yU�V�m���������䖰AQҌ��h�*��� A�P:�Ņۑ�c�3-�QG��P�Ƕ�o��.FBo܋���������
`O��6Z���D7Z�2^X��]��P=r����[��U[��\�x38�����G�ن.GD�i���"�F�N��/������Sz�
�7��jN��������)ge�oI�i����=��.fE�\�h��S���U�@
pn��Lj��Q�zM\> ��{�Eq2�s���0@�_���l�1rkt�cH������$�����]�/�
��u����e.�H��qi¹v~ú�nv9���Z��c�ف���N)bG���`g��6�~"�Ō��)��m}�&R��h;H��"G#�VN�Chq�i���2�P*�[Ly�x�K��%���<���dF�G��)�#��l��(�$��/�X�;m��!���w���O�����Į/�ү�+����h4���f�=��� �oʾ�:�co^�.aO�iN�N��3���؈v��𛆐��ض����ʣr�u���;?�<��{5������ f���/_���Il�MpD�	]�4�[�{N��O������5C�K��^9�m�ڜ����f%��fq;���~'5�2[��t�Ά�=�����M����h0!�����UN�@R3{�fU�9���
�^��n8գdA��WX�r�J
��`���G�F ��|�-���>^�3R����j`�߇��TX�U��y?dYgB9�+<��\�e��2�X��/��{�J��� ?���V����1ѰH�Efb��~UŚ�>~�-8��z@h�L��xk �d�Y�ܽ$_΀fRA��8��˘!��2]֩������Ҥ�����}�H��eq�a�#g�P]N4�Sp)��
�h�:.��}�	���a�G ĥ|���nca|�~D��i�WW�?qV�M�]�,'Nnw� ����*���D���JN�v��mnuLSw���Ey�U�(1�5�Z���?NG��OX�Xtn��u�kWX~��Md|{���
��{�T�Xj%�YQ���)��{C��>�NSۊ�P�:D�����q��/\�Τk�Lr��u|�3O.�I�-����� �j{οRfQ�$:2Y�R�1������3L�Gf�O΂�)p��)��qX��PgEߢ���P���^/1��B%(�?�k�_W��K5�6|��XW��D+�z;��8�hw�
q�q�Q���7X��\&�)�ǥ�w�a��҇���ҟ����I�Nfi�O�����t���l�;�_���٣�a�r$Y����� ��QM���溰� |d���W�Y<!9�߯�-N6���!Ɗk�h�X�����GR�p��-�)u��(��m��B�i.�����,�$x$�6�g�g�����od��Ȑ���V7KK��W�їp�����Wk�
�X�\����'|�;����h&�Ґg��y<�Sޏ���S&/��ɾ�cާia��إ�n��8�����v��0ag߷pR�T2"�Y�\�-9����G�bbK���x9L7������Td�l~�G�t��M ^=�Yh��xW$��'�tsm.��R�����[;<�,���%��sӨ�W�Iʋ����	�K�����aSA�����V�1��f�`fk9ˑ+N=o��E�rT��f���8��:��I�K*���p�i�\��iH�#�������Vu�X?��TʙZ�]v��N}�&Vΰ��,+��Ƥ��vu�2�Э;�S����0=���)��~�^�� �Y�:�����vomiȬs�������)Bg�r�DO�J:�u��I�(�E?x5"{�U\��w(���D����_�bq.[��#��k���#?�G�d�Z��Y��in)��p�w�/sXx�V�i����4�H�� �v��S���M���-�!�S���g�IAܘx��-h� 58/7�Q"<����f���&$ȍAJ��&��|#�)�c�~of���m2RɃ�wgZ�D�i�z3�^Q������_AC� ё��&�{���܃���rcρ:=���(`Z�P���:[L����]���z��(f;�_�����UD�2���s��6yE;��
�|�/��(BV�O���椖��O���:����aN��n�����*���Ng#0�/!�R���ۺp{&]��SB<�s3_���b�dY�J�����`�|ؿ؎?�4,1��!�z#t7`l����<t�K�,��QK%��, Z����r#>�F�����/� ipQ����kMq0��n1�'H��P���㜘Y����@��a]`$�9�X�h�"�_�e(�Dƿ�L�ǿ��0p�n�wa�vfTgy%�k���"@��X�BMe[�Z�8���A��� �K�K{+�~�����I��*�C�C�U��ޘ�Z�8YEW�t��o�0ǹ@�Pc�fs�<�#�A�ۅ_��BY�G�JS��/�=k?��r���-9��(9W �����~��d�����Ⱥ������_.�_�-'�w�_L���ZfG7+[��Ԏ�z%�ҧ�g!��6�<�.rO:�z \��UI��/�i��5N��t���q�[C��ˢ�U#��U	��:o������k~u�w�y��H�BFŏ_<�-*�!���`��4C��1#m����W�_8��!F3�A�fPy@�>���;u�v��)zM��#�Oo��4Q�ŬF4x��5P�*	-.�Co��[�}�E:U(<�g�R������G
�O.�5_ȡ�m��(�*��f�b��$. ���=�r�i�F�Z��S8�tN�h���q/hXý�cF��Dd�!��p��|����Y��<b���=;��C ?m�z�" �<��2��n�oʯd�Z*e�Z%�#GVs�E�:Hh㭯�fK�x�E��c1�e�hw��s�Iy�M ���=��_��T:~��.9��[�6���[P��lv�$�5������"6n}V��r�(�t��V;�����K�\�����`�G6�vcEpQ�z�����O�4O�$����_열z�9?í���c�|�V	�J#t�K��6��SV�����@h�0�3���F�5K��{�g�[qM�Z9m���c�7dD�&�MzO��A6��Y��	,��i��������.�Y�B���� �m/���<Ns�w0��J�7��+;	���'�5�7�x<E��֨bD�E�0%�f9��!�i[������f'+-��L����NHnls©�j�V��]s*�;ĵ�͟Q�B�T+����6�'���d����}G�=N@��`����:�N�Vq0?��p-�����dZ��y �9�略Zŷ{�r��i�\�'�V{����"�{�y]����?/�ŻN���g�UjJO��H@�5(s"(�OQ��� �2�x)�Du����ZsL����p�����d�_H�Are)��"&;��C�x���X ���1����Cn��������
���P�u��J���̨#к��Y�D���]%��zT�*RӾPO���)�}~�j{	Op�T��j��^Oh8R"�	!�%V�t�?n�@��!��/�=�L�'*,��N�$ �H���������[v!8��,�hi��{4�xܮ�#�p�����	L=��n�������2�+a"@�A/O[DM?�G��s�u�r�QB����F����a�����2rh�B4B�{y��!^g�E��olֆ�y]�t<?�x5�XI�?�_�� ��>�Z�ewm^0���+�d{j��*L�����D��X�����Ij��?)�S����tt0��7W���-]�
��y3kO�4(���k���$@O�B˓��/d��	s�����:��E��� �ab"��d��!��y��E�ф��(����iH�lt�wdA���û���C���@��%Y-��m�<P㬱Pӕ������,��{1z��/'�_6�6�p#E�)�o]�XJY���5�	��|�r�PV�]L��W��/h�<틌��Υ��37����/|��Ἀv�7��;.xܶ$i�[Ѓ0���?n65�'b�62{���7��E���
~�{TݜL�r=���ОQ�ޞ�[�9�&���e�[����/'M��"Q���|�5���ʡH�d�v�o>C5����t�XQ'�v��ց�{�2���m�z(�x�j]����.��%k?�>���b���mC@��Tw/^��������jlrMq��Ѷ��G�[fa`������� hnX����t�E+!�r�a%�z_ag������x���=�4�� Q�`B���P������;�k���E�(�e@!�C+Y����IS����Y�2�:'�^.��k���.ήٛ�F�xh0=��3�;�dk���m1��_���1��]R��/�t%�뮗8.gi\S	��n=�}�qO�Bm:	���bg�D������Jx�@�,n������l�/�ZYȲ
��!&;�[!~�Vz�@?��8ugZ�еk�Hh=��\��ܢ�*n-��ڎ��u(��t�K��l��TSvZ�d�X�v^�O��s�_]Y ��̦����s%��.���t
������"���'L�lÍ�m�|�He�X�$����4�$�,�>b4W�lSs!�/�1l�'ࡽ�r���!o_7Ew�&�k��ҋ���.闿���!� Ys��m��oT��i�^�Twu��u�L�Fܻ2��w�s!��~bG�A�\dh蓐�s��#}$�מ�럩ū��+d+]��;�)z*6į:��8��4klg���i�������<Z����}�ּ'�T�m�c�L�(�UefP��e�A�3/Wq�⳼}4��#��_v�<��Ƥ�rSjF������P6��V�[ߗ���&& �|�pV�u��%�ѬEj�?��{�@�-9�Ғo��A6D7ܧS�_mT�,������0S�!��z^Z��Y�O���O"�13v(ǿ���d�1����ͳJcKP�7��_BX���$�%B�6n���44��U������.s���n��^���������9Z�p���r�������1(�1�2|��#��"Y�z�8|�o�Mu�����j��Z�*-8�SD:�m�`���{�k��ɘ����C6�`�9s�o|��F��-+Da}�,�+	�C�ub��&#^>�Ut��E�f�."�*�D��mި�L��%����ó�͆;��hB�����4]�	��م]>#jA-��2�_���ʪ�~�����Bpz�j��"��3^$	��磌4V�ٹ�/��+�-�����BWr�3̈Ś������N+r��}����j�����A-���)k�%��¶��i����gbK��Lm���wiO:��L��������@�0������<���зzC��,Ab��iV+X�G#����;զ�Gl�Kq�R@��b�Ե�p�pl#�>��/sL�r����Ɍш�8)�d��z3������)ʏys��{s���8��nCua]OӸm�5.Fז�tB�߃Rd�N������zz[�햐���K�M�M�xS�K��t=t�.�н��@�@<�
���H�ʔ���nB4%�8�/=�Pg��2�`LV3g2��)ȓP�m��2����Er�6��`d��a�[.�
95�'�ї�Ӟ��ZY�NK�GXJ<��Jk���R��m�}��g㭮��|��۾D���0]�!���8nW�,��o��E��f���=n �)����u���fx+Ya��%3ep�K�/�B���fMH�G���")Mn�!C�%|�M���­j�E��ξz�@Uճ;���oe����%,�Km/7��o@�0)�7�JE7�:7~=�k=vlr~�N'm��М~8�4uL���(�<�	)��&kN?��O��l�z8�������Q{_�Yi�$"�xq�}=�e�y)$��uL7��d�2CÃ��o�迀\\j��\�'kv��4��i�5"A{�B>-��h�I+;3�L�o�1C6�[�/=���L?r�
�8:h���_�JU'7�+��j����Z�h����˔����Y:�:���,_�o�m�D4c]�RMxh���Fsa#]y㠾_'u�#�5�b�Hmlѣ6��6 8�}��M���k�i�f&��T�bu���r�m	��F9-�X��ƽ�$Я��\T��M�b=L|Ζk�5��C���i3�D��V��K`<i�k	��)�2�^z_�O�����d���.�+m�.!��V#�i8l��JNM��%lm���%���)�bDtQ�����6�t��n@LX^�>�����f"�CD��D���Q5�����$G��["�y���y�� o�n�z��$q݆�d队B-��ɭ�R!f��e� f];���iAW�6�z�+��w����!_��6���Y+�~���@P��f�DD�����ܱ����������~vl�F"��Ŗ{B�6�y�Pm}]�J.�Ց�H �}xs �Ȭ�"�Յ.\�Ht#Zs��I�77������f`�;Ϝ(��d������U�8�[�[���a$*�.hɳ�;HBNR��D��g:kt�7E}���3IGY8�i匈Gz�PV��:���hzbi�f��B�r�?
���)�װ����a��ĝi�z����r>�|�����ot#�K4�EL��N*�L����W��A�Y��2Q���w�Z
�՜'U�����ޘ+�|�~��K�$����p��w��_;���ZU'.�>U����C�(ß�t�0D]���x;Eo�Q�[㴗�<��z��U���������n��D��&�>���
'p4���ʶܡ�2:Z���^��,�nܢ�.$�Oo�W�'�,�4��E=h�܇w�!@&wE����%
�
������������ۏ�i��ҵ$���ɦ}�=�`Jb�����v����ʫ����}�S���/�T�̚i���䗼�G�w�?$�4x��l��!�jxI����՘83V�S��ب���ٗ���I�׭��s�P�����G2§�x@fei��A�?jI>��߯a��Pi�_(���:�g1��$O�<�}�fu?����JeU/)��mæw�@����ss�.��J
Uv��0��R?0��`���F~d���-�\1��ÿ�榞�w���%�5x �!���?�q���Lr#ր5�psK�7��`�>�����t/g|q�sQcM��h�n�.�����y g��������QeM,K�B�!���������I��i~S������F}0���C�[�Ɇn���Ӹ�r���,��q�c$U,~���|���A�/���i4Jo�Z�a	�կ�C��DO�>ي�F���`rck6{s����}.#�bjg���
���u�5f�@�PD�f��'��x�Vh�}��q1.��]��(o��+�8����;�\E1)�ro��J����^��W�C�@�J��J�aԝ_�_�L=�̉����ڥTY�ŤԻ��S������)Ԟ���D8��E���,�Hiz��Rw+qќ�^Aٱ{�T�����=����+��uA?#L��6��4�奣!�u�[��$[���L8�,�B�h�:�*�����C>�.�ɂ�6c6@���09O�\��C�:���Fn��]m��*з�|Q�-ьZ��Z؍�bi�_5��`�?�\m����(FÛ�����k-�&��Jk��4���l(d�M�ҡ���F����4�Ђ�>t�����w�G_<ƌ	z�J�L�e�ӺCr���r'����cA^-����Fv^5��}"?W/�,x3^ 4��~�2'�O��"�1����rw� ����"��O[���U,m���5�%qT�'��Y�w�c{F��F
��� x��l8f�������bd���ݠ�1˧ ��D-����ݮ2a��Vd��pK�i���Y2(\9&�Ì(u�೫�V�G3ޡ!!d�M�����6�
��l�0�Ĝ� ��M
K��RXyX�ٱI�I�a��a�39�*D�
�z�|笡��#<|�{� 3е��B�[ �&Dp���_%�D�X�UNk|F�v�X��ȳM�ᦒ�bD9���ύ���fOӃPX�/,{Czzl
f��Z��>+U�3؝e��d�RG�n�(��M���5����ύ��0M���μ����s�4��k�0|���/\��vL�F����*FpC�n�$U���d�M�& �X���p���O��� �ۘ�\/�	OT��<S�$B�1h4��^L-���`�G�y��oC�h��k��ֱcѫ�|ʱ8p��0�5yw�K�� =�.?.��
��z^EC;���9+�(��dg�T�#�1�L���&�6�g��/�� �}k�"��ʗФ/b�5�Lz.���>�$��e	K7��+�����D�ɒ�of�#Kl�Qa5�8�.�$U����l�ڨ�&-�o:�0n�T���_ҧSg(�b/�?�|k�{��`�f�턧�V��!$��������{�T-�,2Z����?���r��^Ը��RY�����)����L׆��#4
�d,�M���EI>�88�PF�������؞��]k�{<S�;�A7VT�GK�l�������J�YN0�z�slB�K���oj��ƅ��e�}�"�s���֭.+z=�)\O偔�}��0�T���`{�Ҡ�H�֦��\�$�BCZѠb99�@N��V�s��3������V�yJ<V�\`�7�z��%U=�J��jU�vtY�?�"����]Z�O�O�3�	5�����^֔��_�|K=��O�{�/�<�f�et��.�W��^��x$8���Q<U�U{uz�w`Ǡo|#����,7V�w6;��5����%�S����o�abN�����7X߮�׬����\�_�:]�(?�b���!~̲֛��h���󠻫�slfĤ�7�Hp�Y�Nդ$���$Hh2\M���i ���OD#���EY��ֱw�?���愯�g��F�̙�p��3#EA�`�"�l��fx7��������߹&8I4���3����?��>�;Ί�;;����Q�R�w�\��5;n���a���� �Q�@�K���`��5H���ޭfGw�K�'���VZ\���}�;##�K�yO�ز��cXi� ]m
4�rd��_�{�2�.�YX��o1d�Im�q��{�����k3�pM���	���?���,���/��'����J�(����M�<eݍ��u��ᄊ�H�5���l��S�b��X�$��n$���;g� ���j�����x�j�o!�ȐpP3$8�"�I��iR���clk��Q��d��"�b�&5� ������gd��f	�+�צ$���?l���x"T	�ۥ��,7e����_E�cS�Z(qMU�)Ѣ�J����90��K�e�ʝn1̩N��e�@ ��.�D5��>=�l9�a�ư���ۜ�dq����v�,�#���'T�Z6���b �1��l�Y4I�P*	��=µ��܉*vAJ/�:���\� |SU<g�yw|�;�q��qPʽ-v�n`8�X���� K¦3\%�'�+q{%�u{8�";e~Q���أ+��>*m*����1_vF�AzW��i�0�]cj��Y0ꇞt�I7E��Xa��T?�����H���6��P��&��ė��X��۪i�E��`4�����}��>�-�+�Rw�ȹgt��EWd�y��a��R��f���B	��7�C����y�v0i��_�@_-�uA���kz�����]NF}q�yT�2��S<��';;�E�/)m��0��ΥQ�� �/�"�($~�$P�;�0A�g%��99c���eXg�-?�B�
��LELiૃW���Va[�}.��YH���9�U`�v�b�+iJ��{1���eR�Vu�~���O�n
��E�m��M�=��,���Զ�B�~p�/���T�����:
����!��R��_�ܕw,H�*�l>yQ�	�k����)a7����I�Q�.�yM���l�1�~�ٍo(M.�	J_ŲL�h��}T�-��i�]�H0�{f�WߘB�YPq���@K�TW�8����Eֵ�S~"/�[����:U-V.Ů��V]����Ŕ����偠�|���#衲?��4�.K��fU��C�E&���M�c���y㥅J�)��]�b��!(K�y �RԜ�倁��$WQep��r�=0�'|�a�hz�����U���%oǀ*#�����^�z3`��rE�RZ��gۋ��:%)l��?щmqS�%%;)� F1o& ����;}�d��R[l��t���Խ>�,"T��K>@R��\,���t���r��\��W��ڱ�(�~ﶝbO��S��F̅��]8�����"&SE1lA5%K�PKyD7�������I0ob��4�b�4�@�%ŷTW¯��R3/0����mGA%�s�w~��BL������
W�J�������b��"#�HIm�2���)�h27n<�Q�Jהm�OQ=�]��)|��F9��c��1�J����;��̳���Rٵ�Af�$z�"���)�:g��Z�g�Z���g�f�O�q��$�l�!O)E`�m�u��p��Br6����� �3$����xB�v�7N�u�د��sO��!��JPC��%4��҂[~���W��s�y�¤`��%֋�x�6v`�+�Ki!����5��5:��z�Fb*1� ��
����)�k��w�JI� ��"����/l����0�6XЛ�e�`$ ���΃��1��%c��(e��p�â�	��E��浛�t��%<[kM;N�b��Y���1Só�6%�+X�
�'�%טEK��5�(���
�v��Ps�O���W�YA������m�2��&�)��z��>7(	��-��d�k@+:U�ya�5`bՉ��[|B�Pl"<�?�I�Stnvh��H�qKr����/L����츄-��\�L�U�I9 �5�'6�#+8���-n6��A����t B��1�i�x���4C���;��OTwJ�뽉�(�b@��:��Zpz�đ�r�t�y�g�\��e�O��dz
C2�� `*|�5T�2���Y�MF�����z����P�0�*]���ll_{W�R��v��y�[8�߷V-��*��-k#X���o��j�Z�$�YL��>��,U�g��hA�1��a�f-n5PO{��${���R� i	rdM��{��o�K+Ay=��y��=�@�\%�O�쿚u<���]���Z$�Ea'LM;�{��/OJk3��B�	sVV�����e�h�d�Lkhk���5=KF�i��r'+�?�Ӆ�@j@�$�e�=�t-/(T��n�������c
9uz����0��z�� ?x\�UC4�� ��k6FIAg�6W�n݂�޹Tl?gv����l��O?��d�}-d���:Ŕ�D�4�ֻC�{�si;�����=4x�X��V�V�$��/���OZ糶�F� M�uU�s����j����XU�Y�j�zN���7m^�rN`K�C���
�/l�yxV�s��Q�K��I�5E����S��`���M<V�l��.3���d���j�Lp���79��s�VJ(,pNE&[Z$�&S��Y���P���er���"�*/��%�\=�w`�V����9��On�4E�	**�b�������;� ������Ċ�� ź�:2]�,[��� �|W��[\`/5YT��9c����Y2�π?X^��9���'-.����.��,��:"TV���X�c�qfne�����4��YER\��R}�M�b�jM �1�n�l]������vqK��x�#��흠]Bπ�V��O����TH1آ l5����ʺ�Ѧ�eH�G����C����GWnֽ��W���͟�gp�ۺ�.u��*��]id�`�׊GWԊ� ���n��"yH�Ik�?%���f>�.�O�x])��g�a�1�
?����	Lے�g�WU�
K�-�Fjp�tF�Ah���> �"���H�!2��K�x��'����Y@����G�����/g�Qt�&���D�È�6�s8ɝĈ�1k�_4�|�f9E %!�3�Ú���ҏ��kh*�^��뵎�����v4��8<9��|�zH�Y���0h�ב�Y t��PR��S��TQ*�zҼ�(HPK�N�R�)
Sl�4R(C[�PLb���e˼���d�8O�dW��%��� �1���V"�����t-��-%:�h�LIiM�+M�*�Uۇ�s2�
؜8O�Q)�X����@��On��l�ՠ�u�9sN�>��dx�n�9���$��
(ƙY�ukn�����09�̼�v��~"�?X)�\v���}��>�B��������pO`�"��P�J��*�h��a#L����,/G4�x����aD9`W��h�r��(*����O�r|�_�ϼ�w{��$wt@{Jh�e�q��H?�ֽ!dz+�����{��=��
%`�� =�דmS,uC�f����?�4?���Z
�PrN��L���'����\lY���\��D[)q�Y>�2�̴T�������eF=���O ��� �*�0��^ u�26}��}��\�� �4S՚=�W/��K�&p4�ް�P[��n�i3�2[Z��/R�S_\۝�_zcB��[�Ϊ�#KD�9��-\��ˬ u|�X���ń��L���Ҿ
3S��3P�X��_Z)��j���PbR)�}�{h�.��_/;T���>^`�Fr�:OQMqY���t��/׿U�����2�N���mH��5���k�����	��@'��u��$�d	�.r�w��sd�c�f�o뢚"�M;23��.��i�A�6�{ �a��5�ʼ�:��9�iN����!En�u�p��q4��z�����P��Q�t<����ň#_�PW%MB�_������h�a�ۥ����c�a�+��J���*�G5k�����qШ�CV�A�����%�2�0�$���$,��:�?6��;��)ӯ��o �l$�0{Dس��<3��`������|�Pb�ID������C���5�����U�@�j�q��~Y.��~\�l��1
W-�V*غ�E�%�2��=��Ӣ�-��n���ޤ�Pt�(��x`�N|;.��RY���J���KxH�>���9FF���g=��7��~H���k� �7:!Zd\�W��)�����VN{�^@���u�ow��L���t�`�7��F���&�f<XLG�����J�����K	�8�~��y���K���
E�)D[Xt�/Oн�[m3Y�O6�A�
\-S=cP3�zd_����q6}��'��~�X�"���2���e<�ڴ�@�|�������Fg��6�������(lk��V�-��,������!]��&��յ�X~��X%YZ�q��?���lJ��黤��$E�z�;����<p�� �;{�J0��{�Y�l���/>u�
����2�e/>;ɝ!�Ox��h:�MTv����e�X�R�"�@'*[�!R4^=�Xj�~�X#���ۏ�g`��w(۞��Ⱦ
�^��<�`��iWd��imvV$��ry<&���#�#������[���N��J}�i|�0�����������-��S%��\��⒃��(bf���R�<��+�#�T4�=���:f6�oXٴ0I�]CB��p��D�|��qD�<�Wڻc�o
	;�v���释��+F�Z��w�U/�ƒ}|��fv�rΆ�4��tü@��	q�𡣪��p�V�ɪ*�=�[��mA����&��"���%G����kp�F}&G(R��	Z��Va?������S
�C�L�>�-��p��Pp��勳��8X˲�$`=AQ����^}&/���U�(�1[�g�2�3i���?�+�a���u/��lI�iԭx���i����5�JE�D]�����D�����2�-��e6����hF̈��^s҉ m��-�q�8����̍�_���ki�����k)��7�B��%��{(X��{g�����
6��vA�ڇ.K�l}?&2�������)�y���p;G-KB������
���y�l�a��Zʶ_]���s�vf{s�A��L>DJ��ZD�Ͼ��e����%�k_�9��+�X�dh@�G����$98��MJ�r�GD�X�~��T�S�n^�J�g�tF����%6�4L!�X�C{F=��i���85���]`�H&o�OD�mE/cq�1��Jz�B�97�����ġ�e���i\9���z��q�X[���,���jJ�;�Q6�O���+��p��uP���Z�FmG��\��"�fM �O��#�����Bgu���-,�HUM$ �L!��彟��A�9��W�s�P[���Bg��%A�/yZf��W�𮳁�*�3}��>�u��TT�%>��J�/
�����{�ϋ�N(����'-b���$*o�H�
@�5�5��/�%��V�����#���� )<�}[͢e�B���Q0��X=���3	�1�#J����M��C���<��=	���1�Hcn7Ԇ4�#����/_���"I�{-����{��,uW��Z�di2V ��`uܳ���:A@>����u���6g�����yXMb*x˶��ې�������f��](}�����Bj��g*+��bȵOG�x�1$���ҡ��"�6E�"��W�=��0���UK�!ߡc%/�y;�%�$.?4��?��W�י=V
�,���2�%�
*���x^]�	�V��cFT� �Ա�uu�������]��J����%�SU��w�	5q�"s�����^F��h�� �hɵ��=�ר�X�ט���O�<B���j���@�{��c�2�� ���(s-��mU$�	U����\� C���l'W_	��Ќ?��2��~����V4z�eY�(��ɮ}�$Ú+~V3jqB���:��M�TW�Z�>��m�\���0H��'�k�vk�n�.:���1$u�� ���qv��!7Q�~�f���4mo�!_�\�͜�ӡ7=t�J4���L+P�W�E=;xtم�+vCer0�Ǎr�7nN���h=��]Rl�:��<-.(�t	:��%��dB(��t�m'�Ap��q�p���q���G�6.�[+mṔ�T'�"���7�%��*���$o~2ts�&�����&0�J�65 �Ů-�y��{h��u�{�Ō�ź���$?a(,��ri��0]*�s�B2"I6�,�+X:,Q�
n�N�e�8%_�����Vq!��.&���n�W)����<3 �����>Z��>A/���-���;�P� d �.���m��n��2���T�]^W9C��E0�{j��<K�+dՊ����S	pi�;]h}� 鬗[~����no(�T��W�Z<4����ͨՉ�������ff���v׍N�kU��Q�H�w�B/�&8:�O�� Dx�{Ѣ·M�����	+�o�ek� a#��?�������L/�t�� �����a>g[m�}o�=}���:�[�x�$�!�aw.X$|mK��mm��P@��l�1}ϴ:�j���4 ����<��8O���ϩ� �]�k����`X��i��"I�q��|�b�C_D���<.��{�AM�n�2�,T����^r|T�&��v+�ˤ	d�ׁ��	$EE��]6�>�� �N�zt}�A��?j��5_i�W�w}���3���u�vc������o�k�_��>�H�\�±|*���G���^����|!��"j�}x��A�d��+dp�*��j��o]B���x���'QE_J2{~p~Z��~��D��Q}&��{�0FDv�唫�|�M(7B�$
z_COnkX�Z����F9^��V�ğI�]CV����U��2��9���Y�a��v��H���zKTb��� ���-w_/6Y��#.u+[ȋ��,@�k�Gʀ�9q5��y{ׂR,8�۷����[�EwiUf����	̥�DH�M!#��{��Vd[��=:!��w���yQ&��#�+[s@���b)�-z��)ܥ\1`$_q���&<��bC���5����#��$9ћ��x�(yP}�BʹR����{<�Ҳ��{G�E_�g�f�������	b�Mw�5��MW|S�|�އ%�,@�ke�+}F��.�ZEƯ��$v}�Sj�py"�2��ʅo;p�Ɯ�m[��*���Y�Ny���-�5�����p�@a�������i�ħ��r�X�%#��t�C��8)u�fu�g[#̸��ۺ�W"ٗpP!����
%X���y�}Rh)DP�ޙ��� �$~_�^��+����7|�/w���Q��6*��*=黛�(��Í��ك�Xvҭ�ՙ�%��}�X�MpBcIl��-��Bb��k{s��
"X��w0�c�W��{E`��hL��Bu�-�h`�g��0�έn�3t�D��+�{�]�,m�BȚL�vH��6i�R�CI�th���qIE(�D�ƒ�"��݆�t 8��r��[�X=��1���H�Dh��Pd�꫙%Ṻ�j��*@��0�߂��o�j8�K�i�=����Ι��9φ�_����j&4�K ݋��|~�Hڷ`��]��n�V���k���<���'P�iC��)`O�#Dxb��y���\VE'ۿ�"3�]uE!�{C̵gj�%Мv��!X��5%�9g�#���W
�v5�ϫo��A4f޴�{8������ńq�7��w��G�p�
��r���i"-�]Q��`��ּ�,⬇ю�U@ɟC$�[�@r��\�,?Q�q,�+�����^���~s�#�f��##>������J����qS�|⨥y�} bn4&Fg#!��T��pþE���q_�z���H���kU�XtPo��su��<%/8��'㖘k��rmiD=�>����%��Z
9��Z�|=cҠ��M	f���B�_�$3��������wD���G^��5�<���x�ζJ�U�ӵ�yN{eP����S\�q���T~�&��ΎN��k宿���̱�p���Cv����͖�=�R��!� h�GO�߈i���a�`��
��U�y��MP\��Y��E�#�~ڔ��n�8c�И՘�S`�S�/>?�0e��q���˼kw-��!J��2�S=���o|~
:� �O��2�Y������:w�T�)f_u����s������Ʈ�I��o:�<fZ�1f�d�7QBG�^�$�T��MDa�y�z�q����ާAK�[rB/��4-���w�+��=��30	|@o�]�����~+�A��+ҡ��\Р��3���;W�(#��D��~@. }������<;L߸�������m�����������"�N?	x�j�DC��Η�~t���Ǯ�9�گ��c��i/!���Jl�^{#�q���*1T�r 1��=�=Xަ6\�`AV��$(��h:�뎗� ��P�Y�+���폜��~�Yȧ�	�Y��!ʕ�F¨SW��n�F���,�}��~) 3@��gx,3�U��;�l
z�'�{���m!U�m��s��0�2��-��'/�]�M ��>A�s8u��yHP%�/I/8@���Ѕ�y5���&y�����w���6�o�Ѻ��\�/�
�!��V��*2��D��OQ"��,!�aIԑG�v�x� ��nJ��HV��}��N��CW���L�8" T�%�Ĳ��m+�f�p֜vW?��qV�bLV �33��|��C�
1�9�5t���D׸��/DP`mm+�O��
{��B�Nk&3G��|���5O��r`�I>�`��u
��G�� ����������@:�����BP�@#��q�I��B�A��ȶ6��*��:I#Ԧ�s�2��T�e5�u��1C{UM�։%�܈E�mI��l��V��4�|xV��J� _�+�0p����#�W�8=�d�i{x�y�]��V�F���FiyY�G�`3�Ca��}'���}�"�G�Gq��ae+��	���F{���(�m���'���Xn�8��F4�]>Y/��X�6��:�3!��p]�H�~���晵*�kf8�.��C��p|f��>�x$c7� �?�jc��	N���uL�#ӈ�h��W��;А<��7K|@	�E�5���`~��*��|�~� '_6�ݕ�9:"�Ome��-���d!CU��V=kS}%�eN&P�jT�f4�q�Z�&Tl�F�0n���[�6�p��7<}3�2s����Z�uŗ�̽eR�v��E�m���J�<�7�B+��ī^���S��H�%����f8�>G����Pg{�YDb�JJ�	*�+r�#�*ψ��xb���U^uH�d10꜓+5�	�u��d��-z����j����j9p�e$�x+�q%�1I�x�I 뇼����QT�q�9ڷ�O��Z`k��v0*>�Z�a�R�L�˲���q�a��+JE�ءC���@�9�}Y�U��Oy���9[&�i�#��8Ǯ.���&�	�&��� L�j{;�V��`;y��TK��d����}N���øU/�������T_\�X��ڰD��c�-4�b���#����
K��')���J�zt.p�r�*[���GRxzcq9R]GH�B�?�����a�!NeHKH����?S6���G0 ��pu;(���,�&T�9UQ�2�-Sct��'pH��b��r5A�?�ED���i��P��}(��X��zX��8�5b���W����<pN5F(<y����}�%چUn\��
�
�$�V��?���TW�Reu�J?��kp־�F[�t1�G�#�	l�I��r&��|�	�#7Uni��ʚ��kpR��@����n��P�n4�l"��_@����%y���+��Բ#0X;�������	E˦����9�V�_\��5�CM�:��w����]5\�=x�<g.�_�Vϧ(::Y�hVV�Eq�k���k�����ŵ�A�O�xs1>!Klh|�|�opJ��}Y��Y���3��K׭�c;v%	
�k�P��! ��[���j);��TpS�c��.]wI|RA����3�
�;�����r2UG���3o�*}�L�)lβ1��<s��@i��Hٝ|�6����(F��W���1�ԍ��#���&�Ht����H����S�����kYJ�]!�C
=a)f�AgD���= H�M`�?�B�� B@=šoH��;킺i���ǛoL��0�� ��BvoZ��]��-�{��>�%,��;�¡&7z�F�l��9�ck)���_�jucۙP��P��5a�#��y��b�DxcU���t�o
	��~�bsE(�OGu�0�+�Q�.Z����T���sT��>���6��EL$��5�ܷ���W��73q������&1ߥ�o�� ���1�-�i��ݍ����"R���t��_[1��=�%A��Q�  I��r��_*hmKx7Bl��;�`$�B��-���1`���P�ʣ'�4�|aB��']��UY����zL��.0��t�O��M�T+�
���_C���Q@7�;��f�Ҁ%�n�Y�u��� ��i�̩��JL��"0��IS�����t�{7o��;4'�H�g�&�>��$�j2�I�]0�uK�~U��c����z��zs����	�"S���"���E	I��3A��I{�h�X�Q7¸�IQN�\����D9減Xwm��prJl�]!yO��:��vf�?�vT��P�JC8�!�9�Ph#�1��T-�%Σ~��a���$��;�4��w�-�:�1��u��r��)n-��M:�aq�rM��
q�m	a��N�!>
��Yt9}�R�!:�X�ϹqV	f����c,�(��a�&�I�2�(��ގ�5lSI���Ĝ�l� �K����'G�s�ɢ������X@�7HO
b�sW�g��g��sP��~}?'��yN2�4�X�����z鸂u$N|q
��$@��z�nJ'��sR�sǙ$���;�N�5Lڔ�G.&�T��1�%�E�Y"�Z4=娫���]��T-��V:��E�ie8E^��w�.�a�/׹?�A�cJ�3�Ϫ�8��WX�2o���N��{!��aݻY`SC�Ѯ	t��SKI֯?jђ�1��m]�;\9�+���%��@�����e��r�W�6�b�%H�t���<��g�`9������/���v.^�{�dJ�Q���gs��'(�a��>�x\�������:�a�Y����i���=�7G��&�NB��`F��*/��:�b��\b��L;���qav���7�k��rxʵ��@����+���,�[�8k�ŉJ:'I$&Y4��a���SD]���_�xy�뵷߽��)bIA���䙓���aqH*1���w��- յ<��`��g��V֝.P
��̓��D��C�h$�s������J:��=7g,J�	+]�L���o�g�zG�?�F��k������~mLX�k�l�D���T��A�lוa�Z'x���;'���<��"|>�b�$���q|�^�@�0%��"C��G�+���}�!���c-~d�9���t�w?�q�M[DB�fhb8����c�����}H]��y��}��|�ԡ0Hyv�w���@ގ�&f��O��K�@K���("�ņ@��QBe�Rdiߎ|曌�MiP�2��n�\�I�.7V~�����BWR�˅��i��.A�u��~�E���u|E
��+T�Z�������~�٩3U����sw�����`��*΂�g�f@��	e{?b��uUKC8%Gc�4�
'�q>�D�q���/�w�X���g�*���pU�.�?Cń�XFV�i]�P���G�B�
i��e:/�nt���K�n��5���_|%�e����x
��?4���I��x��|�sD�.�yɘ����>�r�|��WV�<�������!�Ɣ�7��%zR\�j�)�w��z���^-�E@Ī���^��g�3�� �ݧ)�3����L�h�ȇ�'*�lyu$6D��l���<vQHւ(�֢�\��H��%�����a��B�F�t�;�r/D�җy�� ��4q��Lv�32��}��~��2�g<e�,��*�Ѝ߁Ż���Yџ�(�U�l���͸���8�G�%�";Wb�n�
�Zy̝8��Ά�M�.��̧P� 爡����`p��`�cfu�SO�h�{�c=��cO���O�3�.��:��9��i=�ʷ*�ו��7���}�cN\�k�=�ozQ/k�7��Q��=����T�sܹ���7�Q�t�l�I�m�-�S��ѯb2��~R�Ξ������򲱆*:,�,AE�^?�]8C�otH�m��vƽT�5��Q��ㆨz�X�/(r{�#���>�*.�#�Ԁի��Dl�J�)�=˖��zŧėI�0lGq�!����^�'��X���q���N�S~Ɏ��;!+[=��ɤn��ڙ̈�`Q��W����{ܭU"��΢��t�)t��oQ�ә묊�=��T�������F�d��X(�Ax�ߠ��?�������Z�i�J�C`��
U�,���7�R���� i�zS�7�����F�X;���
 �j�+e�=��������bF7���XR�����(��4ւ������TJb�hU.�i�Ic7j}V�S����B����Ș�2\���{Wq@���Lq9�9*��}k�`�kqc]��(!lݽ��=�������. ���h]&�[��1Ʈ�T�6z��"Pt��M�ۀ����K�y9_���"�s�8p�h�[��gL�G��8'�)1QbdbԄz��z��_��'k����?�L"v��lT�֢����/o��;
*!������z(���BE�?� �]b��ϫ��WHnR�=���&�_�s�SͶ�����0��q�+�;ry$f���
k6~^w��t�w�h��G����~��aF0��l�2޻�Ø 潋��3�O�C����DCc����M��O�k�P�ï"xB�ՖC�R$���tv�|ގg����PW�Õh��u%�h"g`��>�i��9Of�x�=j�kC���֘���A��La��k���QgM)O�998�~��M�pJ�\X�o�Q���]�˫s^�wE������"�ێ��̓-��&��.��S*b�B ��f��!JX߲�$R��g�cUQ
�˰[�B�:���d+S��H�9I�ǚ�;H��i��Ԋ�蒬 <��E�����A������c�gCy��p���&�y��ӡ�����i�����>'3$#�1�q���Z�"qk<m� �>9��/���f��-re�$CL��P��\t9 �%/���������g����8`��*��x���6�#Bn������.Έ��ru�qG�6RS��~���+�S#�D�!�ߧMзj�v����3�N���b�k��+
8������޷��.Qk��L4}3~/'�2�u$�Ddc���%-�ѝ/�j�`���o{{f��\࿁���ٴkBV�
q.����]?d[�X��@x�
e�[��sg�� Y�_������u�G�4,`qv^>{m�~G�rHb��e3������3��U톅 Rp����Ļc������R�G����S}3$Ӊ��cX��oU���l�s�[��9L��Ӄ2c�<t�Ƨ��f���׊� ����J�����a+~�:��Zz%b�XY�p1'����%G�ģ�15nY2�;�f�������_�8+�7�\LVT�o�E�F	�I��]�����N�_���
֊�N��e����mQ�M&ń�$��QV3Y���_�	�`��Q���{<@2��k�j�圼�e����kO��zxsy��ɉDI+����0�̡.-:�;�w��[�#Oݏ����:�<�h�.������K��P��|+�o�
��	ƆJ*N��X4r��ݗ��xɑ�}��D��M�;uf�5z��pD7Oi:��e��ư k<���'(XIka?h�q"Շ��u�{{���&���j�Q����<E�c���9ڗ9��9������2O���!�zR l`�}^��948<ƕ�W@�?��GO��d�X�`{�%i\%$�-R�T��K��b�5�ʞ�r�7l��y�v��\5iԛ���m����`���ŭ�k}����w�I�+�~S�B���P��Dڦ£�BV}u�LX��^1��e*��B��Hz	��=��ء��:���d�7`�_�����h]�
�� ��'��� �B�7=1^&�;�QO�	�b޿jO�/�%�]��ə�̅���/�>�,h���,���g����>�~֟� �ԶAťg����W���_i��h�r0^�Q�O,c��/&�尕��*�IL��)��F�ѩ��{��{���{_�܏S:�*�h5��g�ל�.���A�|��	���!v��7V��gx@r+���;��bS��%�SQ���[�mBU{�28��~ r�	�������?�qQ$���+��~�@o�j������:ڣ��)8�Pv~ ��փJ>]*
��� Y����5�E_�d�A|tf�ف:�VY�ׁK� �)���$���RY
o͚�Q���pt��Eד�,�Յ��s"�]zy�ZI�dE	܇(���Ʋaԝ��vE�N�5"�>�)���g�n��д*Alx�5G�\���Mviu��۝�����|E�q�'BeJ?ta]:�}j�������b�a�0*;���?}+cX���>��)��"��*_�z����H�"[�7*jV�~��ZUL*;��H�w�
�{&7Ad
T��G
���Y(�,�0�����3�u�TL������U�ĩz��/�b�s19b�u�R���7�ƀ|2�|��	����ڈ2QudR����3]�{�>;���V C�oAL�#�������r+� (h�t��'�.��^�{&-I?sy���	���ݡ30$Pgsΰ�����dƱ�Xq+[�5��h�����\<@��q]A�kN��%J�4�-���9<eR�t��O�t�̓�}��!�r�m�.&g�:$�+�IK&�o�3_��#����v�&���s�х����xT���
x*��0[��g��.6��./U|�?6�4D���dc�cD�I6�D㟭&=$/���k8P���Uw�4����c�s��2�.���y��6����̃>qĺ��s�q,� .*~��[��U��x��}�L��=�u���O3����r���%�z�"�w=���L��[v���˩��gh�]�F�8������4��/�0ә��]L�j�fn�J����dB���� 5�=@���j�(�	o�k����g�t����s��p~vd,N��W�7��z�:��[�`^��g
~�8��Nd�ヴH��T�����><��G���J�D��dI�7�n��YjL>V������o���h �iS����>��l�dX�k�3G��J࿂�T�(n��C�v�[!IJ�I�ж�nP��V� G�b�jv)���ԗU�r��L��Q�%QWk����
�����so�e���h���cA��
��I*�mD&���ן�f��ʭ��'�q6�pF��z'd� ��@p�I���#no>���r��c�hM��Ib]
d-���v{y݁}uF���t�--R�<��Ń�L�:'�8�h�d8�.V�]?�8F_e������06�6V�3�MSLw�i���I�ǐ%h��	İ1��e�5�b�JQ�d6�)xYZq�9�Z���i�#ܙ���d|Q?������৙V��z���Ktkh���"]��Ap�R7�8����?<�̛�����n���E�53���HY> a����JF>N�Kp9���49n��,��W��T�*�j���������ZT�'�M��܁Q+��,e�z�������M��������T:u����?�Oć#>�蜰��U�SB���_�LX?D�p_O��n���lF��� 8�y��7J���S7��U�+�,e�5Pd�"Ze]�=Ɍ�B��A\��7e���<�;���W!)���jm��R��۬#�}�7�9f//�
�K�S��Ծz]�G�%vM(��FKb��;��~�^�RYp�}�J�E��U�m�)W{��oXo"u'� l�0�͍Jo��$��@K��a�:����q��ں��������^��F2�ˋ
���2O�@R��g�?x-eY`*��A�}<J�p����<��"Ȳw��F�j�m��>�c���w�I�Eѳ���ސ��s�2�P�_/bv�qB�e�P��	
�B�o{��WG�� 1�=��G���F4m���\r��lZ���c��'/en5_]�� ���mW74eE�\pn&;��ļ�T~�v�/�A+`�SIⅰ����Ѽ��!����ַ�k5 `�A�P�Lھ�2����y�g�ۢ�	ēkE`������驟 M(�*�)�zw]��l:eV�B6�h�U��Z�w%��n���s��s�s{�z���;��d�s�%?�n�� �m�>���/_�Ozi��ތ*ݮճ(��CON2j� ��7�v=�c�	ĩ�����*�Q��]2*�A��x���v��-�o=<.6�Hݰ+�jx9L�����T�K��ރ�
B��V�������@���|pF��c���C��(�6���)\[v�r�����^EE5ҺHS�0��TW�WSd���{�ː���.Cyҗ��d;%������{��7t��9{�V�����d��y�B��C��n��K9g�Eo؁����#l�MKS����Rl>��R9����a�_��ɑ1)�2�qO�r9j���WI������E ea���칤��޺9%��#��&>��71��l�Rk}~�t�������I:�8�f	%���̏5 |�B�8�Mʠ~{ �e�,���y=
Af�����ذ�gNN)��0��. t��F�gM��QүÖ7%��M�+z��^�Jh����i���7G�t���Swz��x���#�~d#w�Bu����tb��l~��*?�goXPx�ʞP��0t��C��Z�#�I.��䝗� ��hZ���-�0nM�g�q�.m�E��&�'1�+��-=��F���b�.5<����w�}u��.���|4�|	�p�1��؋����|D���\&���܋�+z���׎O�{l���<3	0��K�j�j�W��oI[��UXPG��ڳj>C�p��}��KalضLyj}�W�U�9%-#9����^<j�7j��g�={|��B��u���+E�Ϝ)��8�����9�Oqp�r��CV��}%��x�MV�/"���	�C���%#D3��*߄Ff����\ED��;݁�yXqR7;T_�������#�mኊ��<vs[��;��*�_�P�Y0��6=�r\�c��.��p�祩q��/�r�a�`�U{p<��JK�^��k�yHbxyLK8�B8�`�b|�2@(����ѩ�tAdX(����b6��Kpi��I�8���������e��ol�)q��,���k�������R��K�����Ο���ȡ#]XCP�����e�%�Z�,Is��E�^e��nr*��OJ"���ã/O�d�24��Jcշ�o���L�J�dH˔8|����w�ᐗ����d�۞\�X30_:�	~����~Ag�i�ψ7��66MƄ��H���Tశ��7F����d*����g�g�*��ݻ���ʷP�;=B>��@�I��j��$ڔ4/��'�p��2��W�٬+5m<���j����xa���@"�9If@ 8�T=��5>�Ѯ�y�` uL���k6#~�e�5Jt������KS�ԍ{ /)�X�@_�U,�*xH�엿m�1����gd����Â��vj�~�7Scx��\�:db� ��s��=����� M����D�na�悋����}��q��l�����6�j�� �n�<t)�{�0����G�w�OF�r&^��J�"or����}���~zi9t�N��\��H�5�h�籯�qQl9��aۅ�K�!<��|bO�����f��FQ��!����؄:q�;�s��I�A@xv?]?�*�ZH,ڮ�^4�TCv���_{�<;~s�DӝܥH��$:����բ�%��>����d0��2=�p��{٪��P�G�^�/�3�twO��b7*�J���f)̘ľ��j����Ir�#�Ϡ���_Õ�O]���6T|�\8�RM���ʌ4v|��+���o�+G�i�ڎ��|��x50�����l���A��wY{��s����~��W�L�C��rH�U��D�$T�--wB�T��[�Ē-~Ya��
P9iXN�R��6�Go�\]e���Z���q���N�@��)����H�_2�`&̳R�W�'u
��ٱ�� W�����%wX
�c�0� ��k�	p
L�q�ƃ�C�fDf��86!���
+$6��o�ޅ`[�W����!O���gn����_��5!B4�#�U�$��k~�e';�p��w7E�Ep�D�e�BXA���bM7�܄�e��B��?�֗@v�||7�$���Ɉ75_��k��h�	4��[Tږ��;�FTJ����=ɖC�2�%����	�oWz5�3��?5~?�l�Ai*ُBn��N�V�S00C�8:֡�h�,@	��&����c�(3�>Y��%D�Ч�=wի6g���/�B6�����Z��5��eS�M���Z?���9�K}�`�&�\? '�"�g��b�4��Ɖ��Ϳ��2���Z�f=~
��fK�C_UIΘ�� ��T�J%yci����3}��Hn��@�Ĩ�lwS\��/a7��ѵr�f�>]�QS�~/��s5�=�}�(��4�Џ���m���+r_~;f���|�$VK���4m)1�����A��N(%䒍}����jK�6���r�'���-��Zo�J Y&Y8;�fv���ջ�Ӗ��-����L�2��^�Bī-i9�w�]"��B]���.��>��m#�WGE�U p��E�%�:�]B�(�?�O��&;��r7I��M�z�),�-�dSg��`A�h��-��?x�N̓8�ט⺻��+��޻<~���tPQ��^,��vMp� ��㖜<�Y#��so�u0n�*�>^�O�I�f��<�����=X�{uѥ�h-֖T�#�����725`���
1�w�ґJ!3}��_��o�2���_���A����D��'����l�hn�3���·�U��R��C<��v�P6�u2~ �ۃŗ�z�}����E��5J��U��!�����D�V�~GK�R�M����Ϋ�}���Q���f���א�X�T���>d�1TsܬW����3�NX�9�ei��"�ӭC���.2���Q6}����Ƹ��,�OX��4�#娍����:�d�^��	Uɴ�-�\�n,5-�<�QHZ��s"�F�)�3*>�@}Ѐ:P�"y%q�t��E��k�U�m�ຄ���qфd_���w��>�k�3����ުe�/��n/#�>nW��~g��|�=W8�P����y��'��Y�͊�R�B:�7Ӹu��.ۅ\������R���Y!ͫ�.oO�=�%κ>VbspR1t{��M�"*��O�/�㥥���~�ۢ�io��Ƞ>�w��A]������7Ȁw�%�2�Z1���:��n��t[�o�~)����m!A�]ˎ�q{ZB'(�$��ث\�'����?�����PV`���9��2ώ�(�����yB�Vv~���h0��R�q�h��>�c,��'�����'��<Қ�|�r�a�:6U������o+=>��_�$(�Ul|�\��J�Pi�ŦtI�d9���sT��0e G�?��k�[ڏ�Y��)6�d!��[�C�(H�j�=���v%<����nZ�0���	�G1b��g�E���:�> ;Y�bp�B�l����Y� ��/F��)�/�|ҳ�<Ck��u��G��Q��i�G4��`_����<�^�P�]�*�AA�ߴ]Y���+��h�"��ndd[oRrĚ�yT�kM@���-	"�ԩQ�$�ޘ/���`Sl�ccY���i����~�"�h���s��k��E��A͎�y��.s���w5dN3�U��"抆yf�Ƃ�cg:y�5j���Q�0���S����Q`����Q�Q ���^�{@Ƌ}[�&aeWdib&ҥ �$}p#��Ȝ@�Y�Q�X�_S7N'XZGȈ�3��N~9�)}Ĭ�TJ�}8��TQY���20P̄n�}g��/ ��Zs��=��������yܨw_	��X)Мv��DԶ6��R
��IL��6|�UG��pr[��Ky�$n4����9�6��cv��%\;�Ŏ#�:^��]�H��enq�(c�LyK��d��D�۰xԏq���rS�Q�%�O�kz�>�[��g�R�/���<�0�k��(��c������9�����)��<��>�������jܛ��l/���j�6���qm-CK��>H�d��T?�/�/f�,ϝJ�	O' ���DΝ@�8&�cZ')�c��	�^���������l�"��{�CG�l$�K)(�>\!�m��=�N���B�Ɩ;�����[Z=� ��n�&禕>������s��V�@�r��LYJC�w��>���5M^���}�3r�Oǁ4� ��h�A]Ob��r���p0��Ͻ�ĸځ��9T]f,A�J�

F�buj�D�������ޖ˗�>N1�H;Ѣܞ�Y�� C���*tF���d�֯��7�xz�f����vP�����S�S_ˌ�Ms:�^5���l�iT�?zF�)�/$U ��CNI����:��mW�L�q����<�&�^Cբ�G$�1>*}�"
��RV��	��k6ۉ&Nl���&ei�C� ����U�	~*��� ����%�m�9����^�G7UjO��Wa�q��!������M������Q��@�)�.A_$�R5�d.HH-��D!�$�����-&�r)OT��l
<��㸺]��:��ln�֧-!AY���8t���eP��̊�ݨ��ƾ!�
��'����� ��#��+L�k)�#�a�ZBB�q`�*��	*o�x�=���i�J�g:��[�6�8vT��ak̭��.����p�j�Exc�V�`�����ϡ����p���������Q�Q�UP-�E�X8��	곉�g\���o�($��8z��XL��u	����皑#2�����e}j�Q��pWݶ�fk���=\:�7>�^����:Jï��e���*�i4!�������,hpZ� mڢ7`l���6�O��j`ewJ|d�	f�>��c�
fOe�%i�N'�Q̡���u�h.�r�����=?�2��&J.p-|�&+	��U�]�5���@@�%����,<X�N��X�������� ��0x��Ǭ�t��c�{�l+^����
��/+�>E>���� p9+�,�z������و��Mс����(
��ʛ젖�1���ʨ�ڥ�v�O�oӻ���/ˬ�N��^�l��@�=M��6��~s6`�#F��w-h���6j�d�ćw�0_>���"D*�U��#\�Xr�B
mO�����i3��ׄ4�	pJ$R�qvcR�NK�Q���U���I�ᷰ�\{�5j4�����Gt��IeQن#\�Rh1Uo������&�铮����`��	)
��⥓�_?�c]�F��hZڶ�r!��v�?���a��T�i���oN=sh4���h�}����nXݐCn���,�bm�7tD���D�v%�Y#��1��!$��=�0	�;�c]{�=.A 7/���=��MIJp,��l�k��J��n�_`
~�yH:��:<�����t=L�0+fZ���w��+�G~�Ag</t�T�{����O��^�p�{k�e�6mq��t�u��<���TA�4��T
˜���?�Y�����34GϦSN���&I0�����I��h�����8M\A:�"����A�E,�_op�m{�+V�š��F�a���*��$Xz|��T��ԝV~���ּ���Yݴ��������MO�sG�􂸧x�?M�0ԣ�h@�u��jBs���:�aE �`��Yl�b�z��g�c���J�t.����+�*-,�Z�O�G�q�#5�]�O�+P���c����"D���*�jČBHTF��lע��-���)�����		B�}a-�g�yG������F��M�"?k<�E��p�ɕF:�T����b?�V��p+�N���Q�Tۅ3)��C����b|��ˉT�s��E)�`ר
,�L�����l�bx9*�#��.��C^E�tA�R���w���O�3S�=�P�ݴ4��.ܵ��p��RN�N���zB�������/W�B�<خx��wA2b�RE\� t�������~��V�;L�f=�l'~�)���y�K����#��6�G�`S��z1j�C�<��@-H��_�h���!��y��W�=�{���5q��7d���׸<?G!�
�7STKj`���7H���X�׃5����9�������z|߅�=X�g�K��,�I�Zw���{���F6ƣsG޺�U�����؁5kj7�3lY#���dC�c�J�LbO�|�/��ӛ��̼J������'�Z3�������+�]��i���l��y!"=�6����K�{���-A^���YT��J�#�2�Ֆ�9SƤ�� � @���<-�����������T;�Xǅ�)�Z7��7Ɓ�cD�Ab%CU��2�=���WdIT[k*1{�Z}��Z��X�	��B�<�m�G4{ta��jEM]�H�Eq*R���6p~C��~B��Nf��X�Q���I}�\������hx�U�/mx[yݢш���&�N\/��\��R%���+*�v�3�ʀE+��9���v����lf�q��`1W��l���%!��l{i^�9���A��]�I�g�cX����R�P��w$�Ip�l�,>�[[�h��Y"z3�*I��~�(q��\��$���iT��q�S-,�r ���#z!s��֌�F�rK`��,	K�l%Ϛ���?�?�d}��~�:UѾk��y�����*��Z̟}����d Eh���foŴ?�࠹fm�h^a��Q�]e)����+� �I��Xn_�U�hk�IG?!����
��F����se��%ϷA\+��my|�aO*h�P���M�#�b�OnC�!���7���S��["���N|��lu�D�J�k��/�\�C���nǑ�8!�:�m�Ϻ ҹ@�	w�������A��.�이�%W{�������ڭ��4��>qe��V����^�Qt����^`�p�ܤHh�i^\jk�"v�.��^'Ii$i+{.N�8����	�w��Kp�L�@�S�e���#�H�a!h���g8��d�`�Ǖ'��$t�������`�-oj#��^#V�7y)�X�z�ϻ��ڑK3H�t�i��']�4�_ؤ�"��.>��4b��cY�)AE����/�)ޓ\�-�D��f������}��Ў�޽�@�"��X�x�cܷ�O �;{>4���m�qTT�&Ձ�<s�w��!�$�9�sF(�Jp~�JrdT����&�݋���9�ޤ�)�38�%��M��&�f	�Zї�'F�˒��sXi[�q���Qz��a`!��J�	��%
¶SO�@��|S['[����W>RP� ��eGu����
O�n�q9[�T�,_w���݋=�����u�~u��� -��xQ��w�/};�Z�7kz���`�)x���Q���~k6rk���m�C/	� v�i7Έ�4_��9����8�^�H�&�n�ra&�(z���.��|���E��"��)A�&��e~
33\H��?p�ңr_A�砂����)<s�Eoǀ��3^�{�	93}��Sйc�!7�Ҁ!��Q��DER�D��hL���v�?�
G�-�Fm톔�g�]�~]S#l�oζ�j���2T�AC���$j~�����t�� i�*	\�~V�j�%��qIJlGt��$�h��ޮ��g�k�KS�٪Mٯ�wM1(�+��j8#��^�6R5�%6Hg��OsL��%� ��L�(!�\$�ԝz�T���-���4��*qt5Ԁ?a�L���F4��|'�8ό�0�s�<��.���E�՚�������)�Z(}�(�xOk�V"]�ϞQ�_�Ou�^D��"R���GZ���v��k3�cX����M����(K3o������c8ڻ1H1*��=D����1�]�66���,�)�јI��0בMR�R�ꔔ�\Kq�����?�9�~��V�sƷ~r	�s���yJ��$�ޢ�U�k*u�F�ԗ����:)���+'v�;E:5��Y��5�3ㆶ�|n<��v�?���?�q9�Ī�P��&��dǫ��<|5V�Ń �(�,�	ӪPn�*�h�Uv�&#R9R~��,9)2���:[Ѣؕ[��7�N
��җ�~�w#��j�����@Rƈ"s���|�}d�B�4���G`zT#��CR.^S	#B��i�h�T�_[�/#�� �/�/�
�4m�.��@ vM�YݸQ�ъn؀@�D���9<'}6te�H��Oc�~�A2��pص�E���PS��@�B����4��$g˙�����l�h��F~;��~6v-�7�K�*�?4?˩$_�
7������P�7BGn0I&y�V��O��D��D�Gf�F�����jP�2��x��⫲����>��0�,�UH�iJ�L�Ҳ-=2��E��l#���T5���>�;���>�)Sa��9T����
`%WQ��(�!!�����)��!�?����ԉ
��}/�8��1��U4u�y@v��Y��E=�y�m��Q�i���|48.��˄t��Ϳ!]T:S��M������ݏ�g-��K�#7��F�C8N�S�V_[,h1�&��s��ҵ�U�ܜİY����T����s���x�rSJF��mW������`�4~T�N�j3�+�y�S���r�˺3�Rn��⟜g81W�e`�A�<%��؈�]o��EYY6�BA'ԃb��I�ݪ�x�¤<$e�f�V���m��:+�©3[�L�áA�Wm.��㲗S��g[YV�-�^�Yf�]}N..�|�EJ��IXܥ�h��$���%�&U}0Ƽ��d��k��DE!n�2��dU<�v �H��5Qn#����{�E�=�K���o����(�����u.Y��� �'�+��=����s6M]���(������n��Tk��:p�b�W��!�����R�H���FWe���v龣l=%kOW�!����k���~�Tv��0Ջk	�[SW�$�%�_i!%�d��Fܴ�PV��%;��px���
�/�2Y���{�p$�TR�f̘4�ε�0��
� �����<�$A���������^aU���h�c�_��#\ާ��]�[W���Ϙ���A�?������d��%_̬�����	�tm9��{1Py��:�7�c�\�Y�Xd��u��?��h���Y_�@$L�����Z�?����@q.��h~'�����|?op/����鎗�"ϳ�p��4���-bsUDo�����!���#w�;"�p���	�B��,��4cX�Г���D����(�1B�kj�	�{�2��t�K�zv��H�҄rt6�!ٱϑ�m�O��V�p�n,�����i�S��(+�NYx��+�������ՙ��b�9�?nK���vC< z�ǘ�M�?߰-�� |����;�X{/HE������1�����C�!2G*���h�����Q��Gw��1|6|�] 1�/��Echf�#@�Xq)Y�yj�fY/�2OC�t�1Ԏ�h����u޵��ړ*�W����o�L�R�)1�p1�Gu]�fF+l{Z1�Mhe�nlH5H�:ہ�G�����q��z��oT����H`�w�\��u���W�+`�5��� 9QI����������7������/g�^QQj��k����]@�
���E�AJ���ox,eT�b�[�9̜2�t�j�7`�>�zqQi��g��#(s;y]���]O��YD�4�ꁁv��*.�i
�g�ii�H�6"��ϛ�%�,(�h6�5���3!=I`��G���C/�B���^�0���M�ܶnH+ҥ���r�9�FJ��^�ʕ�������\_��'v�|��uuN�C��Տ�깁���EO�NpN�����]Q�J m)�O$1�(���f[�jsM!��v�!(g��E腌�;u���]B�
���Jm�oz�s��/V�D�����5@I��m��4}ķ5U����Vz���p���/�pH�d��a���D�����D=�X�|眃}Y|��w�xZ��X��6��q�&c^��Ymk˘x�/�Y;?Q�P���r�k%���6d"��Q����2��e����;�� @���v�tЄ
��U�����RB��r �T�Y<�9/�g��0�����c���`�o���+~im���R~s�1�d�C��?ǫY"���r�E��߰��q/�Qz��l��5C����k�ꯊ�H���l�"�R.N��"����:��jؖ$��qj��v9��x�@�I�c� ��S0p�`����2tl?�Щ:1�!�ZI��A:G�S��T�aTЈ[Ԯ�����Aۡ�]6!v��R�w��4X6(��'�f5܏��"�	�W��Օ	�����
~�T�M�+ƚ�_,Ղ�~��l|ϥ�&�ǒ-��^$�ޠη���sh������"��X��w�)�t��w�.�����HV�|�K3�j�i�|n�I�����hWٕVɘ���nt���'YY�����p��ʺ�����peE�³0��:����������g�Z�{�����|3����iN��7,�g�N�l˅8M,\k�	==�紞G� o��	?L�(=���Z�ϫ5H߮��+����f^�=��"�+�X@<aLTRJ�cw�N�D��p��~��K��V6��,���kpf��:]��=�5փ~�\;b��XJ>�"�*�̱���	
t�l� ^� �����38�?FloҵN�!�<��%5��sV�C�H%��%��%�ݮ!�b&4��Z��~x5�Y��[=E� �lT��Ud4�g5@|�ߒ����f�%Π�QG�tF���~)$�n�v�S<�)Гg��>�(� ׏�<)�g�b���AL9��o!��-����~6��	�-�)0��T����,��:�=5�Oh�o�]���䧪��lT,�xb	��n�ju*�m�G��h��
�h"������ۖZ$#i!�$I���%!�a��K�U{̈́No"s+��9V3s��W��k=y�|�<|>��N�v�s�*~���C�sh*>%+M�4�[�����vi[�>��D� �'KمÐ5�A4��l*�t�Hm트�:�Y�0�9+�H X����v�B�@жX�4d	�D�ю��d�+�3"^�/�4@�A��l�-�i"":p��I�}��h2��j����t�}s�v&���I�l*;-62u��مO��bR26�b_���E̼�O�E��=`6����˭�h��.���c6x��M����7�_�bd*ǯ�A5�����9]��Z	�_�ei��F^����o3�-s�nQ���Lj���O�������2��1�r�(�?�|�Oc�)��*3^�g`ne@y�I���Qf�˜T@Uҝ�5=�:�D����)�=�OH4��|�ው?�ţ2H��f��1%>���#tq�F! �m-�Y;�lN;���X���y$�*s�����)ÿ`B�2����5�_@�t�÷ܦ6��c�7;�.e*�Z�#0qR��l�l������\QLA��vͦ��b%c���q;nq��ʻ(Q��v�0��aaB6�o���={�^GS!���f��{�������k��;C=�;)<P&R��ic����ay1�S2S��e7iCҜ�����Q�XJm�	W���>�<�E�t?y���x)n�\(�#UΤ����G�G�F�/�+��B��T���9~]h���b^m���Q;W=�b���[��Ð�b2GZ���D�UC�N9���.��pZ��M�ϡ(�p{��'\>Vt#�������ҁү��iҲ~�_ b�.�o�D�+��S���[�����*�f�|ɔ�2��l���n'�`89��np���e5d Os�÷HR0=a��.s��>��� $⩊7
��T�f��j��Q���/CG$�WG�$:�W�n��W2��8<�I-����8^Q���fa{JO��$�1:�O������~���gӤ� ��Y�/��>��h ��������;$���Dh�J'zٴ2=������f�祸�%q$�B�(���R�j�&�,�y|A��*	/���y(�j���r51Qi�ϑ_S,J�W\!���kϖ�W�R|m�&�n/]��Weœܻ�w�4�UE�{B��љH����R+�����������ǡ�gá��(_!�h�@y@!�p	V�p@s�����(1t���e��V[�l��Uo��j�s*�GbI�3A!�0Ä�4q��؁���t���D���
���&l�	T,�>��w���nw�K�0  �t�]K�.3z�����1)M*�Fd��.��O	��70P' �Zp[��GU'#QC��3mp"6ٲ�r$ĪR�4�P �p��G��箻j�@Gl�8x��%�:+���T��� ���m��,��C hX>W�J�hN���ex_���l��o�쿕��G��l͢r�.��,8/���Ϛ{v�>aÐ�W�=擧d�c6�@��<=G��O�4��]��L�dɅ���c��8s�8um�P���hK,>���ϑ�\�� �� Gռ
D9M�>�L���C���Uɪ]u#G��/g)ۋh)�X��R�LŜ��Z�p���]�h�8|��ͺiz#lN�����&�22�/y��:�A�GDHQ������	��ɢ${t�8�j%����~�bF�s�0싍�'�a̓�8�#�����4��o�3Oj�}�K��>D���<}�{1�뒢Ҩ"z���b!ٱ�Sf)��8�X�'Mp\)�'����_5m����l�#bI,I�ʾ�Ű���^�JC���}�"���f:�Q�/��l��*O]��i�#?]��싶��B�$��v����A�6���@��9��_'_�'Wl&�&?3��GU��l��&���kw��������=����۷T��˔�f��V��|���Eʲ.@$��Q�|`�(�{\���%��_(ID�p;ǣ6�/�K,�ő�3^�{c��1.��Q�z��'�w=R�?��0w�r�F�"����QcF�n�XB�qh؁@q��U���c���{`-�NiaB�Q���>��7�䳒jP�!Q��G_�#���"8Y����kp)�J'ciU%Þ>���ĺ�?�%3��ի�ILP���\vF��[:
��˺�0��nf)"�MŅ�73�1����H=���qMA	y���Q����-�TN���l=����mg}�!�f���b��A�POEw:����3sS�]ƴ>c�*��u**F���R��
�ԂJ����Ң}���`[����!Fn@^-�<�?+ʨ�kӗkyOf� �T���{+Z;`Mmף`��YWk�#��� }��p{����ø�H	��~u���8�L����uR���=m��G3O9&�
�����1�I~D�f�}Ba�ȶ7ਣ���Q��A�v҉��/�p-�q�6lgI[@��Y-�PmfЯ3^5K�(˱�Q38D�J��W%����m�����cb�6���Jf�&�.��Z�gh��C2 �xvQ�'C9#M�g�B��z?q�E0�Ǫ�K��.�/�6�?�&0O�њ�d��l&7�����q�ͺp��lq�X�V�<��Ϛ�u@�����g�'?�%
����;���_�a��d�u+{�����{P0f�����G_h��_5b�6�b����9�;�[��d��91��]��3s�[����^T�(�IZ�5K{�5�|;]BvH�]���h�@��Iܞ5��=[Mk�ƞ|D!����j� RyE��n
��=�"ep�!��d��İ��8�J�hh�*� �c�׳PU�$kڭV��n9��
{D���g��x��-������8k ����F�:q���i��b$'E۫��#�$��ġ�|Z�p:�7qZ�(�-9`զ�����s�*:S,��� m�-�J��LW�Vf�h]���s���7$������엘�'� ��Q��"����3�[�y3������2(�a��,|E&J)ڸ���2�ԔQ�W�VZ�D��ʪ*��{՝���S'�����:��WLۯ�������4�Hzz��1��]3�H_%Q� �@�cC���Y	]+�Y�n�8ܬE�|S���6ܟ��,dvY.�fP��2�y(t�c᛽L�D�O3��g��9m��@�q��;0��哄��������e��o�əy
_�T�\���%�l&'�z�lҦDf �(/	�����W��e��m=��H�!ҠgbPw`��Cr�Ŝ��:��<H�_v}�C�X/�LڳM�c}�k�jQ�9�Հ���n.��9�{.A�~;z��Ly��"tPk2߀Aݝ5�W %j�s]b'Vd-{�J1���eq�N��3�<4$�c��$L���4?o��O�cZ���q}$�	�]���w6�T��w𭒳��q!��׀7��.VȉoQO�;S�S��5�k~���ۗZh�_��O �J��������*U�O�)��Î�������p�UAlLH,ľ�c6?`fh�í\�������]�|������� 4>���F�����M�C�eCi�4���AI�6�]�	�%���8�&o��1�+��u��\غ��N����g�§�M�<��:�B��5�M�s�O`���3ŏ�s�0Q"5]
%�$��Ū3��db�N���y������_�w�:h����_�AI~"�2yO���m1��H�������Y�S�|a�����;�?�ar�Q7��=kQ��� ��Eҫ*������Β���Q����9����"B�1�Kg[
�وh)�d����y�#LJVz|���� ���`�R��Zp��C-y����p7�1N3�Mt�֟�E�b��3�95?q���d�1^>����n�$�e�� H�u2�MϺ?st-v�ET�=��9b7Dr�:^��D?�So��`U����� <�;d,:id൒6R�0R�������� wm%��ӂ��� ��uz#^����Z�_�����\OffI�,�LL��l�i]�ccz=���P�`��h�VY>�@�;�����l��HZ���Y�>������O�[R>u4Y��۩�T�^DN ��mJ@m�	�'*C[W�kh�O�3a�֘.��㔒1[��∬9�70��S\�h�ǏHgP`�KZ�2��G=��&6w�;���v��t���Mz�{����̾�gOmF��x�:4ʥB���`��O�_�F@��s���~j,2�K����nj���IC���	��BN���~z6+@'I��W�P�*\)k��TZ,()�r�_�(��)>}}�bV���K�9j����R�b���W��j�y��'!�.�Q�36�)3����,��C��C U���X�+��Y�A>�R�E�C����a>g���i��߁�YdE�/&�ϱ��2bi/�|R�TQ"GR�?Msgټ>��B³9G��h递�����s�B�-"EԨ�_h��|\��B�؃�qQM��b�yΌ�	�e���`�����O>ԓ���}j����+��V�e�\frp
�r�_}����Y�L��P��O��5�����G��=$�HN��|R6�$s�ƺ���_�c��Cq,9}�ː;o�r�Σ�%����j�۝"[�v��jnd�K�ʤP����I�+�Ϗg�~�7>�BEnW��ܼ�1��S����+˄ŮQ݌�5̖zkG&�`Ė(�PءW����?�6}s�Go����%�ct~y(ڽ��d��=��@������*�����%��%K�\�xŃ]G���C�m��ɐħ�Ic�{��D��q|�>�Ag��`A����Xl�9�6�8`P� Lp��.� jx|l���Ϛ��;:|��#���Bz�W�BG������c�0�JVq�fn�=|���fX�-,�d8Q�sD�;[�p|�O�R�@�g�<� ��յ��_a?6i?p�C�iU��N�I��J)�b$�e��PWn��	��b�QO��1!�lP`ߚ#�����Q)�m��N�A'��V�7[�4
h2'���o�&mF�`�u]{��P�\Ils��\�����fO����U�pY+�*�N�#6f��v����RXG��q��9�f��ݭ�&��۹ö�xq��Ns�P��s�sq��N���|P\aH�ף�i��tF��Wu�"��	�t�;�B+d|;B�ZO7��k��^��	`��dFʂ����w��H��k"�4���.e7HBQ���k
%�p��|���.�j�&�	�'c(]p�G	(�� �	�G(;Qn^���}y'���B�����K�Y	7��6�	2"��#Ƙ��{�Bl��m�e�OC\�u�?�qn;���nd�h6d���^�mb����ϯ=�Dg��ܔ�Ɯ�T��O8R��g	@���7R�Pɽ�Fh�j�
״�f�[�	Tz�+ ��W4��	���Lm�C��Ř�]��^�K)؇.�X'��E�*��O���d��Y��n�b�#��R+F��(K���;J#�:˷ۛ��\�uO٣��	ӄu`-�Dn[��c�G c��f	���))��.�}��A��o�M�;���O>���է���+��)e%FJS�4R�xتU{^(v���68o1��]�w����4���K�����0o\l>���N��m�;Z7G�i,� u.{8��fmA)�\)S�I��	��u�M�5-��\�L;���"���OT a�ҍ�H�ډ� �鸉�������.k\E�A�f�6�h��<\8̉*IOc��<q�y�"�;5kr�D0"�N:#��	���.4��G��Lwn�����Vj�%3>�Y�PǗ��	픰�^o�y۰9�N�&�y���$��8Y�s��Y����]�������("�i������lt,Z��|D.�w��`�`���~܍i���&^L�ǒ��7%�}���ֲ}�?w��mZ?J�K��7�2���Q��+�li�G��v_|��;&���z>���CzK1o��� ��&-\t��<�����7f^؀�nKY�V��fBYoq<��zp�o%�e��)�85� ����3Y�`���{�9����dVf���x�나��ѿ:��K�Aa�t�2��5��"�|ݦ\�����7ҧ97��ݓU�0=В����%�P�j�4��.��h5u�O�'�����#�H��>��Z�����P����#!ֶ�����`���j���<�mŀ����V]k�s욌�]�9[��ZǞH~����K��I}A��7¡�\�
��Ya��u�����뙴D0�!�es4^Y���_LU,w^e!�a��^F� �6�%VXG'��
nD�T)����P���dl%���� ���ܥ�uM08���oe������I��zh�!٦;�C`۸1�m��G��+Knl̖��~�9!ۺ	�#�R��Ug�\i� KAT���;q��3pC��>�Z��O��B��G�5�(�m�Dњ�<�B��j�s�]"�Ы�����=��=W�hn��M0��U#0S�ig&.fI>��F�S��iK�#� 5��&�l#Y>�U:��w�6?�\���  SS�{>��·� {�?#��f�N�g�٭�q��/�fN�̱Au���f��i��d�$j|^���aư=�X~i9�)�����x2��H��)n��)�"k����)F��+B!�`j�� Zn�Z������+�։�
�*�
yBS�'&x�߅ g*Lч$�q��Ut��^wE���<t1�ع��B��}��)k�B*��T�9_���O�|�[��y��fo\&�f�4;���,����t۹��F4���� ��Z�r-׾_�Π*�J�l��N�m��+���];��̕<k��z�*UT�\|�30Yʄ�%���#�=�D��*���f-W��D�������9����_�PAYgHY��Ӕ�!��c��6��op�;?��Ϗ��q%�ޜf��x"�@=�O��k�������f|H�~.��o�y��K�����t���Է'=�_&��u���=�u�K�2���Qΰ�#Ԓ?ܬ��2=dE+�2��G�7������a�A%fL�xzK�&����d�!-R΍N>��足�cR�����@7��v#"��3'J�*C�|�����M	т�%0-5�35�%
?�_+N_�)rJ��/���
�h�M�@�aD�{�,ё��T��[5Rr��&��t"Z�**O�I����ʩ��ƚ��y!�,���U2��
%[E0�[�ѳ��ګj=�:�j�������@�4pZK�8��C�v�fk/.S~ٷ��#��?��~�l��ҋ�>埵+�Px4F˹����%T�r��\�i(���|����N��&�n귪{�LUM��3��+Z�C	�6�g��bέ���+�J���M���)&��>��c�1_��6q{wA�r�����c�v+�fɧ���3��|��&�dhX�<E�c�85A�	�\(mvB5c���H�q����Q{��i�U8���VD��D�أjPQq�A���3�,�;�iީf����J�����M����=�r1O��)��7GX���1jL5���6crr5-�^K��oy�[�Bp��&s�B9L�WGl��R���R��sbO��n�!
�ͷh<�<w,��AD9����W�>J�i��}���m{�N�+3� f�R�]+*�[V`�DA��W"�	��G�ڑr�Ⴈ��L"�Io���g��O6慙��<0LVF	p�ձ����*�*βw�=o<��"p	�W�,v��J`��<!n!��lf�6b��U	��/)���d@��׭Ϸ�C@/��������_�fw�|�c <�?�R�g�^B<�y�r_�QC�w������
	������s��V/w�V�h�Pڜ�|���2�0m~�jJi_z����Y��67B����b���d�y졘�Q�فG�KV3nz�����l=xC�2W<��s$�I���7�h����M�2���X4#�[��!�=r�У6�L��*~q��!���c��A�i��ς,B��I��<���7�f�.���|�Y隸Q�)ft�#��MQ�ȋ��)��
y�D��_mw��;�kZ�fh�N#�6]��9�x\1�2I���k���B�39Ǆ[��t3[c@�^�� �
�������u'�����K�����T����-E�,6��.#�����X�����Qp�^�����U�V*'&.�C���~/H�5\�難��b�[�MO ov<6GI�P^f�� �n�D�Гa�8�3`����o�C��1�6��D3wu�[B	�`�b�>��m���Mc��w̲5�5F>�\�>�)0��&HS6��ɤ*�M��%U�$Z泥J Pވ��]���l��҈���+
�yB��a;���!�'�3�OdN����֭���Z�xh2i����:ݗWy�iKI�.��n�,U��b�c�'���0��s��b��M��#/|�r�:��!�5��.�4b,)�w�ݱN%���$''��tl�=��}�4o����$Y�k��¾4�p_�3�M�.����u��1�ow�$����A�Fs�c����/6���.4�q�nA�[ZX4T�%���8�Kb��_!��;��g6����k��cn�� Zm�YG��i�V�C��L��p�z�	�b`!�;�r��F����|�J�p,���Q#��>Q���=�x��w��G��������6�j|� �Z_���'�����o�n[&�zr�f�Y���>V_�w;$Q�0�e�1�E%��ɳ�]�j���Y^*8S�H}3�a��4��W�W_�=�_�ҹ�!I�H����p9�i`��hvb�ٯ�s�����u�[�CΧ�Vb�p帖` A�z�F����9oO	Jg1��$D�+�Ci'z�qhxcc�h�[Wj�� �xs�k��w�uE���^��28�'e���=�+÷�A��$5�A��2�#��:w�;�Tj����s�x}yXK��<�"�F4��+�������YR���7.��.����o�؁%��}�rd�V��V��$U���}ޠ�_zT0�p���k����X��IUTt�}��ͷ�z�����.�X}���/��RP"?��xGB�JGH{�ѕ~�i�j����7Ǧݨ��9��5\\c��8u����L}�X�)�j�aLM�����\��Ih�cG%��ڒ�t�IPMj�^�d�x��b��o��D6�N[�c���3#T���qx�qi��S=Uc���v�|�,��b�?�L��z9�?��%���ޡf�&�64�����!����h��5�����<+��dgQqD�*�������R�t~���!�"�+Y���'jI�72�'M��z�b�"0����	�w�'hc�Y�Ǟ#z�E[�Y-@]�]�W����^l���C���I`-���R+x>g��?t���l����D*䗀5�<#�j4=���]��k@�R���5���Ϩ��r�b��E�X&����0�v��HW�����Z�+����O�/��1�i	~�L��p�'J�giO���z�t�@ �!��l+zYyc9f���Fx����n�U�x�E�~�(9�V����bj w%!pBצ�jd#��_k�un���~����9;��q�3b1�$��%%�53�5a!L1�տ�����~�XqFv�;=�?�<t�4as��y�������#b椛<����o	g�7�B�^��4,�F�q*^O��j@������zY9.�
E���i'BRA�`fL��l��D���ɻ49��I&ʀĴ挐L��&��"d���Qb���\��-I׽n�o��"���a)�>;�mb]1I!�2�+�1��0�2�gJ�ʃm+{����ҭL=Xޞ`z��n;�nx�v=J��}���" �D��d����E��ub�V��Wh����x��~U��Z_��t�]v���05)l�@9�tt~N����i�0mO��[ܖݽ���*UuŐ3D.�s��il.�+�k�I
�6��t8�,k��N�x�ш#����q��)�3���!���Ο�����(�P9���i�E�Ͼ�����"�>�����i���_
�ǵ���lR~ov�UEA�#G��~�oe>�����-C��� 1��1��c�!=w\T��c�m{�r��庍�p�����mj�F��Q₯�XP���Zl󆌧c��ʐ?c�`���G��eF�YʿE{��������J���˿'9�7U�@�u�i4�*x��J����-���?��L�|�0�uڕ�)�W{َ��A�+k�ӟ�<%W?�*@�Pw>��29S�qD9�)^v0%��~�^����<)�Z��:�E�%s'��R�T2&i�ؐ������l`�l������@� �����M?��yp:E���3l:�WH���EP�tI�!E�1$����[��l���_.���x]~���r��@f��暘~���+�0�Ɍ;8H��0����U�*)*���Iz�����.i�9��$��5Q0u�W(�?G��@Kr��]�,-_�KI�m|�	����}��m��Ri���)��O�˚���ͪ�QX���?c�}�a%b�������Ӏ\xPL�e�3aU�*�fJ}X? 'l0*��翡���߬����,�ת� (�pO�9�£� ��|��>-�$Td���m����,���%m���ڶ������%?��(�u�i���,"�G��lRW��G36ӫ�տ��5Z�׸rI�'1�Tv�kC�ͨ�8o!FnI��| ��c	�M"�\
r�.J=�yJ�V]���v7wl;�����2s�WD#�wߎ �̓�X5L��q)vA��X[��W{�[�(c�[�Uǐ���E
q9��j6Q���͇q��GAk}j��)��F�4�V��$�3�  �8A������k��n���|�cV(�ڭe�B��e����{��p�$�����K�jU�,7��2��G�7�9߬!l
X�)�Fmb��TT'S�)it�٪i�ی	t���=���nCb�ƌ�ӸUI���j��^� ����"(	���}	8�!�"՛%�~�}�xzH�+V	�%�&EV.���\��C�H5��A{V��Ex�H��R@3d�N�㭚x�J�x��X���?�g �%�X2���tC�r�2�Q��ݦ����~�`.�"�H;��v�^��A��+ޞ�v��F]�.�/B��$���&�P1}�������J��<Zvx~7}Gv�S�ԇ��"AVw`_��t�����w#:��ڼH��rP�ZZ=���0�X�т���g�သ��~F h�D�����K2���v�HҜ���R7L��J��fq��x���<��T�R���0�?C[����L����/ ���Aa+s�zC�8�&F�8���e�E�7M����:B�b˜~eV��L1�X/38�y���Vg@q�Y}�Ri��<�U\>��B+�d;	�N��� �oŉQ~�W
�ґI���x�-�	��y�f,�
���[Y�[���OR�S=��هr~�#�VJ3nUk�J�k�a���ч��JJ�i�	���KX�7;���ߚ�?��%�=����v,vq��Ӕ ���ư���s�WBh&/��v�f��(�� w-�s��'�c.3���w,�����M��#	G �s�JV���/8���^��0��2�Ѡ����	*��4s��/n_E�Z0J̑N�(��g���`Is�7�d9G�#o�s�+d� ����Y
�Z`�T�o��XXFr�g�ī^*7 �3�֤0����F|�g}��7�6Bw�d����i�H����wj�,�y�H�Q)5.b��8�����L|�R���/�� 1�Y�9��[W����E/�{���M�J
&rX��v��rD�T��`�0N�1N"�W3a���c���b�[,#=�S?2����-K(|:X6��aⶃx�P-�����L0���6���DI��(+�E���?���
�<��u�'�@�ɏjk���"��h���Q�-�o�İ��68eb]�V�¯�`8n�E�{�W�J��3��/�w]�2�ٴ^�
�s*Z}c}��~��n�c 5 Q���>�7�l>�%�F�+�UA��a��c��I�U!7{)5n+�1�S����舕�b/��FK�{�)��oR��F:ú�[n�*����IQz1���"6��������H{B�X�nU�e�����9xx.�ۢ"V�'��^�jY\�e
�8%d˨)<��k�i�}�Im���0&g�φ]Ƞ į�a���R���/yVèWC�\\�fM�k�C�<��I�&��VWϪr��nL��1j�du
�./��8�,���Ƣʲ'l�./P`�C����uk�^Z��;	V#'�?����R�N
�TP,̱�������;�cHrə@�U�� ˼�r�L�ͺ#�IN$s�HG��.:Do0^/�^���H����T���>t���{,(�����v��6�!�n/{�F҅�R�G���Q*���|��4.)I�%�J�]�W��_	D��[�Vq�] @��!k�n-�[
��5�B?�!*l�B/�T��,����7k��&~��(k+G���c>��?�n��W܇}
��q�w���W�^؏_+���N�w��'Q֝�{�A��|�5jy:G�d�)�w�]�֔��_É~��0s�����C� )�b������f��w|�������'��I�z��ٜ=�|, �
f�C�؇����в}��)���?�5�a1k"�-Gh]�!<{�?.��Z�C�h��;�D����#�]8d�d(�|h3Or�`��bσ��f-���ׄ��]���r� ��TM�t�(�Z���S�w�1q��3�d%�;5����9��4���ؿ�n3��ȴ�~����@��#�p�
*B��m*���Y�NJ��3I���J4=�٧)�ݮ�F�	}��]�^Q���f<��У��	��xC�����g�iF�X���-��y�5���֧~���~�Xκ�ֈ���c/��{��]Gg�H���j.��(�o�S��~�����֐L*ŊCC{���a���ŭK;��7����P�|T���M�"D�%�7�?L,`���d�U�,b�0�����ҍ �L�qX+E�$�y1��������&o�0B��ST�Ox���H<?���h���>��m�plQ�lZʽ�#xR0�1�4{�XbǶr683��a哀
�j�S��J����֞��B�Q�-�(�l����[�����y+3+&ZN��O�;Ik�q� X���?�f���U�ey694�{��M�yɐIƊ�<w�c9L2c-0��6Bg��J�C}�QTֵ���*sYf�q��x{_�}?��?h�!�or�/�»Ƕ^a��qhm���^�ua0�N�׮��Y�7�!uUD�K��nm�*[�rв�(�!w�7ڊ�=	i״ta�@H�\��޼���v{�0~�_�C�"�({O��cNh�	�(��E������.��`{�������q��� �uD:��f)j���=��ҙ���3>kvUhnaZ!�Y-�tSS,��{�([3z�[�$TP���^��D���e��3��e����Aw���${I�Ig�7�
�'LV51��,R��ϴ����|�m��Z�@Ȓ��\�]�eCF
��N1���r����a�:\/細Ì���Ԙk̍��V�����A"����ʈ"tf.�`��t���kZW�䡃�9K��	6��>ܝ�5�šn}�i���J�7o������4w��Nrʴ�[XW�3�ѻ#��|�m�;EQ��d�|{̆���k�t(�ø��O0V׵?z$t�nE0�� x��2�� GQ<��)	1�~�y��ސ���5����"�~-����J�N��=�l�e�4b�-ʷc��������y�T:��|-L�����UKp?�ʯG�}�k���N>�M�O��p�qË�c�8ȟ]-��٭�G��2:���F�eQ�������xM��muf��]c���6�(�ѫ.0t�4*�E;bN��^~�:�|(�:WG,#��i�(+��[A����Zm3����gV.Ӳ�\�����dڒ@��sw�Vk�qw3�G�J����-���	��n�M�!��j��xg��n�q%Py�>��/;hz=�(�[�ݠ�D�wK�>��M��۞jZ��[�7�*X�%e���$E��<7n�b�����-��(��!�&룺M�K�TI�U��Q�i=�ܱi1�,)>5���JB�e�6e���"���)�eE36y=�c9*���7�4�<�n |8L���W=�훳���a��`o2���۩�A֛Ե=r�5��A���Dv�R�|�na�^Z����t�v�{�-�u˗.�����pا}�7�&��[�� yIU|8{J��X��H�}d>�a[\��
��h�kmo�(&�O�3�k��Y)�0 �є��Z�K���!癘\�K��&�K��	$�������Z(}�d>�8�Y���z�zt�ۂ��a(��x:̆_p	H�LC���hkE����t�A��أj^|UG@�ZF�j����s�jB�I���R�D��+�R�d&���Sҍ^"�8�=j6�]Z}��6JO�y
��F14?$0W�֟)ݩ��ci9�	c�Fv,�Ɵ��Swqx�n���Ej@��E�+FB��I_��s��7I��A9~N�Tk�SVv��]z�eZ:_z�z>1��n9V�*|\�`��v���y���p^�D�O�A*w���C�QY�{�c�{o�p]\��OO}�eN-���T�|�,誴.յ�-�*�kx����?��� l�4u�����&SgR�(q��y4"�#8�,i}S��>�9�c��]�Ls���H���v�p��v���|��4�Z�$�6)��9��KX��8�TKèT �bֽR�\��|��#��5�;&scO,w�	�g��1m'Aj$���}���\��'.�0� Dx[?Ư���wJ�_]��'R���Y�1j.x[
$�>�T9�,��'�m"U(2��q��
	괍�bX�Z����:3��|]�i�o�� ��Cb�����[Q�Q�>lR�t�A���J�>�tc�B}x�� �=����Z����%Ͳ��bx8�t6j�*�Y�AY6����_8�z���QP��"L��B�	yM��Y���^�X���t�ˎ	{X��Y��`�K����I«ܨ?��� �ð"�h2%���$S!��C}�a{K2�
$�h�
RY}r���J�f���A���NE�K|'��Ξ�)z�Q�H�������J�M~E�"7����筩����3[�0��@��;hf�ML���Rc�U�2j���kt!h�e%���4gM8�c7^��d���l�Q_�	-�4j��~����_�T���ëOq�#5b���;�]�L7���2�wF) ~&�]���B󌘻7
�}�d)ޏ�D��c @Lf��9�^�ԃ�P�b[g2�5sE��_�5�7�V�˃~�U��Ih�;C���o�=-�.[J3�����Ϝ� �~�4�)2�
Z���;�]�	(i��7��}�O���=��F:�-�m���H���U55$QJ�Ԗ��l�P�HTqz���Z6%�QT�s��p�0�%+hP\���I��yl9�u:�ڲ.�&��n��IC��ް��h�9�K^VHF��X�H�u��E����G���D�{��ۭ��[�"����U�<&��%�CϞx�:,f8���Ӓ�y�`�ߡ>c�$$\{���1B�)�=l�d��^a��(����ԱH��o�\��?��&�yz4H%g�Ϊ��#D2�]M��h���n��r
--UF*а �Ԋi��� �ྼu�n'�=���,_���� ���:��W��N�5�����.�_11o(��qv(zaJ����ia�ON䷖K����C<R����S�8q=������+��`�>���"���>{����&P��(�0?Ci`[ ���Aj$״����T���8j|��y灿����T��Ղ���%Qd��lHz��>�)�/=bo�.�Ѹ����
jg��H�B��K�]/��.֘�+�z$\s�C�K>]X1@7�)u�L���� �4���ߟZA��� ��Q������!b*�6�� xw���P��X�a41{Y�n7�v�,���\��OP���Uh`	������bni��w]d���hQhg�P�+-��kN*�
������{�&�E
��]��n������4DL�OЃH}�8�N.���h���*�(
��{>(��:ĉ�� yJ�Mӭ��=ۈ�/�}��M?CI Rc���us�2��fm5n��(�01x�C�׏a�/��/�dj�	x�l�|��!�e9�����;Q̞.-}��_9D�M�(I���#�7�?t$��f��N�ں��8&nD���r��Nf��뉰�g$N�◷���UŹ�����]�5Z���'�?)c���' �hR�X3dy/'t 仠�wvB_�U(&e�`5Y�:&��eQJ�P_��w�֩H�IN�ă"i�ҥ/T��o�M���g`%����`.���)T��c��=hG�lO�2^�\j�B�������
�3�NHz&;s+E����vA!�J���DA��c�4#JDl���x�_R�$ĿX�7�z��F�`��A�}%C�vIҔ��"�v2
�=�*�\��c�E��
YQO7��7��B��QA�n��\;0�Sv°���b��-�y��!�Z���_?��E#�?M}�{��pc��E�h��Հ�	F�j�.a�[�@��	���&��_��\`�0c��'�u~�X!� ���_�^��<YL�T����3�Ph$�g��`,������\�U����d�~?�;.�cX����q.1zn�c)������:����.�w̆�⅗�S� ��O�>	K����Qď��4LG��&R��@����3�*WW�y�<�8O�r5*K�)<4����d����"��4F��4�R��4���~�K���|�yk�O�t�_�x!��4P7euK�<�	)o+�M���M��R��F�=&rڇ(�f2�m����6��TN���V+=D5��� ���n�͎{�Ϝ��#!��CG�gx.}�&���E���1{4#�5�������(�6��7+�Z/P���r�ݯӝ�.u�Y�T�''�A,gO��j9�<��Wc��Αj����ײ0�L˹N�p����Uɪ�)h/��O1�	��.	t�i�ݦ�$��ws�����}̩�'��!iP9_"��+ <̪2�'�&(��!4����Ҡ�e�7�F�k�w�����#�7�.��s�e}�^��o��į]�rn�)�y4����=�$=�/s��]1�t�<�܌%'��D�)�@YF,�Η%��l��2|��'1/G-pK���r� s70�E��>?��h��jޅ
�t�F�b��.cW|���Gut�A��!�_��ɫj�u�9r�
8Sg���	I�=�W 2�1=!k�n	���5��(�?�O|����=q�����K��]�p�^,���V�vx��2!
}��*�>0��iX��p�5�� Kp�X�9� �"FCv�40�݌���;Sӌ�<�z�ݯ	�(�B`��;�h�[驧#��V��� � �dj� �ّ�� '$F���5ܷ��8�*aG8�Vj���ݍ��cDhOYı_���� �@�l&Z����֕�%�FI�P��36��w``�3���H�g�x�����F�O�E�m�J�X�|�j=H��H�D"��CЍמ� �N���������'%ǧ1�Wv���R�L��$?a��:'F����J�����e�B��sE����z�_(N�_��וy��0")GO���lzW%l�Ɋ�8~�DǗ���L�mت{�L[s�{z^�"9:c��S���:v��6+�#�j_�ʌ~(��wE]@wkܖ!jl��k��5ys��fL��9L�H�Ϫ_6#��v�-:O��$1�E</��f���Д����᩷�9t���5�Gu��vRPaα/��)4>��k��%����OB�4ݣ`o�j�{腋Wy���41�����=�ԗ�e�=�D7�œ�.A�k3�j�����:��Knd?��XSo�)��lQ?���V�j�x5s!�MD¥}֒<�"��>
�|�1G3s5P��9��6��.�G�1��{Y�e����{hw}s�B�[��svۉRwG�uy n�A�l���|Z�O)�_	e�8/�,c��:�9�c*���é�v�͠1.����GS��zd�Dn��a���ч��] E��K��]tդ-#�:f�� 9��������d��}gh"�z���Ğ��%�mJ��Q9%Z⎲���J�8`	�/F@1����5��>��C�$e&�>4��|᎞�6���S^���]-�'Y�v��2�p�Į,����YRz^w����8<��Q�إ<�a�q�/fk��V�܂�&����~�z W���KԠ�U�[Li1��ݛ��s����"��t3SSi����O~�+�}��>�@�c!J����V9��b5�}3��Z�m�Cj��w�MrR[����͙Њ8ő�K�V��ۙ��N�B��W�&��g�\%9���7-1?ڑ�wMJ"I�[2yz! �@	��i�;��CvńN�R�-[��	'�X?�tQ����g:[���D������[& 2��U�L�t�d�q,�m�o&��X��G� j#�+�0�`���j��$�Ʃb��}�r�l/���N!�q1s?�0=r�e���>��C����F��"��Ʃ���#i:r?�`�/鿕�0)ht
'<6K 8�DA貚W`m|c����sކ�(��)�T�1�����0g�"Sl0�$t~��u(�EeK0��+c�a����;g�2A��$P�<��� �4Mw�;l��*74�X��q�"�Nʹy��:B�u3�������9��3���~ �]ꎑ���!T�q�;ge�a�>��Qi$;%U�_����.|:S@s�ԗ�vWy��`��'0��>���˃�F��qi�BG��l��~YX��ʫ!,گM޾�7��T�*1�Vx5Q�&��u2�ǧVk8Oh����݈����3F��?ߗ��$����gQ�x��L2`�� ��Ex*X;9U@�7<�;o�ܾ;�/׈\��R�Β�r��˻v�<L-j5��
���֠5�^5�����{Q`SV�'>�$��r#�C��L����
�|v6�Qq�b�&�?��K�v�wz�1��!c�0�SwT��T4���o�.��bn�hlh/�OE���#�¼S��M
�b�zM������K�M	�<�Ǟd���R�f	���*&]r��P����S�2��/����I�o����W��&�p�L�Qۊ%hk"_�"�M������B�2܊T�!���d�T��8�˄��i1�0h�5�9����dޛx��ȫ�dY��(�Ho�Ge�6lf��q�]��++r{�o|� $��5�&����Y�1���U_c꘳!�G۸�KH+.4ӽ��Ljd h7��\������wg��J��S��}��J�v��a�[��,'����[�I,�=�y�@D�� ���?+أ?�~����%D�'��H_�_q(h�W&D��E���A�"X��7"��@i�iY�UZH��02��Ø��d���3B��?���[�6�@�K[��m�����	�(�䴩_�x� ��:^掫���&�޷\Gt��ךP��>z��|'\;E�q�ƗQ�:o�!j�������"�G��rG^��S�\̎�q��L�(�n&�Ѥ����5[�%���5�����д
𩧄�bu��>'q�˴��-�Io�����������>Xa��;R]rm e�'�T���ť�Uo� �n�9�%V���2gw�{^�o)=�6�:�״,U
xڏ��Q�����W_�xܶ��(�^+Y��,U�B���vy�K1����q��`w�K��z���V)竄�B��&,��tc���U�m�(1�,�	c�I�R[#�m����Ob��C��SP9�=��ԛ���Zwl;
GLωJ��ܚ�R�QA�d��5FC�r�M��.�����Vx����ms�������Wb)�}d�t�U��|�H��驷ۦ`�J'���Nr*��,�q�r}�2�M|���q���֍����a`�#�N�(��3xI��Í�kyM*��X��� Z��ߣ�2�_ٖ�	Jp�Y8r��o<���a�C�>>�Ÿ�axʂ;�%�&@W�M�s�f%�6SR;h�AVoA�}�Џ*2(0�1g��G��A곹�Bu��C��˕�C�6����l���3\�qx������bK]Y���M�B��{ *�.�a�޺�� T��4�߀������c��?_7dc�6M��里|�
@�����w�t�G�,Iq�����Zm9����B��k��"�R�Ԣ�~�S��s&���n�9�5K�Ph����@����rr+BŠ+u�i��G����1w	$�^?���?:$��n���m�4Ú�^�7y�c#+J+��K��eE������O��?�Xf���h#��:��Y���ß2N��E����
8��ik�Ǖ�Kc�+l7���^�ReD%4�v�����Q����X,W�0���x�U���x���Z�cP"XF��P����$�Ӗ`�|Z�����PYjݘ�&i{�sK	|�>�fY�d��*�r�jk-�P���K��.=�8drRМR��C��ld�^)�φ����{bs+���ћ0mE�(1j�xiX2u�壬�j�AĘ3��m�~l~�L���Ƀ���/��/+ܧί�Bvs)禌��_7��MY-���]�p;[���N�悼����z��"�$9�Bo1$$����L����������1��V������c����<�Y�.�r���ю��t�˷��Py�[ �g06# 3���d1�z�E"t�9����=����7;G�e�
6�ޙ�������Ӧ�pş=W�;R�%>r(6�0��	�?�@����=T�:�Q㸵~�u�����bP��R*mùlRw�No_�:�1dC�p��?y0d���b�+��l8Ï�����f���`�+;H(T�w�}��3j5u΍�"����e�4��=D��@l�I�5��S.�{O��IDU���s���l�A�9��m�8�
/}s*um.��%�Ќ5�2N�1́�ٿJ��'�R9
�x��K��)��i��8�(^u�KO��یH����X�6Eڒ7�����iy��}���{�n4Q"	� �VH�� S�X���Kv��忉�t1� ـ��"zs��.���F'�59)�x��ꘌ/�	�&N��Qs�zf-S$CX��`ը�A�z�d���]���mU�v>�ܴ�/\7@GO(HȀ�pq��P4HF��M��A	���/1b���Z���8ie�,�VP���4�-.耇!ԙZ �.<fu�F]�<��g'N�����S��O�t��ؚd/��4��/_!Ue�`�L!!Ȋr<�@�z��r�&?��6Oy���&Z{䅭�񪚇���bL���`�ysꛡ��D��0���k�����t�p�}@�èd�B��K����}Sn_��:�>��)��gf�P�=#�˞��:�T�f��'M]l|���`k�?���˻Z�h�]2p����,`]���j@����:w��e1'aK'�7P��e��Hkw�ߧO�K���T"k����s�$�<V6����K�� x��# Sڀ	dz0<,��.>��w�
��v�rI�W7_x��y%Y��%9%�q�N
����{ٵQ��U$�6����Y�-l.\���޿���] �A0e��8��ߑ��A[ꋄ�ѩ���)�CJnqy�������?=���q��S��Q����d�>s� �����o/6>��I�M��"��f�b�R����Y�
m����C�?%�ҀM���;B��u���x�/p>�"�O]�VڊJƥ9}P��`�k:+(v�.�TJk����J�=�V�~攺�9���M5���F�;�9?[T�h���Mwj����O�E��(��� �n���$Ş��	���7Oz�N�ű U�Ǻ�X/ln�l�9�U�*/������"�R��ڼٛ�AS�=�7����V�2���eV��tV*v�x��wь�	.�E]�1�Du��^�i���v�LBr�|jS`��kYa{�;r�Z?��홇`�Mx��؆@U_��!z�_�C4�pԯ�q{'Q����P����|�׷QK��^�#�]��Bf�~��:����6r��$��Ly��*�2��į��De`�x�"�F�{���N��B�3�M�^$�Mu�8��n9W�P�j����C�ߩ���6�b+Ƭmu^����q�߈���{;�,�K	v/vU����2��#���\�σR*�k�s(�ڰۺ��E�
'
oo�I&�#��v��T����	|I'X���͇^���7M���ف���E�x��(;؞X�gbJ.��P��;x��K���q)���g��I����!�l�U���<'����C?M<|;7���z�h	xv6g��uу�~�Kj��q��xOf�'�|$����i� � ��8(�f
�B�9zI��XZA�eH4|���+��VK�]8x'���	X����̀ĺ��롔�xsih� C�h�1�E��{r�`���gF=�g�q��g��t���8�$L"�h�/Cu����;���0b3V��w�7�kRu��L`y%�k=��V�MQ�d��ο+�+$�����Kw�\"$�Z�cZ)25�}�m��� �>0��ć*y�1܄�X/���ʻ^.�?�l����L�Q�LK����W�G�"a��j��)|�M�,r�s�z��WgI�0�n��W���{���O P�W�]��A���yԖ��M��:��#v�ÜY�p; J�<�����y�:ùd�b,��}a����Z���lb�a��R�Ub0�O�,�xH��^I��cw�ak��2��q9��/�Ym[���#�ߢ��^e/̥�z3�d�/���fÇ�) ��I3���L��+~��u������9	V%؝�O��v|J+�	&��&W��l�:�-͉ϙ�r����R3[�
Г�PD4kX�ݎȍC=�C@L�� ��$��%���=���l
-���=̡�H� �D<� s9���1Xe�����X�W�Q���BEM
VVy}g2ە�s��3v{ ��ۺ�/w^���L�����5T�V�a2���ߦ�␌�Q>�̓��R�R�-�z;#W���%�,5�Y|�vB�������x⶗�ӿ-��9�'���X��k��y]r�V"�7�u"*�;H�!?�������#{�^�Uu���s>�_�`������j>>�.�d�/E��W|)I	kT�ۿ�ZĎwj�#v\V�z�+ߚ�ſ��P�*wR��[��+Њ��i�֪�����hS8�7�񩉽`@��t�-p%J�C�p (k��H/����J[�Yڦ�5b3g5��P�>�����v�0����P.u����#5o^�� ��w�'��2$n�r�^?&7�������'_ Pg����¤c=�
�l��'���v�|'mR��CQ[<[k�ddIs�D�mk~��|#��:?4q��N��7WZe堻��y) �%o�K���l�+�oJ�L��Ķ��-)��(Ip���V~me�'^r֩�F���{y�S���"	$���<���E��/ Br�Z�����kJ�-^M; /���3"�����qe��<����~� �9��Х�K��x�)|#/��������[�=p�<��� �W�aU��˔��՝�g��x�����Ww�ؚ�z�y�'�jv�����ސ��p�6&���-Ln��^����X��=����i��L?@�x�e�*�^ڞ_ĨY|�c�wf������/�3�2��=�
�/}=�-��<:���mp������Q����B�������܊Z�&�`-)��pYFI�Y�R�H�_��	�b��5S� �5�22>7ݦv�0�o9�Y'�(~�/	*}�Z�3Y	g���<���$�]�D�s3#u���|X��e<�8*M�����1�Epc� �%;u�:�� �NeӦ���2�L������8��?Jw�:�O�O[�ۑ����!��X�ہ�l�P�t��
��� ���Q��@���&�l�/�Hj��Ή�p=*i����>$�o5?���ҬZ��3YE�"�~�*Xy��Gxּ<M)�U�.��}�������� ��O�1����b���\��n~dtj����k�!�
4>��(ua�l���0Wu7܆�]���3�q!��7��$|��{.VB}4N|V�9��0�{�@��"��-��q���#�X?�|ut�E�$dħ�%��)k�F�I�������)X�m�E���HX~��i��;�o��;~+���q���_
�����]�y���!c����mR�?HnS�hN�s�o�5�4T�����d[+��d,���}M�j���4�~���l��I�dJ-�ñ�bj%����Kįk��]�$6���p���ؠѳ��Ɯ(8�$,�'Z$L\�h����e��p�cd����\"�iW�sׯ��@��JH�����\*�-�F���&j�xC4R)��s�ZRv�5����Q�}��9gt�9HI�[���.5��ѹ����^Bb��0�}Z�D��Q� ��W�f��T-��D:|��Z1�b�_�������d�@1D۟/�	�����ɫ�.��̪��2��SR7��М�m�:�(Qp��b��S�b�)�.���9��K�Æ��"!�DlX��2d�}�"o�z��蠁@�Bd������ �m�$H]�,��[i�ׇ:���j��_��LB޼P������ ������F�yEʂ�Я�.%�ۯ�z�v�cZo��p��#R��W"0ޗ�i$!@�>M~.���9!��]����zS��˅a¡^��j:�	g��:��@ �tM~iA�E_���%��m����+���s��Ӏ�%��3��)�?�����r2Y`��##(6���O6(�p�d��Ƽ�td�Tf���N
	��E?K�?=����c�+�Q��Mk0��o��Z�۶���SH�l#������Ξ�0_���M�f�׵L��rᒊk:�߮�Z���/l���N?���rf�q��w�<���?���ji�-E9��[�)iR���Y��K� %��i�Ά
��c��5x��e!�7H^

uzX��$\}
X��ؕ,(x����ΤK�
�Z���ً�{Eh:&��E�e�,/���3�4Op14��ݓ�Sq�47d(�zB�YFm��ȉ����1K�OmB�V�^���	
�>gY��ϼ��Lc����-10D�9�r?��LZ�hk3��3Թ߄���U]�2�
T~	~��R�h�I�(Rp����\G�F����N7\�^�Ͼ������J�VR�"��Ż�S��R,���,Rw��
���-�2Y���0��|�Y6���g��G��\dl�ж��$��R9�܍gvTӵ	�^5F�׌��
`�(g��W��:��B.+g���-cs�DZ���1$.���o�0���|������'���V$��Z�9�'��M���!l��Ih��A.�$�h�ְIOt��� �g��(7�h�b�x\�)z�lQN0��X�g"��KH��۲�oٱ��mi����B�6��H�t0����)�kW���a�}}�[�&���绝XNf���Ud��l�zҋ8`�A����$���T���t_m�|���u�Ҩ�-n�}�#Uޒ�&6̇��p�qO"�v	]����x
��I�_*�-�ł�����ƾ.>U���ֵ��j��4�IsҲ���6��p
3����{��g�bՏ"�&����f��!z`B>?��p���o�7�\̅oZ��v��(�|Z?QP���Vs|�(�K���CN��*��^Zj�`�ڏP\x�������-Jn�u ��0t� �g<����]�v#B���k�y��94zd�Tņ�i�p񒎲٩P�R����K��s��,��=+��f�{Q QA���l�d����ف���V�fVG׋�¬]S}��;�4;~�2y`B�)oC����Kc�8�Ʈ��L8�oؗ�p�&�>=����bX�ߴW(EKN�Afww����[��NBd	ߪ5;���	{�i�f�hR�z�<t�0������Ξ�C��M;̗�/Ҩj�f�qpܟ���F�b��
s� %�ar]m����������BoN�[� )�\n���$Ϡ(�7g�(<�V����2�Q	5�b�;�;�M�l�}B���r��������:�O�Mk��J�>��6��+{{�Ox7��MhI�ŰG�m�kY�I�3'�xQ�ןi.a�,+��'�ɻC���Yf�/������hr�����U���5Gs*i=phb���I��p��N<�Ry�S(%��üG����1���b?��Q@����`�e~���W3E�~�!>�x[�1����)>v��D"5@o���i�G���"�#ѹ�����c���غ �vGXK(&���L?j���l�߳��<�������X�l�<F�HxR��Xǣ;�0}_d|v��.|���,���yϏ����Y��8�-.�ps�)o��� �u(+����y��"������r����9����#%3��|�Q��Ƭ��v=h�R�y��U���"�C��0ޝ���O��\Έ3����k\��V�/�*���M"Dp~C?�+���;�g��6��Fzg��3�eM,��Azؘw$�C)ݚ;\s)HzViM�7F�p�O�b�_�)k/kSdh������:M)LBF�3���q'FsUzD�����@ӌQ,99�ӂ�wwP@�	�����=���I�)^i����ͣ�V�s�w�M:���Ax��$�y��BRb�j�@�㯪f�� ��U��Lׅ#��i���L�d�!"!lw{�2��K��f�{��Z�\5&{z\�����A�?�h�z�Ghy��R�c�b?��ݹ�+���9-�>b��jRI`C�g�6������J>�����'��>��3w�f,j��r%�+ۡ��/S�<l��~'�8�?Xv������? OVk�Ng��<W��x��L%|�@$�;�`�?�bK�{D�@~8#Y���c&���P[�f?��o�mf_ڃu��R�����}��<����BҼlnC�l:/�ўH�U3�:49Q�?�_1F�� tHc ��5]��SD�6v�fIr�!6�J ]���寔�L�t�ӣܤޘꝷ�V�������i�n"\rP'픹]�:�$]Qt V�O
���x=��*�
N�J=�T�]�Z}�w&�}Y�v�d�8�t`�"�������"�XU���#��+-!�ǩ��=L���ۺں��_̪�<��m���,����?��O��V��K5l�c5?�D��r��,|) ���n��H�2]h��QD�a���S��! ����TJ������) �����Z�Y�a��d���@�1��TD��!R��.H9��Z_z��{��6�}�0)B��Q�.�w^�8 8�ð�,	����^�:��g�W+7�+�FMѣy�G���&s�����a���N�&�Y�����v��R0���;�Dm:�^K�H��n����:݇��XR�D��k���J��A�2򯣈���W�o�N�Ӂ*Y�Lէm�)�	�)7{���XM�d�߅�J"&xnb4.}���dQ%��XO�Є.;|���A*�<��8t\��f(X3U��dE��pJ�6砯���_���Y9WłE��W_��g@� G��l��V�+xs�n�c1�2�Z5f�O��'{��,�3��\a��{�Q���]Τ��DzC�9o���}�@hOiڣX�,�y� q ����#'��4�!��Z�F!]�$��NRy�����¥k�үז�F0�6��mj���߮��	��'q.�o��v�8��k��}�Q�e�����1��PM������^�,yS����)���[S^�g��Wy�a��wm�|��Y�1�'n��Y��BK4��q����Lm=�'�T�����"�V�=�c�����E=D)��Hu#ƞ��� '�h���'�Qr�A��h�3P9�dL�9�(RU��i*=1��[��\�[}*�pK ���8�c�-ҁ�^���Y���x%�Ӹt��C+�]��˫�z��][���q�7&(+���A4c�G�9G��$��n	�^��x�:��&d���T��eR1G�F\�^S�?NAWN4(~j�f���Tޑ�>/�����Y+8����g�²e������pzܮxL�(��/�2,�ȸ���V�Ͼ?��BQ �'���j$����tT��"����`���Ye����<��	���>�l�HWnl-&+�h�v`wp&�y��@r}�[�R��oD�J�Z�K]�wxP���t��O���&����1���@M�V��|�85�M[a�&�lRX�,���B�4Ii���W��`�A*��������!����b��;0.�{H�����\�ݠ�0Mi傈0�!q��
ǽ�*��I�8�����H��י%�����#��j�<���6�/��=u��M%�r��fv|}�j����,��Vz�r��Os0W1�ɴ�]�ދ��hEU�Dcv�w >ѼF��$X�0�k%� �n��O�%�F����,}qU�YHr�ų����N��]�i�M�@�s9��QƔ��~����Wd��h�2:(G���>#d��m���^~ǸQ\�L[!vJ����p"�)��2A?�Jc끐�,1��k��V���l'��H����b���۴�6�鈻�^6�YL���Z��FS�,Ͻ,G�A@�����K�]T���@�bt`���R�j
K.Jsw�r�?�P#���y�A��4V�F�=�h+�6`�m|�G[ܾ��g�d�[�xjP2�bogV�� Y�E2���nJ�lড̤���!A�G�����
P�?#�C�/�u����@�iP{�^��"���0a���mGX'��W#�M��|h2��ty�+�8�(�6^K������B��<3ua!P6R�@{����t`��[ѐ�&�\���qڄ����~g��(�����~�d�XB��������.��z1�j����03����I:͠cv����Z#a��e�X�@䳌��b��q]�I��MN�ۧ��������t�u��!��������$Pv�yi��Q;��)8A����vp�h�ϴ:3tJ�9-��3z�8x�y�Vo8�ğn;�X5E�����/j���;Ϫ��Z�j����`�{��.K�Ѩ�w����]O�u���c/���3��_�@��2����^!���ׁtv��'�_�/�.&F��Z���6��Q^�'����FH\⍴��T�Z���6e�W1K��n(�ϋGz{��d
�<�!t��!Q>d(Ny�c��Шh���-�]�)5c�m�O՝�+u%�Z���Jd��md���9� ��������!��W��x�h�s{��m;<U�u��*�M�.4��.�3g$3	9�O�q���T8{k��}��㨏�;#�d���\�,Ǭ�"�W�2���E�# {�sпy��D�5c�N���[�a��ZZ��h�ݰ� ���M������~��&��N~_OAaj���ڼS����
�f�PWz�P��ɧ̋haQ�2��Q|ZeEؖ��~$��%z�M`�������sP�͠���]��?ͼ�3���+��=��	��;��	ƨ$�2�0!{k��I;fv/���`�����hh�)f��
�hoDk���y���j�f���
��5~[M��׵z�����������ʛ��y�� l�zh�����)�n>i�� �Q�����^
:�]�h!	���� 4|<���W9>Ƈ�	R+l>��l�֣�x��/f�㕐���J8��L�`P\���	o��\h�<rR�̩���N��~��2��dH��1�_��Sz���� p��.ݳ6N�'x�*W���Vbx����ⱉ{!\H��X��M��u'㎭�*0M��K�r����k��
c��/�wc����k�*�>�F���N7a�Q�I�t��u�T,	*� �1�3hy+�����"�.uS�[��xu2�2+��ZV��*��*�i]sXd����E/2���ݰ�Bf��dc�D�R��BYT�j?�y���`g��>i���7\8�Q{ф�ݣ�&#I��R���X�����I+�S��Α��{;�`��,!ڋ	[������"�H�ݰ42�ơ 5��l��|*�7� ��4"��}p�f-iy�p�N�+��.H&��O���C��;�C��߭�I։~�\جi�xo�jq�!Ӯ�J<�3J��$�tP���IE
)�Y��TU{��Is��QԬG�[Gp��1���BL���]��@6��̟�����Ȃ��P�^�� �����NV�ϗ��o��g��q�aɽd'��t��E3��J�h���!�:����B��
B��B�ÎOӖ��P������nMS�]�\�0fH�@� �����k*�k�m��lP�ó�����jo�f��{�Zv����� Q��¯�>l��<��;�������K�i�f��]S�6�������[g��W plZ���"��YI��.t�R�L����;�\��~��Ud.�<&�E�gD6HKX�'W���1�S�gQH9oc*7 ���P�Ȗ'�k|:�6�m� k��Y��6`_dx���s����9�`�4�?M�el�X��ci���`,�<�}l�~��=���(��N���	j4s/��J7#!�W��Ј�2��eؖ�z�׋.PE�ĺ�+��T2�&}+#.�
�b-�@�n�Q��<�#p���7�~�E&���5��8���������&��r,�.�Ψ�#����Mkʿw'����y�����k�lj�H�;��O��5]������:��_�z<�|nyB����{����!���q��l��5O�Xm;��P�q��܃"�/0�<�o7��w��HY,�l��"^y/�Mׂ4����nu��YsJ���?�R�G�V�����
<���R'U*��Ë�-j�R���%��W�p
qG�i�,�7�@��5S|��q���V���d֑Hz<��S��F�K�O=o��_�o�"�n�P�,�#@ۜ���]1;���v&vD*��P�+B&��K/�����7qiԍs���m�Q�����zM�~��4����S�&.Lv)E�$�I$0�o�9�q?��P����|�jǸ��Ğ"ZD������}��o2����Q%-�hE�dZ��KK���gfn�]��Z�o����k%'؋+��A!�/](����)����U�!br�c�7WMX�����8���y[l=npbOO�/a�����6'Gp_P%2�r[�A
&a=��j�a�~x<?�!M�J׹�H[O���O���q嗬��Y'd}���~PjM�gM.p[�j�a�KC�B���8o�4���,J>ʡiO��~3���	� q�p<����do�t�5���m�,�>�#���#���M�Jz��m�ĉd�Uŵ�~XŎ���q��yE�l�2͏�3�UW�݅�(v���x��=��=w�m]�����kN�7��3<0������54~K��.�S1�3�؝/��U{��0�#f�ߨۡ3n��D【�3��q�؀?��`�����ZY����1�0�
��"��f��#On��7�dwz�"���Ch�Te��%��� |��q�n��1�j�t�aT F��R>;�g�k��v\�`�J�`�X�nq��/>V��>�lgr�d]����Z��vT�7a=4�@�z�h�;2J`�~��G!������"�-N��z����R-��q��>=W��:�(a#��$�êz!M�Gߞ>��@.Sf��b�Q���l�:�%l-@�|� v��#�~�I����e�Ud
�O�2֍���ih�i�!@�tx����D�Cm����/�jU�y_�
D8%:j�9.�$�U� �"p��K����((�T�`����*Y ����e:�N޲�N���8�|���K�����5��_��D=>�k~������� g�-����7:w��r���i�>த���OOt� �]���������ܦ�/��0�ZVi�Nx�FF�hY�XD�qx
�Q A^�,hW��;�O������h�m�'���3����q�n��<��̪�z�Ʌ=*9����d����]����Z��U���5:%K]4D*�eQ���q1��i�-�d�?�Z���U��m~70_�Җ*�	�"��dD��2������]5ģ3�n�oд^��(���/���a�����^����ǀ�D��Ϡ�:��`�u���~t����Q�����x��p���T����IR��s �����W�b�`�G�yO�()��9;�O�}F��9����^�z���)z����� ����qo~4:��ަx��B:��Ì�}&%p����<Dƍ����g'��OQVaL��7ڿNƈ)~�w���@��/X��������+̰ɝ��g5�����=hQ}�+�����ݕ`��;�Td�/�FJ1Ӛ���_l�0����������ؐY�U��\_�tyּ�&��;���]c�G9�䮒�\Y妄)�vAVQ�q�����N�����C@�=�i͙�wi�DWQd��X�D��v�!+�L]w��i�SɳA��X�F�C��k�)L|!�<�ӟ=��ޫwLW�?/�
<��M���7:��Oz���2rA�]۳D�ǰ;�X=(pIr�5Ƽ��K۝�Ӊ�G�k�P��L����L�G�#3�B��������O4p��q�
��G��/:9c*(H��[+���w�[e*�M�/=���U��*x¥ǃLR�X����%��]5�Y�w,���������H�n�|�B����~.�d�O�$o�f�`6��a��b��M�4X=g~H	�f����4:�Ü�4��h�TKH��<�S�j��-�xJ���[Dȍq#m���T�������[�((�k���/8�1b	��f�.n���䋴�5	�d�n�c&��,���mT�a�H��ع�c�N��]�}�^|&�p����6R����ĸ"s�A/��c�������L�m�� J�*7�}I����#��X'���;D����jV�
��D�ql�hjK��S�����|�A�$�՝�"�v慃�ta���#Ѽ/k������c�~���k��e��r ��!�1邾��E���ҫ';>Ov��B�0�D�J&���{o�q�_f�Y�pE���	�E������?�z1��D��:��b�ob��9BL�|v�T��ϲ�D&o��K����_��w�6���9yc ��í�����oEͿ��H�o��4���q�I����P�(�	�S�DU�ȶ3t���u#��ԉ��I��
6z���'"{�ԏ��&�"���`��8���.�ɑ���� ڌ��G�o�����o �#=A1J~N���L�L��?����1.��[9���!��#ѥ�4��j>q���"�
�=*���_����|���x� �j#�d��]����,NGsj��'�qٻ�ٶ>z*�A^�D�p�$&�.Y��"'����b�,߉D<�9-Ik��N���y8զ�^��j?�(j̇�I*�&�H��6�����y�_���.��]_�Dו~��t�^�ϝ�wB_�K���.E�F	z���̓��νE�D�?lgƘu�q�x����ҡ&�n4��Ghs�aq��#�^��~2��ז�QJ�]L q�}V��T���+��%m��b��~,�c����M���Z�x# ���n��1�:"5��'�`��.�r�W�6zx���n9��2��%����Z�_��I�۰s�L��⍣'��ȯ%(�K�CR0~�=�H���(��*soF��+�^�g攂s�F,DܨX��Vi=L��U~�<i�ǜO{���D�G`:�I@�T-N�Tr��[<��,�y�zv�k�Z0��MP�4l3ì�Bl@gz����L�(S漻�~�3+�w�C���f*G����:%m��2h,t�g�VcL��9��+?�4}޹�� ���p�q!{��F�D�3��A�E��Gp�?J��"�����(��W7��J��r&�.��6� 1�!E�ŉzYN*"%�w�Ս¤'�Hu�b��&�Rl�Q��oA@�.j|S dZ??���Z8�uj�[m˲�>�+�����wXE7mz�#�! A�L�s-A�X�ڿs��9b	w5��qP=�ZM5ܤ�T�XҶ��*��V�r��G��^�e<�[e��&���c?��V���=�}>nM�O[c���cuyiN�{'0P��h�M���V�Ҕ���޿������wH+3~U��>y@�?��L���Pږ�zc��;?�>հԯ|�&�4�9Г��A-�dL:|!?i�@�.�6C�'Zӊ�9~=Ƌ I�M_Q��)(F�CW����so��a�ЛҐ`��;]�@��$V{�P�ڡlK�F�F]t.��dVlΨ�����3+p�z�f�E����I����<+�q�r\&
�$��Ѷ�<�$79}1�qōRa�^���(x�[�k�݃bjCi���T�l���&k>hg^e�N�;aAc���w,�����r>�>�e��qO@�c���0H'�KZ[��ʄ�o�`jf�{s��0Q����LV�ha�M�уZ:�\�����"�ۦ��K�&^3霫��ާ��e'��i���2��A[�ļ�7P/���K�����M� ��V|��ԥ[צ���Ǽ�%�^��չu_����#n2�U%���5�����z�#���?�E"Q]��i�{ �\�tP����Zl�	#����pւ��ԓ�(��7�C_<<�$t��=&7g�d�o�^r$�z������*�?�l��S��K��!\ƈ�Zւm�zM�`E��SΨA*w�EH>��F�O�KmY�ڱ�g��s+��j*kZs��{>
��2pڡ_TFR����<'�&����jv!W֚w�υ��ۇ[D�W̶Z8���ĶK���b�ܧYZX��a=��C�
u�W���M�
#�FRW�&��"g}�❜���#�8����]����ˬo�督|��7�l���-%�+��ͼ��-�#�_�鬎�Z��9�!�����[4���wD׍����W#j�I��GR����"c͌+�$�&�����FNd����u�.���f���Ȁ�Yؽ�xJ�^� <Y���+2	S�t��Tm��/�X��-��P�/���Ʃ�wMR[��$}
KNT��mpC�'�̒U` �kA$	�:��8�M�~f�I�W�5h1	+<1 6T�s�*Q���N������4�]��~0]��vO�A���f�j��,���Ͳ)E�4��I:��s�0����Pa�����<$BF��t�-Dޝ������;5*�AE������Uh�}�8h�N+��(��L��L�� ʋ[")cK��S*������/>��w��め��~GF8��yb�_�u��UfA������N4ʤ��r��4�jw��4�UXC��(���2~�eZL=0�� ��)>���|pܖ}q�K5;IS*hf�He��R��*x�U##Ǐ3�{���P��t�P��5��1Vy��!vE�f����ST��ŧ��[�< �5:a���`a��y���u��"z�D�]���z�HEW\�� ����nT q>d1��ª�iA�ɜf����$S��<NwЊSVwg�Tzs�gSދ���K%=��	t�w��/���\��5sy�"�!�p��*l��v�D.�_в7ϯL���b��T{�;DvaK�H�[$�붰){VGE|���%8D���c�=�44�P���?��8�]���s���'�A�q�^%����I����p���)�9�Ŷ&sa�͙��8��g���\�O��~
��+�L����0-�{6e}-�0E'�w�[
�ԁzc��9�!H���PT�����B�5]�KAԗ��u���x�X �� 9���q� =>�(�p��t���m	'�����:�����\��/���#�/�����SJ�θ�:�Q�<nCoif4����\O2QRj�?�):�0���DM���b-W�j�pJƂ�o�>;�*о�8xq?�/C�:̫̅����,��CfR
�!d�IG��b�?^_�w������5�5A�L�_�U��C���Ր@��a�������-�+�U&k������+e�3?�D8.(i��A�k�ι���9��S}EY�7O��%Kz�.47��T[S�{܄�毡�u]�Yq]�E�7��'��C"�8�I{-޻j��ilSف�}1Yc-B�= �'-�9xwx���)M��4���*-���X�K�To��$��p��P�^V`�y��������TU��E�(cŦ �%���F�'�w�6��ef��c|����'r���'�m���U��,J�����j;4�K�Zo%q�Q�Nᛌv|nC�K�����U�h�L���-�o����Ni�{��q�3�m�WQF�_В�<�J�?�ZB&���yx��yi1i�B�J��wtQ�C`��A��r���!A�Zs�ۢ�_��x����+ i�y08�X��.w��p��A��7[��LtT>0����|3"Y���	�����1K�Y��Q_��vh�q�/�~�T��f0������(^�1X�WZ��2��!�`$�˻�ݽ��;@�tsv��ſR����f(*lG�X{�UT߮���!A���}"e�ԉ5�"�x[F��G!�k栮�?�I5��2�cQ��u��pŊ��X�*.ى�?����f�Gg�#�b�#�4,C`��9}o7L��N@��CP��՟�a(,��|�o�E�tܔ��`*n�׷�8�_Y<��g��|��u�$���C->�=�܋�0 �SМ��Z�c�=�	�����A4������&���<g��+�s�MlL��+i~�e�*���ڌ�$�ĵ	��
_k�� �~�4�gɿ�u���̨�u`�n�9>vp�r"�|d��x\�ߓ����M@ZC�}�K*���r12�ܜ"�A��k���Ѭ����9_SXT���+$�e��~�N��ċ�ט�r������J�D�����#��23�6��#��ye�<�*��G=�U��\sN���~��vГ#cF�#L{��چ��|13���p��0��Hۢ��7D��;�a _f�z��8)ذ�����g!z�����Z�d	��a�̮$�4�ڸx�,]~!�$���ssw^4[��/]�38��6�E�CLl�Š�����zޠ�A�o*.	(�#���B��m�#�q�tz56�����50��D�ێ	� �2���Sh��G�rXLrÛ/B��ukj�(_�`��0�4� ���8�@8��@� �8�F�(�1�bp�v���>�;���ln/r �+<Ճ�LR�*�$ǢΕ�[�^/P4A�/����Ή�����G���aL'�#���x�NP�K��V.�`�W�Lr6��T!�A���e�F%n ΂t��u���?'a�8�\����4�w�h�v������~x���n�oo��a`Di ��i<��ǈ	�\K�*m|���r�MY
i��T��y&��<i��C��\I�|�P��N�~g@[s�.3���*�K�,������o��������EΫ
�p�\���$��:�^?(y�z��E��*��8������k��i��Δ�'Fx��+o�H���Ul� �K$��9��Vy��!��0���Rͭ0��x&I�RkB8���=o�a��hax�/Tg��wٌ´��$<����+������CnE�F<���%T/���F�H�YCi�v�s�]h
<ϖ�  &�DdrB�xo	6H��	�~K|�F�;����%A�tT �����Gf�]���_�W}.�g����*:)j�ʇ���WW�ނ����ƴ�p#�(`����kfAv��x�zB]~��A����E�P*�����Z�R�Q�y��5�9eiB�)Ό�4�j�Ec���ؓmx߰c����@]N���dh�VI54���n!���y><H�O�V�ϙĪs+�5�E�<��^��z^���5:5�<�����^0�C�=�	�[�ٰ�O�m��Q��$�c�VDzʅ1��O�*ab���x�:��v�F%��i�����J��GE�PI7�Q�LYC�]��Iv�\DE��h4�Aa$��c��/��_�f�o&���#�	s��2����_���\%/���'�n�Y/��4	
�a���'=�~��(7�9G�b�8�����xӪD���ךk��Ϯp��C�B_���*��������v��%�5-�HyT�4��U9�_��u�Zw�Q�n>�-�V��W�a�Z��\�"?�$3����ϭ>��0d��>���(���t�:�r>m�Ф����+���3Z~ s��CŲ�=�k���\���m��=ڤg��	�r��(������?��a��j+�:��k�EEa5������<\�0�@u��z�G�>7�쁙�A��VV�J��#�-8l5ى=/q��ɓ��͇�;w�@���[�a0/m�#[]�����,���;���o ����t�'��%&/�.�ց[�6�Y�:?xu��0���)5�^T�x���?2�Bh�S�[�ᅇ��I�S$�HxMi0j&�9�mʽ�ߚvd���Ww(��U���ɥ�`���3����F�^]<3��h��0��X�]{���5MQ�D��3Zx�k�Z�-��NW�t�\`�Z��]�+�K�bG����� �+�V�VNx�����Ș7��݈~]WA��g��(��)sY�oK��)�F���]Z~K�;��s��'x�.�e��K�!��E�D�0 ����[�j��/�\�y��7�\��í�%§�",f��^%�L^��*���a:qg����wg�M�˱�썯���a~�\}'Й��g"�[ŵ=z��sȣ��%�0��%d��9̀J�tX�����oDȩ�g��Q������zD�Xx�{˓�%IQ��2���U�d��Q�h�6k�aZ�^�{����0h����C�i��������3�Ay�N� ��)�X7���b�/{��m�R7�,
�b�3C } �_�ifo�7b���5-������Y'
P_}���+��֮��v�;�
�׺U�7�q���Ÿ�BL-�/��`�~���/����gq#E���/ ^������]�� 8�X^�휟���Q�ܑ��K�4����a?��s)��mmc94����=��\=)< .�U`C�C��*}�$YQ�n �F
>Ǵ����'��4��P��]�L|�f�[ �蹽�w�d�
� +d,��� �*"U�d�Ȑm�[�|)Kw��v�'e=�	;Eİ&�1�A��du髇�j�Ik�k[���L��������=���w<�� k���=�p]R�v�F���(W���/�1���?P@=
�0p)#���H��u��!U�1+/S�ɩ�n��:rq�Y�M���V|O�����%��{���@9U�xJ�d��{_ʭ��7	��g���x.])�M��{w��`��u7&+%b��@d��7�&�
x���][�>�/h��5Q�B��N��mM�h*�`�PY�Ó���:��e���@�x�D������G4�@����-2����-���K�f�J2h��1��z�^��I�z~<�('L�A�L٘s�oF�L�M#�)`_����Η6��S%�Z�ɆA����Te~G��=!C�H��0�a�r��]0����J�n`�,���A�\_�M�4� ��$:��\�mqN)�6�~R��@��k�I��m�!�Ë,곝��U�-����8�fg;�ѻ���	c��n���Y����BQ�B��[jп�qr�T��O�Ձ,�%���x�X�04�m"��4���$����6���=<MX?q�v�*�Yw��~v�����!i$��	l�S.�F���!�J(���;7��1��o+�5�ٹO;s0��K/�P0۬q�U]�A�Q2�23�ws���#w�T�~�S�T0$!Oͺ_�&�ҴP|�={�5�5$��
��.���C�'�i�=�h �ݺh$U/q�s%\CO�[Sފ"���?1Q\.Dv�^�i�F*XA�9�u��
J&��2Rx�H~G{�7���&	�*&���S;��
ɥ��0�*Ǳ(�T���	�_�Z���V<n��H���R���bE �
sM�"u��u��s#5���"�����ћ��2r�ޮ0g���rg�(^�BTc��C�j�҇��#�����+J )��b������N�y�S��q�k�;���OQݘ����#n�q�����!	��E�m!h0SѼ"�6�'����+���2��}�y�,��'_��09�gj!\�X��b4&<�	y�W?1��5��P'�AM���7����������C/1�	���抻�	닺f!2��O���;�xX��W��&�ce6���� T���-�����+=��H�Gl�"�[M���6:��v��m�}�Bc�dm�P��:�؈��\�WX"�uك���6c�z0����nnW^�l���5H��^z7aj����Қ/ќ=�!�Yx���P1ؔ%� �7u��h�ӓv&k���o��;�/���"|ޱc��@��c���<|/���JҞ��mƒ2�G��[Oxf��=���K�1S���?��ҵ{Q<�f��.�����,����2YW��见�,=Q� ���I��g@XN ���#�C�n���mG��~�}�����gRiM����� �s�v#QY�#�Y�ŗs�Q��"����Ʀ�w���ʑ�����2�+��S���Ce�Twq�(��Y<귺
�ID�&0��=ia�\te�@ߙ�o�a�$`ԁI:,�q��|��'�?t�Y-`�2��Iz�KAqأFq���u�iλ[��)���	<<�k1j]3e/�u}�v(�j����VE�����x���?`M��"��#��j2
9��������H�i��l~R��U�� ��%D`����޺#KK��%#�1r����i����2�GW�i�6g!�M�GʔI{VB�5�|[xz���;ؼ0{�Љ�6"^��)�����U��*$�z��0��%I�	�"�x����M,r��`�?#��'�QT��5\8XVdSo�<�@��1������¼ #s&d2��B d�℀���Ƞ3��C�b�+�EZ��k]Wx��������i�ݜB*:��,��:��l,��F@��уۭ�t'��e����5]`���+IK8=��h�@�Y���Ĕ}�/�_�����2�����,N�I���F��`�b��pܶ=&TX���CWZ��"�T�������?�6�]��_�r����s����[��?廏� >��u`�o_��]쒱�G���ST��5M6齾�P��c��@�2�}�o��λ��e�Q_J��&�Y�-
u���ڔ��/�������!cr��T����R+�At�y�sE��۹`��"��a�)M�pc�V�	k�FȽ�ƥ7Ɣ�z�Ӓ��_��������s���юje���,>
�Bk�{{��3'b^��k��qO���`�E6l�%"I�	����Ǽ�~$�P~��4m�A/s�;n�����c,���к�x{�X�z�16�4Lt�Q�T��+=��g?�WŶ���� o���&�n���2������9��f,���#4WX�!ߔ<'��$�N��qfl
)����Çw�D�W%���2���"�(�>�<��Vh��j�(`D��+�QY��AuP^F{L��0������/�X��G�&����S�Qx�}��>���clRb�}Ѽ�Kg�N?	��-�Q��7���q��&�;��@�d������F"�߳m�����v(#��ћ�9�J�#�W&��[6��6�$2�R=�������H��-�'���	^
�{d�F��>�W��UseZP���/B��rԙW�<����Ù�o����I �խ	J�d�it�����E)�K�h�0��@�>��zt���|)��b��h������H�汰��H�{,�3�Z�b� ˠv��(���6,xQc8�������|~����L��]N���������I�O^��f���H�)p]�5]8��7�S1�N��;)�3.a�;�坰�Y<���y��
g�j���Ik%���4%�ʄ��0'߸^��c�i��G#�*�!l�n��c���"�a�uQ�BrH���ׂ֦��q��geq�ζõ�2}.t�ɾ�nZ��-���0�}�a�UC���IU>~�=�~k�e���n�U����OE�3�n'P= �j���F+�D�n��
�=dNRl��@����!nb��GP��aQ���]���p|\��?��z�H1��^Y���<�l�9�j 3��d+"�7$�h*�-�����F[��U�L����>2�c�B+7 ��U@G�A�`b��5W���J#�F�� ���MVx؁��]Z�+��V��z��- �#Y�t�V�v;1k)�/
�R�ql�C!�� �5T�8 V#OgW�nJ��\�teds<._������>�h�n��q�|F��r���P2R��/'��q%�X���2%Dbr@�	�F�r�*횢.<���,�|��/�@>T��D��-�Q鳈>�?��l���EE�2%^��N�S쏭[�.����c���B�f<����*�������_�Â�@<��	z���*q��A���=�jYՓ�$�I��+��g����ڋ�g���i�IZc2m��s�u���"%���M���&�ȑSj��G:��-���2*֙+�$���q��{{������=��a�җJ�b[@ �	� ����TsMT�`�RL�4��&L���E�D��L{�Z��v ���hn�4�r9�Mǧ�.���97�4�qU�K�+�&iG��V�/={�dS�^�I�ŠB�^�m
��Wh��C�����������,^w�2��6K(b���Q/gę�t[=Η��|���j�	$��������Qc�T��N����������@u��哱�xI?˃]a��9Ή��X�`k!�:o&��ܰa��u��j�� Ǉ��Ffw�d��'�2H�C�Ȫ�Z��ئaZ��dL�m4S��,����fR�C
j�UQ�X{ ��)�o����O�f�pf��sH�p�iG.���M`M�������iU��X�H@0�M���z��#��A��&�-��e���M1W��f�2�]1lM�����y���zd	�P�FL�6��W�����[^G.TI!i%����!F�Yv�B08N8oQ�JQ��G,]��9	�e�X��d{+,�o�d��}Cf�gv����lѪ[�<՚+��)6�����ѡ�ق��h���(��
^,��tݠ�^ء,�XN	��ᥓ'�E�����|̈n5}�J���~	_o���}ܿ�n6k��"B;��|���H�H����{�|o���.u�q�u�C���R����Ga�g�x���=�t�	��9oJ�߯@�1�P�a�g5lK�L,���Kv��0bϥo�I���7�������C��%������6�	�K�5��0�\�`wV�_�Q���O��YtD'��h��>3"
^ˎ����ȅ�K���I�CGS�+TD`�e`O88Õ����!lf��
rޑ��9����YVn�㑮����^��Θ�]Ac���q¼@;u��G���P���ї��K8��	�zB �\��X`�q���+b��/��	z��z=+cT�3��}�+�vuf�h%��5�w>I�>?�a� L�x�����]��VWP'{�g�L!"N|&ֹ`^ ;H�7��}�\��V��ݭ��`];I�h�/$�������h���F�4X,!C�,��f�x'�O~��d~TN̘�^*��<+���U�Q�]6�y-f���+KD�cN*�!��/�ܻ�l#�wwf�H�F��|U��Sc�b^(�;�g�BG�Z��Ҟ�t���!����nYZCQ����lՆx�Y�R6dU������Bl��R�.0�lU$V�Y�Q(�S�$`l������ugہ{O�QL[���W3����R[�~�o#���rQ��qr6��Z7!O����z}�!^M2�L{Qބ]�|@���̳/�o��G莮�d���0��$@�`���Y=ɞ|ݍ�"��D��9C[\������h�����2��LıbXz6�U�
�2D)2�P�x�ﾉ���`T�ʙC�����D�}r�C��b�kk�`yt�U���-��C�:��� m��; 7*T���D��3cۓ�F�e7�>�q	��V�b]��P�����u�N8�e��F���q�ۀ�2����$$`��o������8Z�>0j46�f��v���I�c����_�ي0��xP�(� ��G���V���e$�F��˵j`A+�k�MFC���F�s�`��������8��&�L[ҕ��n������0�=3Q;���D|JԍHH�0j�g@��b�H8f&�'M���{#�	i�]rp�"V�����@��B@����Vi�=�XO[O��PV�\�`�#րS�2M���� �p3�TP��w�B��܋��>���T��P]���G��%�S�hV�a��9��OLcҠ�2��U^��I���)]���r
��;��l���d��~.�'P4�JX�QO�.��S ��q?�!�K�M{ʫU�n^9��jB��#�1K8Pq۞�LЕ=]�ʑ��
��LZ;�kNi��>zx�y��!<�r��c�a��疔ܨ9�?X��Xh�'��h��t1VmE����-�8Y��L1��	2�ue�g����V����n�g�����A	h��,Yt�� ���u���o8l�P��/2d�z�$�W�R�)t�#���"�mV	-��0)�6�m�E�����zZ
H](p�?�^��{�A{#k�K���K��^rM"���^�R|�dDbpiks"n��2�g���� Lf�ӀL�/f�(�����43l_���X�<ZP�Z�>Ϲ]f�+��,�@>X�P�Gy;���W�����Ԡ��u��]$
��%+�	���'n5���پl+�I�)R@�ӥ=�;�j2	���� �u��1H�	�R/Ɵ��x�b� ��S4x��1�5^�YPn3\
�ar�S[;���@r�DYv �I�j�f�=�P��p�;Q����)	��C���	^��#q��`S��r*��<�^������f�&�<���j�
��_��l5cZv<���:/�"L�ۡq鎗�	�"�Du�Uc�O�����`�
P�������"�xٓ���=�-��g1y]z{�ށ`�c��V�$���-�K����,���\Wn�4
M �Ǿ4P:S&�Br$4)�@����:%Z���:�uΎW<OF`�9����G�s)�Y��p��Ϗ}��V}7�A�����d=�'���as��uCçǣ.(�	�T;KI���Y�N����Y��7���Akm��>���KF��>��!�t
'��m�L!�H��imƯ1\/����I��ms��}��5\�Ik�!��z,�N����=*�x����5np�1;O���/1������9������6r�,NfUt`��=է�.� dꡋ�_��7Q}CI�u�p��ӷ~4^Y���A�I#9K�����rK-	 #�@0�$j���	"2՛�5-�Ub�ӴԴ�F�S�->9���F"�lXz�w�k�88E�,�!޳S:x7F�(���5� �ͮ��Y��Y�����?f/����J���/*P���h}\�'@I�u��a
��.HҪ(52Oq��m�Q��I
���٧�[7?B�g=�e�򮅦��ĭ���<|&�(4��l�R�-]Ԩ�X=�!���㧭�(8�[M�����wY��!��JS��8��ĊA�T�f�д�zDJ�$�T��5?W���Cg�E�NN�-�\^��{��T֨�ڑl�$��?��%��Nq)�����|B�JDq[f�u�1�n�|��;ڔy����KE��D��^���3C¨��¶�E�R�3z�U���-v�;D�u�&������6��h6���R�0+�٣ܜ��T�Q�$���TL7��ܞ�������;�"^<1^>��ƭ'ʀ�L˛�B�	�z��[���Ρf��I\lRx\ �Dq�jZ�
ew7�-̔_��z��4����HfB�1�J�4��o�~�@X�H� ���&B�J]~A���FiI���oZ>�X�	 Y����ޘ��aȶ�}��+[^���=cĦ��2�t�!�wa���K�O�&��5�|?��;ҁ+� o9���)ʱ�y�f\Jih��mV	�i�9iŋHe^�В
�ݿnn��zU0;�Ҩ%9L�ýk}�Ik�k�W�Èǲb��OI���.L���LG�ZxJ�tʛ���Z�K3�d2��]<��1=p�%��� �8ke����	��\��ፈA]M��uO�n�e����%�Y(-�p>�.|ϱ�=� >�z�:����ӗw����p������+<�	0�������P�CgU�fX&��M���Iv�R�Y �����]���2	��+ ��`���Q��91B���Wip�D�SyD���e�����:� _�E�G��?�Hg��ݐ�h��*�ν]��a�&QHi�'O�ύ(���C �K{�),%���t�j�h�7��� �:���l���u\w���=�϶���%�Ϛu<�����%3�5���2�;>��_E=m�
���/v$b�Ⅼ�D�8�UV�ǲ�|X�S�*�����R��k�/���8S�O$���&��!�O���:FEH����[._����o�ax���}3�X{wB��y�����A����~	�߉�:���0��I��`_�TVD�48�~fV��"���OB=�u���:�iǶ��#!u��ҥ�v/�l��X��m%^,	XYW���	��cC'���(f4���Z��t��qy!��X��~{
pT�չ}o�W��B���m�}�P���١h��!��-Y�}� �!FH�^x��Q��5+7m��]w�x�c5VY�`/f��^9wp�q8L�84r��1���K|ӹ���5}�|ꇐ@ ���:�rM��y��E���n����\3Lzl����e��xwk#�WY�1�������X�[�9�[)�]+��;�AS��&��B���o���F���ql����F�$z�(H�8��<�^��������	����ZAaG>j�����jƤ}C�s�jQ�u�>� 5Ë���|�ɠ�рF�����A�$3���&X�mM4f�ځ܌)��;H�<��Y��7�b��f�rkb�+L�,������ٲ+([)�e�%�]�~KI0�DՅT�[&��܍�5Zk#�K�t,'�~���i��}�W�zv��� �N�)��}y�X󮪥�;��'���t��)�i]n�M�G+��[��ˬJ]�_��U�w���(�i��
�s�����r���&]�M���s�G�Y���Q[���V�`Z�K�Z>0-�`s p�x{�w@s�,��-,X��hwՌ��~�AV��U�P�j�asc-I��8>�ޅݟK��`(@�-̴Eq� ����Eqzd�2�۾";Dބ�V���#e�*A<��i3�D������������B�}�8��t	ɩ�*�|ڔRj�����To����`Pi�x >\Sd�N�Y�ll�7�n�fȪ��Кt�bբ`.�-��0M��E�T 6�O�钒�b,�U�7��H�������U#��*�>!��zߕ�pV'��v���lQ�{U(NH���������;�����u Y�����<�veC�^�U
��h,[mX��BrcA��#�����Ņpk����8FWի���t���@�-4�/�C;h��������"��
UF��^jV�٣���J�]v5>]��	�P�1�I$��U�����(,�/�������~?���0h�=���֝��v�W1�£�;��%�ӠT�MƯ�m(�M,:F �_S��g���1e�1��KO9H�p���X5�e�/�#��9o��Z��_��5���n%�"p��=�<���1��V#��
��5��"����۵9O�z�[Ɍ���r�D@���!�A �m�Ie3� �|B8���J0�	2���u7M�.|�9>���nr?�&��0�)=�D�ȵ�B��u4�]�0d���x�>\�����)_��ʃ�jd���Xз
L��߯��eғ�I�BFֻ]#�
ݗ����:l�$��ֺ�M�r��[�ج� T5R��:MǇ�)�O�+�Jhz�ij���h���Z�^�B�Fɔ˿��2��1��Z�|GK�vo��1h�}w 	��H��U[�;���}�b�[��%q�q���t� ��+���DN�X�S6�g��EQu�j��.�n@�TV�A�ꡕ��q�O�ܞ*��֓_ҹk����̃�.��轘���[fk�|�x��!��F�D�Jľ�I�!5�C�d�B��^�O�r%��_~�?�x���Zo�uދ�d��Ld����K/|������,�A���2�I��,Ө���1S��>�em��9����h����4g.ތ�P��d����X�I8�y31Hp�1	,���߆��Ym�,!c��7�PF�j�� X���&�3�� �<*�5;j0#����k�y	2��Gƕ���;��3F�_T&7P��#.�
�Ɩ�����v�����xI_���4[Ĉ/*�^|�m�Ѳ�q�83M�Jh$�&��P�s���+�@bA���K�����da	�J���D/S�a_U�<�k9c�@,�,��C!/�+Gճ�h#'_��\ᐄ�?G�;�Q����rR|c�cͿ�E��D�]E����O�/ʊ��4LG�\{<���|_a�CH9�ĩ.�P"��0'tHj{T�}r���� ��7�l�_�3��X�	��+[��}�{{*��m��k�"�r��`J�.�/D٘�X���&�s8eb<�ӹ^	KFV:e�~��
��-�����u�1G�b��ȓ7���O�8�di&A����Uل����_,����)���s4�~k���B�t��)P)�6����=����c�}(��:a�t5T�Ga�i?%hy��tf���T4�45�5��t��~�W�q͝֐#0y>vE9]JK�͇.<�ݺҬ�+�|�ײ�SC �p/��C��惮�c�S"�ǉ��;ZG�@��ӆ|7�������A�l��@���>�l�2!!	��6W���U4��kp�z2YG�̲�`���Xv��;���<!N�8�q�\�B4�]��2d�I'�{�F	����6�����m����1x�Zю��b�(Pct�[�8Y�x�
i-��6v9���u�����R���`X�{I{?�0b���*����oN�>.�	�{����R�nΐ'��A���S/��K��M��t�Ru�	��}��%u$�r���r�hk)�P�DN�D �^{ՠ���67��;�W��Y�W@퉤�%ya�Iݗ I�N~5�i���rs��A�Z`�I���͇.�	���{$�I��m^��CX�:�8׏KC�:����i܌`�c�4�  �`|��=A��a�Dχ��U���}��4���$��h'��w�wf����.��ua����z���@���M�6
QɽHƽ��"���V��T�_*zN^Y�S��7�[s�"�V�����u�hю/�е�݂E�T���ح�[��[p'�dM�p��|^�)�6�Q���cpY��y+J?�2�̠����'�<t�i��?���X �)���\Z-9��
R��4g�s+��9y��R����}]�wϸ.p�>�\�t�#���N(D���<Q�}	�h�L'���MMXzIy���l��P�O-�����5DbO�4��G��:qxbr�	��ۚ�s{����oId�0�����t�!TY�&h����w��i�6������3�h�H�OX�J�a�]�g���@Lm�Ϫ�� ��(��_���L��	�!�2�U��%%=B�mVZ�^n���
�*7X�-" �ӑ-� �1P�G�KU�5YSd�Z�X�gP�1�lǜ�+���V��2������y[3�@���n��z��)��SHz�|Ҋ���8j��^}V2�B�B�B[=������V˚�̉�N��q�/[4L!!�3պ)�u#˷k��cr��L�-��޳R.�I�''k�)� Ep���q�uæ*�Gh��	}j�X����a�(]��Ě����}q��rT��R��Kכin~��#x�9.�A�H��Bn��O��j�g����E�e��g��"%[)j�N�<��ʂ�'�߶�'�v0R��¤�U��t-�v݈�aJ���\�8	���S�Y�bZK���Хu/�����8l�#��9�BxZ�֑�&���tmi�S�j�sM�r2S�:(d��Jk��������e���_`�~���(BBÝQiA/�[�/�՚f��0a��az�>��������'&f��Y�Rb�2늺���7ѱ�C�×;�; f�؄$��I�S����ӣJ�k4i��������4I���
�P�cS���hvoFM�n�G��M�r�I�T����ךVj��h!g�����dO�-��g1Q��k�g{[Á�� i"7?<
!b�[U5� ���M�V��g��^����[��UJH{0{��ª��H�F�2�	�eM"�@POLmMжo��,��]��o��W_��}e�%)#Q�ͼ%����]��I�6��<ɶ�55a��"��xS��5��W��k���}�>&(�.�v�e˗C;��Q��ڪq�z­%e�M�3n���W��sNJk�n(Z�M�7ɤ� �n��:�%������&����{&Q��:��iz�>���\l����+@e_�����������X��^�6���7�W0��bx�Ê�Nh~M�m�K$Cf�N�N��"�q�á"Ȓ_�1���;7@��<,E�"5�f��iui���BGϭ�Y�JR�.1=�U��g?i������"Ӽ'��1�2�o�]đY.q�s�ֳM(��=I|�t�8qXՊ�2�TU��h]��.t�ENb*�rMb��u�y����a��$1�B(���L�o���*EFc`	�j��#����!S<Sg�z�by������Űu&�����F����`��̬6��ڥT��C&/�
��"���+�3cta��qB����v�g�4(G��X��كi�f ��4FK�%Л�BS�T���C^p�8Z��I=�n�4�4�5�M��dȊ,\���y��/e��ڛQ��я�:�%��(�w��jdZM�v|;S`�1f Y�n�9U���K~v�����(��q#����)?mg��G�6�Ok�z�r����{Q�bݫI�Y=�yA� 2��>�,"��j�{�����"��<�#��i��������d~��-���
��]���rO���^-+���4.�	wp���lU6>g�Q�Q3B����f1~h���d������:��Q����o��oJඍ��� r@�.���g��R���Jyi�l�6F!��)�"m�ڢ��拖X��$v����I�pM�Ж�*�:}*L�MECNG��˜A��,!�
�;���U��Bc����[8W;�Iĥ���+!@������[���N�F�5g~�= �}ǟ�g�=;����Dct_���F󷾮�x\�jln(~u���AZ��R?�=�Ϯ?\~�Sv������Y螎���M��6�<Y�?}:�)��; �b-�3�c�K�(b.W\�&֥���S��A|��O?��v�u�k�7v��T~Nږ��(�}� 7�C�)��a��n��;�:�b���H�b���4��(�.|����O<;b��OE��|�YV�/IS	%h/����e�1g�U8�m)�	
�MB<��'9�ȍ2s&�W,R�2{�5�A Qˁ�=sKd�C��<�F�hM�	M�r���S�uK�1�yY(	�䱈�'����4�^�|ELn��7a��Ml�%�O����#>�^�FϦ��F��'-H��hJ���a���j)�u��[\��d�|��N�q� nq0X�������VƜE|����H-UWiҮ:�f$��|3qkB�< !z�3Iz���'�[j$�R_Dl��oe��A� 3�kk�F�݋E���� :��j��U�r�l����d@\]�.�<��������[M�\H���"6��\P��5�Q�e���sy*q��4f�3��3um�]� a���iK����0�f���%cטg>6���P�=4{mKM^l�
=c"�^�1p���Qi'�ϧ�4��"����ymIat���
}�t�Y?��D_��MS�iH����ʇ�e+3�͆�����b�����:�=��N[��/� D��(�Ax�*kTU��l(�s7�C�Rr��{�b��ʍ��5vR����i+ `�|=]�p�2�:#�v��A:'� w"��{X
�t4u�+��j+|Ÿ�F�8��	|}���C�Z0�=b�V�����Kt�XAJ���2ƚ�P҈�n����)�Gؠ⧼���R�ulG�&���پ�ô����Ē�1��f���:��uec��x�Z�6���5�  
��JR	b
��� +	�,`�� !�j��C�6$R�a��%f���X��_Z�&BC_����fo��d�DqiA���?���m�(�	�kg��' I��U�]Fޟ��)=HR�*�_�e�K"L+"8i_>����D{�&e����ܟ�!V2{��d#�7���	�n,��Y��?(�ϖ9D�3A�>-�%s��QC���ͨx��Pr����4H?>?ͩ�� 40��5��@��������t�D�����y�b/lq�|����:_����m��~�qۅ��ej\�qk*~ G8����}���Z&�ue'6~��;�q�,W3��#`�z��R+�>��Ep���y�@�����) A�.�������HFnQ��*a���H#w��u���0��@�ud��\j� h�Ȕ ���0<+<)��d��rN��0�6��Zӗ������t��f�A�B~��27��5g����#�?�q��\bD��]AHlE�ف�Et���ԝR�����n��_���!�U�$�6ͬ�y`����܊;x���nF��ʆQ�D����B��`\�,�CQ���MwM�d��ӓ�UK������� ^(.��y�TIQ:�5o08T$E���d���L�H�0x���:<OQ*�zN�]2*��������[׋�o�-�0�Ft9�����"�P#�OiP�@$�s�Q���_�<n(�˞�B'��8�����M�r,�{�sZJ	����Cf�6����f�-K�0G�k��Ϸ�
3L+���o+Sn��.�q��#}J���>������L7��^jC��&��`��tɓ
#:߭� �.�#\���!)�@3�����vT��ym�`�9��B�.�|dn�Ⳬ���Z_��5�Z��!~`X�қ����,�"�����Rw&Z��Rvdsf]����Հ?G)���n� �j&��Xb!��oj����-oo#1c��t	,B�謦�Y ��l�GIB(���|(���H��i�ᗥ�mq�1�ZW�b��Hoՠ�A����3�.�l�3s��vKǯ��ۄݟ��ݪ�,�3��pi���Ё�� ������ ;A_��!&�ݥ����K�/�?ܠ���A�14+NY���\O�8��1�[����{����;6Lۺ"�P�4(�ZA�T���i�����.��ѵ D��haB��eU9IQK�PM�e��Uj��،MYi��Ӕ<�K[E9�����"t���?
X� $�G k��>Y����G�����`*���+����?%�c�o6v=*|�m�%޿�L��M���4�̹����,,���IR��0���ٚ/��߹sS�N���L���D�*3O\W6��~��Ź�ty�e�I���\�c��d2�HdT̉�{$ɩ���(Cā�Q���I�K�X-Џ����T��2�xs��&l�E�z���=J��l�Zh_��ue�@�B��@x>�?
ؚ0�t�?��|�R�\���2�������!�L��R�/(�kB�~=/j�>��Z�9g�˝t��{+��R9Dw{G��)�۠
�]iKZ5))w.£=�t�v���#����ǋ�*˚@SJWV�w�:
�I�ؾ+6ّ� ^�:�eZ*��R�e��o
��iMP[�C?|8O��Q����y�ʠF�]�_SphD���f�9�g�ȂC��2N��T�� .	[�����M3r��kh6���˭��E�ÿ���NLGT-(CHF8\�BȺ{a�d��e�ۯxd�e4���g����\69��j�P$�#�}B^k��6Ӵ�n����ą�/�\b;�ً����t�2�T�\�5"'`k���g�J���]�}���j��5.�nrL���c�%��g C�[�+P;�aDb��9��-04�7�|
��=�w(��wzw�.E����Rm��ծ�O���OKh�� '%ut�t��7i�΁��܉ҡ��p��+�o�^���	�Z�H\UU��萙T�Bk�Ni���=�pȱQ��x�AqC�er,5�Z��CY	7���X��O�� P��Q�P�v���B'�^�A4o���?�D\�ۚX�T�����+�K8]��~l$��eH����\�ڪ)���Da�aPH?э�+fyh���i���2
�I�j�����-O��]���AN��^�貹6zJ�����k�I��8&�9~�>��fm!=�	\�H1%����jF�_X�ε�˶��ء���4�R��\��Wۮݜ�Q�YU��m�gx]�R]����G`sߡ#Ô턳�ߋ�, j�_;�Q۸��}~�3���l[(
��KPeWBU)��ՏX�e9�1��x��bM*�{d�[�]�P֢J� oZocAR�6���5���|�V
�C�n����M�2��B�S��m+ֈ��ݧ�pk�馛Q9��r�i(z����Ģ	�����})�V#����HJ�?@*V-�T����p�H����1��K��29ˎ�h��fI��2�{��]I����!OD';m�t�����E��Ϙ�hBA=s�)��\脈 0"���9�A�Ϸ�������R`{�>��>iB&��v�P��Q �3��ޠ��P3���i��3�+�iXi~�U�������6���^,	S�����uD�`�^2E�4n�mټ'`�	����ޣ���Il[r�X��	����M�Z��CXy\�0��S�L%���7����4ɚ�A����¢ph޶�����Hk��G��,�@����8i
9�%��*#C{�R7�'>#��`���8Zn�$�O�?MM��a� {�V���/��HB��s?��M),���@����uw��"�Fq
�����|�v����lnWoK �&���w��V���Y4~[Q�Z��~Z^W/؛�.F� �����ۢ�xv6E���\M��n���1�V�gG�Ѓ��,��@ms�jm��,ER�m�A�,�ʷ���?�7n�5!=�����@��מ~�=��]^���e	�}��&r�'�B
��>��5ǀ�<��{���=G�\�q�>Hɏ�}��}[�љ;D�owa��:ȥ�'������LH������`cTN#Lw<A%��Y� �r4��+�.$�"%&;�����Ia瘰/������ UstLK�[2(A=H.h��ʊ�gd�911�����=�N!��qsW��ł�P;��n�Ԟ�xYKF;a��pC�pr�t����`�ɫ(�HYb�-R9�]����D=�1?s����c�$p�k�R�j|�i%��������<�5 6��P��ȸ������C����O_UØ������o|k��yC�k6�	,j=����w$��M?����S��pƶ@�XOL�QuR%Q�"�l7ZF�+�?KU�A��C.�1xc������v�?�/~��IeO�����G]�
6*T'Ѧ&G}:ɏ��>fl��
3syG�A���.�0Zs��`�,��ؚ[d���u�G�+�WL%QY]^V� �^2l�~�X����`7m9)�O��y;Ԣ��b��of��'�`pzj����a��Ϲ��.���J�lQ��CeZ'� $��#
F�+<ّ�:+�h{�����[�L&0�|.Yϱ����ZZ�7�T5�(瓱8��;4����K"��Ӥ<�d�k�)z{g=�v��Q�&�S ;ly�ޏ!*g�Qtۅ����Z�q�����T��&�V[�����h1]?�3�0�n�Q���Eͩ�Ժ��0�mk�V�[��7��$��%Y������#���o� [L��3T�琊b�%1�0�\���Fg�[���&�d��@�z�-[����=��]6CD�����H��ۛ�![vyj%�ʇW��FS�bF�����V�p%ߢR��V�e�!�������	�r�ޭcN�6�"�'�����3�>�у�U�zO�UW�q��,���}��LD�H�3�R��"��K����^��_U�]��x���+��䦆9��	���u�����?��*�U��R��n{"�&�� �!���צ�2�4vˊe�G#�s�w�5������I6�Ͷ|����c��e��]9eǗ�#�ʶ��*�%�ɷNm�ۉ-�����կ(w!{�ؐeĮ�e�.tY��*�ĵE�a�d�	~.�Lo�2�D�.�l~��gb�H��M�M��#���"�XD�6��^C�SģK$���I=.�zo�1�����.b�7�����C�0ڦn;I�>F���VN�"����L�HΣa�jC�RH$s�q5B]��?�.i�mFk*�Z!e#�G�$����Q�*����Q��7<�F~6ת<�]/>��ӡ��ph�S���t�*��v���EU�U��&��)}x��h�	���ِZk��b��M���	�n�!����u�k�H:G��>B��6"d�Z�`J���{��dg�H�E?_!��r,��<�jڨ�G��ʶ���,vcRwC��~&̮�,N��s5�]PO�1�&�=�,�ED���3m������'O9MU�_���[�Y7�V(
[�\�dtdl?�[Iu`��iS�N��G����[u-�x;N���4hpo�/��	�p)���ڹ)D�S��dq��$�wb�_ʺ�!!=�����E8�L���ϻV��$�@�%yh��Ԑ5�(���곶v>OOr�R]7|yՂօ�;�P����)�wWB��%��t�~�X���frmg�,ܽ�:�`��I�(zF�� V�Q�KaT#����i4�)���Pth\��e���Lsl90�@�^���[Ƹ����I'U�)�"��bv:e��ƲU-���������#_z,�9��`܋Mv�g!����2ԍ��zO��v�ͦ5��Ćt�$��6��x���������F�cln^��PN(����r��������E����D���Jgpb�0�u�����Y�6��O����Dg��&#i�������/�Λjy�h�j�6�݄�����q-���0��������%Wd�v��P�0�(��	69[;����ҢI��p�|0�����N�������ߣ�S~~ҩ� ����m�g�뭄���cN%���k�T�SտΙ
�q�PCL_��E{�d���k˞��|&@Ͷ�@0B��D'e�"�ƒ&��~�^�ɉ��xjz^�a�9}$�Y��K�'��y5x�����x�_w�%��oݶ��d��Q$�Y�4s�\9`ȾkȽ�E�PO:FԼ��͟�3Jegc3L�>]0����7��1�@Z�Y9'�+���BVU �v�+f�oUH:m�7HZ�� h�f�Df�y�B���T|E��<@�a{ׯ�7�>�c�d����I2�4"#	v9���?��L��Kײ+�-��PQ��Gm��\�={����D�C�	��$��z1�����j�8x��8~�_0 ������R��F��GS݋���)y|o�Ů�j-����W-�ja@g�PpC$~��[��c�̸���*E�&OY��J��[�l�����7~����L&PI����׀(%�6o�"��:��E�`�ԭՊ#���h���g�m~\}�{V�n��}h�����I�u���e�`�tJ�	���V��HE} ���ǮX������~8|ڼ��~=�����`b�	U�K�{`6�v������t�Ff�[8��Oq�8�cћY2)S\T�0>��g2���)*��u��;��a�f�NSr.���Bs'�ˬ��䝁�\;��r���Zǖ�?�!����U'<[#M�a<t�N�T5�{G�z��(@�Tf�4m�Z�F���XQ.c~we6��_�Pߍo��J*S���a��!��	b�7CD��*�i���$�j;U���ξ��޺�h�NL��a\��}�X��E���z\0r����r]H3}I;�J�d� ��VZ�#��	�9�P�y2Kn���7=7�L���ky+
�������ʑȍ\h��+�_�$�^Wҩ��c&]~�JuNJC��[q^j��S���]�B
������Hp6/�"{nH��v8}��,Ϳ��������
a:�El����,���x�A^�Oۣ[�kxuC�t���4 8Bve���mxOA]d<S!�[���42��'��W,�VT<T������[�̽��^!�xT ���H.�c���8���,��ԩ��+Ĥ��������y�-�VC��Ԩ��2|S!�,������?*��=ľ� Րh�kg�kF��6)��AP鹳�\-f1���?���}<�&���ͳ�O�$�f�F�d�w��-���oq杽��q�|c��!�Ǆ3-;��RK�/�. ��Ty���_D����$]�yC��.(��E)��%�s�ňh���|l0pMT�!�dy-�	����}�`	�ׅ���oC]%�{ܖ7W���`����o!�n�ޯ!�h��^=��q�M�񉤞{%!��1�=�PX��!���'+��:sr��}�wR�؜�B���$"x{���CQ�R�R��o�RK��~�:s�	Mj��NM*�̔�R4��U�zQ��8\=�,�į�pG�{)��iF�6Q8/_D�_����e���@��(��*�4;:�f�o=me��S.>uA����:-Q�%��k�c�G!"�M����;A#1�Ue�]�x��g� �ױ׵$��߈fY."D�P=.B��k\��!y�#�eG	��h�G/?�z�	������s��;�|���z����k���`]�հ���~��袃yo��.:ϩ�u���/1ޔz��q_�g�(&��F��UM�+����j��wb$x�O\���i��"` ���KuJ��C��n��x6/��������-�6�9Ě���V?�\�v�����ȊY��σF�8w��q�%{]邎�ȗ�4b�D-@y0}hM�=i㥾o��8�bNф=�c��ev�c��ʼ	��;詤��'�R����Y���ߣ<�DF��tһ�K�Ug�BA���l�%�̊%�b"��X�W�?�s�;��I,�K�q�S~�IF8�F]FjlN�}�0nz��"1��Zc�	�]K^:�����,�jk��I��H{V�Y/�+�ӆ���;z:MJI3r8!���Uc�Տ��ܝ�ꧭyɤ3?Y��y�G�m�A��*t7+���P�����n	}���^���I#-�Ǯ&����I�-hhd�@���khA������:� |����9�/������d�9U��If�T�����WqTT�.']%S|�V�V�w��#�*=6V���z���C9�ؓ�^�bM��3	�����H�,����'�KtZ8��&"|�:��|	A?�_����OΚJn�㊳"j�u�k	B�h�b���
9"��7ш ��qw�F���c��O�C��:�H��\�x'�1Z�%}��V�̟}2�I�Rvg³ ����pG�(~�'ק�Ts�U9k؄������I��5�m��ƈ��J�Jn����J�[���Ko��{x=�#��auZ�)[؈���A��j�7>b�(��rU�d�
K|��+�߷uW�D��d3�o�澂�~c N񃋃@�W��v|?�8]��gx��.g���1��Qp�1�A�)#׈♠ ���'���/��#	�s�hZ�R�)W�+bv8��#�ﳵyYx�M�Z|�u+n��ҵ6�i&�Tnv��$S�cyq;��fÑ,A9P�Q��n��c:g���p���b�(�z͆�M�u�ظ�ڴ�W�V�p�Nϖ9l�j�5w4�t��/[bڝ�	��S����5FR�,Q3��l�.����S�wqQ ǮT)*��_n�D�͈�d��S�ZE$8ʜ���э��gѡ)e����Pg�vˏ+
Ŭ\��fH��Lߠ�����kx��>{�d�6UP%�6�%���s�l�XO|e������*b$��N���������?��E��ľ5iY$)n�!xa��}����<��u�_���)C��f�l;�S�����PHy�e�^I���v�a��
Gj
�U���Z��}��5��Y�ȋ�=܊9`�UY�<&�5�F�a�`a�O�.j��:Ŋ�M��������g�N_L��2���]6��� Xp0n-@S���º�qJj���޼��+�T
��|ދ��oȟ4]�Ҭm)P��� �������J��3�A�q}%�~cow�&���iu�J�#�7XC1����v��gc{Fk�S���� Q{jR���m{{���kR�wK��?1�s���G7%h���3F:�z��c��v�G�t��b��8���8�|'XR$l�Az@P`� ��	����k��E0Yw�A'�9�T���������_���hs�sY�� ����A��Ņ��h�5|#�Һ����A����o��m22�2qI%���
�"��Z��P��Aj�ݿ��F��;}Ơ�`���]�-��'�'Kt��������T>�y�y��R�? ��!�3��(�!�i�'�a�L�X*4�M5j��D�<�)�W��Y��Ĥ����.E�e��8K���������B��\�A\J��E[�ڊh����Ο��4L�)r���Ḇ'!�d(�;�o��Ԩ�H����Kk��ܕO��w#���K�q*Fӛ:���!�e�9����m�l�S�ÿ=�������-�͟�ķ�jC*�O1q��e��ϻ֍ʯ��%&�G�F��п�?��� <��T� ��Q�L���/H�K��q��m��h��~��Yܞ��]A>�κ��HR^��O z(���g�%�A��wIX����- S�+��փ��f�Ѯ��!�@�d�O~���9�"�O��?!@ܟ�*�����S��.��
A=/8y ��)�v5�:�ٳF��R*�|��Ks�>S����BP4�N���R�x�*8.�Q����H|S~K��s��d�Ǿ��� �sq�� #���uvˏ:���b	C��n�6*hB5��3^9��lޠ�PlD.i�\n�t �L@�е+�Թ0c9���X9����l����l
"R�eQ'�W����q�@������$Cw�� ��.�H<����%��m�׏�VT'Y�h�,q��3%��B��µ�ޢ�i�ba̘|.�[��l��L�Gx�8�q�ͫ/�xƋ�-�63��1e ?��~�^E���e��R��HFc<�F��Y�x���Ŭ.z|Ќ�|H6�`�!TX�*�с�:�����񂎲|�Pb��aH��rH����KE���TW{�#�!�2��+�b1L��Qm��e������@���Y�8[ ׎��	u5�\%��M?�D�ߦ��'��Bm*�=��(%�x��u����CF"�`c�,Z��HqR����*%��^O�ČƐH������邌�Fd�uj����׸ŝ����e������{�����ԕFX-�)ڕA29'2�G+C�U_d�(�����8�WX��z��lm��4�����������'���S�����7,�<]��0��G�N}Gґ.RZ3�$��������\߰u��%7[��Jmt��B�懻m��?�@;�Փӝ��fK��g��՞lQ(�:MEm� ��s�����T�����u����^��|���gJ�fO��7טxҳ��}�o��X����ބ*���FV�m��Iqw*pU���0K�m~��'�Á�{z7�D^D4Hq�O	"�t�?�|����5�1]@��F�ZrBwq7���>Է໋Hg,x�ۅ�/��Z�1x\��w�_�������9�-�1J�`���>������H�	��?�-�/����=p'ROs!o^G�X�J�'����x�9ʞQ�.�õ�0�?�H������%r�y�y�(�$�#&gC��N�DL��q�9r�q�О�Z����kxG�[��X �[��N�*$f��SWE�#l	�c�.�I,�/~A�LUhK��I>g��y��z{j�]p/;���w�	Ε�_�`��䮈d,�4�p�Q
��!=��<��H��f���>,et\z54O��DV<!�������l�7i�E�o���^�s�������^�A�v�K��,G?�4�-64h/@���H)������ċҔ�f,�����H9����k���{����I.��a�oV�	�~�X�~ֻ�b���R�d�P,p���5,nt�B��)�'�vrV�$��>����7�޹����,�}�[<�
��%v5ƥ��R�
��^
�!W�@�`\�y@g�@���jרk/g�IF0^ۻ��(�D|w#cX;��^y��/A����eپ���!�3�ol}[=�����Q�y[ �t��D*��d�H�h頭x"�(^�����3��Gg��)h9eu�\��r04n&�Ť{a,G ���l_��^�M�^�O@��t��}��BX�;��4s��������+�[Z����i��ie&4||��9�H�j~U�?M�v����4w/�bũ�wg���*8�M
L#�����#Z::�Ĵ\��WC�ܘ��wh�ʟ+RU�1{�ĸ�e�E{�0�lU1y�ObY�VR
FHC��)�� !G���n�ݹ
&�Zs!H���9��[���u�&���Y��" ����� ��� ɴ�K{��
Z+�9D2�@�{ƣ/U�>~�������\��֍˘��x�����U{k1�9I_H���s���g�j��Z�f>�^�Պ�ݘ�bM]0&m�����8m�>��p 8����^Yy�loN z�:�(��g����	���ݚ[pn�)�blے8a�P���DY*@X$R��72�J���?�P�<��2�YP�sA�"b������6uv8����=������ɹ������m7�,��/D^a��AOC����^� ұkb��F�x���`�ܓ�pW~U�ߐ���ی��VԊ��������4�+s=;w�@H��|;r
;Z�˓ȭ��cZ	,jb�2�'$�7�n_J��;���42/�������&����]��(G���QLZ��^���$�LŇ����E���bpA�Q{>;h��1�M�����s�O�N{`k8��+�4AE�.����>�r]�Z�x.��	3m��]j[�!͝�Q�t�%/�������v#���j>�c;(�����������ۭ�PV!$$��';FY)�������>��h�TT��Q������$�l^��^ʃ�u#q�����t1�NR�l~��r�7�gz�md�7L�S��gRI��[t��Ѡ���[��yS��;�����-i6N�� ��o{�4�V���7̻ U���%EU�i��C݅��9�������7�J`˟&{}�%#T|0f�u��n��
��6~�J� �8D�	+��,%�lk|�y��=XPH�p�3ݻ��#�u/��(��-�qd���,�Iʆbu����H����'˲͘�G������o�]��h���O��v9��h"��A1���D9:8�f2�n|kM}u��
�7>S�E�b]gQzCg�(Z ;;i�XAZ���L�Uh��[�q�����uw����iʃ`us�f�v���U�Oj	y��T��^��2};T{\}G�}ۗ�P �l�8��Z%y��!�%��fo���G�͏�g���u)����&L�ί̀��T^9�l&�Q>]����f�όރ>Ր��E��lU1r9]-������:c��&TNz� #�?�>�=e2����/�f�������:�|�z"o�\������	K0_��-/,ݟ��B�����]\�S�3(o�;�,�89Sc������ᥧDֹ�����.��[4�w��qC<w{)��Qz��N���d%d��K���}�z.$*-O��%�q"�鋛+j��9�\�{Id\���\�Y��qc�,���F/tj!K<��]TB&;���V�_���/"������饆.�_�]��A���:Nb��i8p���� X{c�"�f��зX�t��Ɏ�r5\~����ȋG���^p��.����y���TS��B�Tr�(xٚ��L��?k����T6)��T�B��uCpS!k�d�T���	|OgY�=M�O�sǦ&��P���GC̨v9������𗵪��$�����W"�KuP��ϕ���?G��>o�^���w4�2M��6^l�J������/,މW:{�hYӼ�K/�5��u5�,EPdQW�B�J�z�û<��%����Cp�*!�����_u�>!�����S�kd#��pIy�幻���!r�ͨ�By��91n�+5X4�B�L�,������B���������	�O���zw7HGj"۽��_�cz��"1:�Z�}5N+4	{5+��Z�5WƓ���×Hi31*4R<<}���J4!���O���T�Kә����b,�2�g�M�6}[���q/�m^2���/����(=�՟f���xJ����Ђ�p���V�s��r��킌}ּ`��ر��o�?�[�xO.��ɹziks���
��褡q���ӱ���8��J�"Ʀc��S���N	�a�JH�W�d�&ڳ�b�j%d?�м��O��v��B)�ҵa&�?��>��_l0]�l ��IC��eԇib�n�(Z�XkDso�g�,ɏ��Ё�dϞ�ѨYY�,.03�4���?%�9��u(K�+�U��P�y*�����9��'��d[I������"K����c�w]�:q��TN��C侴,��@��	(6�:���f&_�ׯ���'���O���e$R����-��r����w��I!z�\�w�7�I�KC3i �4�P�M�:��W�?4;S�eh�5w$��V�w?|��/Q	}xr����}n����4@�ה���_n�z]��Z),T�UZ,>����wo~�
}L��1,�g5�%�1���x�6��-~�	p6�f���I���P����p�t4�Z��'��`1i���6	k��XUVT\vԖ`�j]Ι ׽�����e�b�T����<Rx�Тp�;~S��e87��"!ؕ~�pJ��6��:�\Q���^�Y��R�0աO.A)Ug�6:q�CM�Aɽf����]��
��,���>�`p���䨅r���W�p�4��浅�
'3F��]���V����"ɖzf����=/�^�q�d�\c#�7R����_������r�$Y�>�{�a�]R��z���֘H�8vq��{_�������OCD
�Z�0�U�YJɩ��'����U}6����>-�͐/�*�-�\M�qY4��[Hŵ�l�y�W�d&1HN�$2)�̷仕��U���� A�_����I�BJ�`-N&��)A_6-A�U�j���ܕ��zt������Nq�Y��nq쏞��J��dj�2���t6�{�����g6t�����9r|��+H�{�}Z�'�*4F��֊f�����N�X�͍��+����u��G@����h~"�%��C�K!���TA�6����L��?�#�uQ?Y6=, da��[���Q�}z�t�~�`�����TD,+5e��ep.e���#-�}$r�W�|�X�mB0�-(�>��=�{��#�;'K�js	���yG �s�a�|֡*RFh��)��l�y�������m8��1Xk^jFCHxCb�����UDn�����S��s�Z��O��۟���}*[z;�	�J�i�nY��]�����6�"F��=������1vl�s]���P �B��VY�5��~����O����pi7��ʑ�9�0g���K](��QF/�F��:n��q�.2��s�W��[P5��� �"�W���ꃀ�-�!	�y׾%�0�׏�H���(����'*�-������ &qF�Od�n��/�~����|��vs�W5�d�Ã�hM���s�V���c��U��Ƞ�O�U7����Ex]�0pu-ބ� �A 1 e56��y�ƻ:㤠p�OjNE/w�D�Jj~x?]�U��6��y��q�MF�c�A��	��z�@Ѿ^��+�����h��!'�O�K���|�Z���?G���fJ-��Y�o�� /T[�]��&�׾��1&�ZS��4��SVdO�E�zT��u�5�Q�5�Ē]�CN=�^@L$
5 �bHmJv3n�U�:�(X߻K�f�N#�0��1뚑Q�P�C��hh�;M�ܜ
:{e����F׊����lz�\ ���R����+��gP�]���F�&;���MN�%�p )_��u���O���Xz��H�J֙5��}1kg�ݟ�Ŧ�ȕ���l�����T��.���Ȋ���I���4��ju�%�:�Z��W_X0��V�%YFHr��ҋd�ޡ/�{����A��ݱ�H��������j	%qG�)�ҳ$�'l��
�L�\_�Sh3�K?/=��"���{c#�?����k3C���-6��/Z�_�ԊaPA5��I~d�6�R-c놗U�d�������L��hvq�$�9y����t4'���⑻��pʛ6-�? 
N%������N:��N�Mwڂ8�k��Ư�1�};h�x%������L#	�o��\ ����UL�~�z�xU�!����D~8:�G����nT�O�u�G��Y�8|�H]p��0o�2(�f�s�<�}�*g,b�IɢKq�*"��Gt\��%��J
������L*ɹ&�F�
��&Z^�Ž�^!�J�7p B�hP����Z&6|��R�(��چ��g
��]O�
w�n&Gц��}LǞ���K���9A�<�~+�nJE���� 4֝���MS���8��]0<�����7��"�dn֣fu-�Ӗ71�wT�9�Il��F��8a�^ϣ���9>�4[CBH�{��zJ[�c���X���æ��%�l�aGm��QN�\F������}hD��ݒ�3����մ�Kk^��f�[��6z������Nݑ�\\�;�-0���`��u)d�	x(+��շp��A�A��1���g�b�>�F!lп�e4�R���&p�o�[��xm��eJ�Ѧ�۳G��L�Elj��T����eN!���P�<��LL����F�el}֡���H�����_��Kk��:+��8�-�_������)N��U�q�����#�$�*�=����KQ��i��o/�N��V �0���`�k?R=������7��'|�����^�B-��صQw�Өwi����Ĥ!��D�}��;?��>쐈iz��+�}fH���4�����}TwT(�yH��x�<}�F�;���|�"�Nƹ]y%��K�5S�秡Yr�2jt�ܢB>���xE髙�nn\6�`)ѺYU�<[
Lr@/N?�U$-#�/���<�ۉ�A%*]LG�q6q/:����:�vx��� mL3��gǶ4��v�{��e�v/Fy�.!)v1�6l�Z�=�{��q��0�=`�hs��h�$���]j��x;��@r软iO��U���,�"��D�K��On��0�@ڔT�?r�]�~�M�O�ސ�8���҄���	#7�	� �<�m���0:��j�i/�y媶����Wb������0v���e�`�Ф��#�W��\�E�&�O�n%�Z�\���b�- ��ۮrt��|q���@�W"[R����x���l�'� $;/_��w��Ϭ9��9�O��G�/Zb�����k5�c=mE:0�%9�"&td+�'�Ib|ښ.D��Ub��ǵ_a�p��z�M�|�'ę*�*�T��}N�������܅Pp�8�L��Ȝ�P�.�j!�_,ˎ0�W�|o� #z��l���5�4���V���ƾo��&�[�{5;5��)2ۇ�1�>��f����<���`!�{�5bqX���bc�Ƣk�hm�����bL�r&4�30�u�&�� K�D#7��������}�:�Ӕs6e������!S��οk�kx���pJ��&�kKmkc��;}�hy�b?;��u��8�(�����gy�U�"-�	f�}zJ�q�^ז������" �O��� �*�F��&�˃���zd�:{���Y��Г�qX��p����j��È(n.қ�� �V�E%�E��K�S�TY�U�[S^�E��#���%� �a�(� �9�y�ۇ����VCw_���zJz�*0U�K5���������]���d��\���1�)�����HY�.����?2:��J�gH�f��rG����ɘ��1��ŔGM�
W�1X�������AZ�����@�#vѓ����_yWѩ���s�\w)n\�+���S�Vtt,��}�j�8���@�n�F��հ�a#���5锎3�<�n��%N"���r6�	��&`�1��g�Uf��:9tu�C�B�|�}�Q��C��u�@r��=�N��[?�E?7<E��Ie�F���ω~I�.3Ia}��{RE!.@:H��A-n:q����Wa��+�Zm..��q�-�Ɔ}1^kΝe��w�!b����֔�|׾��TRp��t�r�*�;�&�e����y8=���Q����@����{�G���wXWZ�D��-��=�$���pw��Ud��~�3V<Vz��Si-1�RE>j3�n�i�u��O\�\w�W�r@p��
� ��a����>��oN�w;�ցOF�e\<EDHy�M��̜���)S��9#����df5E���^�F�l�ɘF}�o'Y�XGx�f���$�I��B�����\��ZY~���x���p��1v ��d ª�J臊���Z��0�ݴ���^��՗���WS���4��zUԒ�)u�W~\d&��F�A;��K�����rﲞ��8����+�>[�9��t�B-1�	�?<���}������կ$����>�3�b�P'6�]N����݂֥Ӫ<B
��X�#x/�Ɠ�]o��8[s�r�	�%���4��Mb���[ZW4o<�|�����Q�&;���R|'>&5��|o�b@�{��d���*΂�v����$.���fb��U��>�ǿZ}¬Nv�[PP.]kv��.����F�P�r;�[2��z��u����$f�oT&PC��l~6]e�i���D�>���T<MZc ���d0�@(��G�7/I��"����m��l�$��ɰ*�a=`%�wVZ�r.�O��0���Ugw�*άƥZ/�����|��4t��,�uy ��.��Bm���Z�cl��t���]�E:p�H�8�>������m�'�#�2~^W����F���`�Λ��1n��3�;ሿ�-T|e�f$��	EcyB�d�:���؞�3�<b�d�Y�7�r{�y�y��a��z���<-�lz��+w�P����J
�5����ci�D�5�X��ׁ4��{���)�����\���CR|o�n�(����ͣ����Cc%���=3(2�!"�9��~�(V�g�O*�$����R!�.��<I������bY	�u�v�����3���LI%[n�>���֐�ػ\: �J�䌎3­,'�0���:r�S7�>;���j^���h����:�\>ݍ$|f ��`��"�?/���8��A�d�y.sN�7k�s�P��`{ę�C�-����@;�7�XzTv�w�c>А��`C�� M�C�T14*����V�e 끀 }o��j�5�{�dOcΩ�'H���[��5NԚ �����v�~|��&�{k9[9k�l���Gh�k�V�+fҕ󄖰�=�P�ӓ|�D\��8U�@�&p�`F::W��2����YGUm�q��F8��ּ^��f��^�g�� ��!)?�z����t`���/M��r�U<��=u���m��Cл�W ���{mQ�ܺ�J�B�U$��y�����%;�� ^��2mYƍ��y����#iZHCl�{k���t`b��0L[��đ�U���v�W��q���y�Dз�J76�\"�rN\Y0��v��w���W��G �	%�-y��֫h���YT|c����EWi���\)hA�!�0�6�L�k�I��I9:�	�U<A<Ƒ���S*��J$��}-�Ά3��$Ǥ!�{h�1_D;I���s�v*�RP�|:�:`2-��j�v:!�����3=��z�����[���F�#,��+5����ϛs�p5J���I��h.vV�|< �o�<ړ_�%�(T����/�?��F��HF�IE#ش38q�A�@��'\@ 3�Ek��w���",�]�=�w�р�fA���A3l7�'@����U�Yb9�Z��0Ȏ���R��p��;x��2Q�g�+�|�!�E6�h��e��K����B�:�D�%wK�H�tr�a�~E\���nF�?��](S�/l�z��^9h�m�M�&�ۀ$���
���m<��0�]���F,"�JL�������V�.��i����|0��e`��X������Jo��I�Û���
b"	�����r��_ʦh�ew��۴c#7����V��_#���<�;ݔ�����G�
�w�.��[S����vͦ)6�?�9��|=��b���C���(Bo=Qy��gQB.���C�lr?��dt��
H��T�@	6�5��4�ܜ�}\I�-����3'�!,��M.���[�.�l���U�o �Y��e��۩%���݄�=���wW�8zr���>RvZa�{
�)6̎�=��_(J�G<�^<���{ގAP�����m�l��>Oͻ%�Y�*����bV���̄�`ZN��6eќ.�gy��;>��}d�nR�V�3�5Cr��R[��Zg��&�e�\}u_[�ː2�-���7���g`�ET?�<Rx�)BY"g�;#c��#�ʸ|,}��Z&�$׉×2�y
qWyD
�@tS\��],���28z^W��ԗ����7E����?�+똵�Gb�O�ջ.�ã����I|�8����9r~ά?�Zp��QTe�_(� d�
7Ǯ�gB�SL;������b�-�<�L�n'����	��Lef��?�����c*�����lR���Ŭ9�Q��j[�����sU�{���~U��hd�cj���D{FA�-�HT+����L�iF�%��6X*�ifP�ҹ��#��?X:֭��]��L,�ecQ�e�;�x2�)+�7��ɚJTQ�ρ[��Q�\��(��h�K�7	y-�Va�5���#��آ
�����F�07"��C�%f^Jv��F�ҁ�){xRg#ٳ�(^�M���b?<��؟��?Lk˲��ߋM:�O���\��qD�X�z�ho�=1@����(DEX�qyp��k� ���֍pR� �F!�;���=�d��e^�U�I�|�d�59�mA�S��»�ܡ٭����n��+�f�_(�����7��ظ.L���_dq���Rb�i��i~C��Y|���o1E��!Vw�S��P��_������6�Z�w�_�L�:��@sYWH��*0�p1�'�[l�
�>`�|����}� �T|�/�܏�i8$S7�{�%`U�T�%n7���&�m-� :J%��F�a���6�r�IQa��(�h�	d�Pj��1.�U�SK�e��L��Ȑ�,�˿g-�y��]�d������|7r���T͚I��/�N�F���ҍ���������xU��S���+���֑���A�j��";;���fct�[��W����.a��y��Z���s�ݪ��=|���1"����t�\��@̺	�T�;@�|a��B"׆�TWm|�z&�B�Oe�s�ʵ%�����)�\��v��ũ+�����}�4�b DHAj�ڪ���\�0�#?u+q��[��h�~.ͬ��Ĝ��������/�$]�t�pn��/�ڲ+����q�vExkɲ��O7^��'���(��+.v2ҤwUx�2;�����c5���s+�8v�Aoa���ꤰ��3�ޓ\��R��mhԨ�])-��h��bωN&`�k:��5���Re�'&狨�d
n���}3��l�+�L�l��U�vB+�a�n�5�knЬ���̻g�����z}z���Q�F*G��6��q�b|���C	<FO�u n��,� �?����;��xva��@�� �2Sq@Hj!BzHG��?O��p�%���E���b��S^l0�y(���7�2�i/˗�J$F��w�ey<�H���K�i-���՚��p#�+,Ă��t�Jwku�O =!�֑��z�sD;� �	�^�JB�/ҷ	q:Y��	A<�kձW,0�C�Y��CG�<T����/�R!Ȑ_������Sf�~�l�5���5�	=���ڔ�n�mE�?n(��~��݈IC��y�i��`��sH�ĥ�ɥ��9�bb;Gf�#\X��-�3�*��M�e.�EEY�tQ
�!T'���[od^�ؗ��B�D�^e%iI�ޠE���&&�=}�� ŸÇ�F�ȇ���U؎�g��2��́���l�^9A#}�y�+i0�*j뢷�Y�h%�u�W�+�l�[���l&����m�>A~��͕���ؔd�)��x�N����	2��4��t �������
�q���P45S՜���.�K+X�m:)"� 7�0/��!�����V�Xy�	+�_^R�l�2+�}5r)bP��1k��������н5���X>�۷���8G��ey�$��"���4�S4�]�$M���S�:��a��W��	�U*r2�=8�1�`w���zc�E���־d�ьb�dP��8���LG�Ps�pS��^�Bo������r��J ������Rxf�b�m>=��� �a��~F�Goo*�0$��f4�hq��U�J���7~�,'�)C�l&���[�d��Ml�"�{^$O��9oeA�{����y�����`#��e~�D2�牙�jHq�=P�u�J�W���HP8/���@d��-zI1�vp���8/bO�*�;�:�`��(�"��]�DNB�/f�
PB�.�)4��V����B�K�Ɍ���!��X]M�4ß�
��x��,���*���*6m�{����8�W����qS|t�n�e�����P2�xd"�/�{�K�s�����D�,R��*��rdUP�u�'S�t$������Am�Ȏ��?��<� j��=UA\4n��$��J4ZR_Ŋ��Mm�[��Q��PCm����d��_`
�o��� ��������������J��rlznW8�+Y��,����YH�LxgLE,���u-�p��3}�{�.����v ��I�-�N�Ѐ1x�]�)�a�4�f&^��k��UY���2,�͇CJ,�R����\mDY�٥I>V%��� G�"X�P�A�E�I5�a�f)�K�$����_-^L���]�kB�����9�Xp�~3ƨ��sHR��oE;��e)H�� Gc����b+OLs�N?sg>�|EA&-���Zģ!��U��t7���ȕ1�6_=}�����֙FV��KW��<�5�aݠ��G� RRFy��F������*��u#�7Z�jo�k�����)��Z#K�
����=D�p�'����>�)D��E�B��uD���I��?=%�t���T�r��Yu-�������^ݤ�J�T=v�6Q�V�G��?�-5��jK��Pm�Dt��[[�D|�m���UJ@ct�<��j�q�=�+��7�s'��+x������{�����[���u�5���I�F��}��j�#׬૧���y�m_��h��ĽFf}�^�.<r		�1���aI�h�ƻ`Ƈ.��т����-�w��U��m�*fh��+#n���Rkq2�E���yHyH��-��$y�`�ZՋ-�ŋ�����Vl2��3}��lvP2�޶�g��=�y��8O�����a�_2+k�s�K�=��5(�ʼu�Q��8�i��DО?a^���v]⦗��>&�}�G�@�LW�)�7�njxQ���7�|m�Q|;���-�_��Q�7�<R�bi�QP���?}bl�����i��2UI���)�L�5-Dj#NC�O��.N�$�S���r^,�H�@�=Cu(�u��Wr�Zf/��㖺us�Hz��?�r���&�	|iW�m�� ���|���㲒���s�� *���/\s��2��� ���K 
�c�%@��o�����J#O�=��qF\�6��J�_��Y����y9n�ؾ��ҫ:k=�,�f�M��z$��]P_�mn�R,����{m��%�����^~uwM���e�oł~O���g��l�n�T�nĵ�b�K�Nŕ�j�S'��Y5��[W�G�mƨQ]z���R4������{�&�Ө��l�����/-�	O�1�����<SZ���j�3p������$K�ò�Yb��m�é���m�����"Q,�$�ñ�pԴe�a�@�Q��w����IZG�$62�������-}��3v���
���H��Ծ��K��\"�&{%L��W
J��K̜��dC�~�.�'�]�<��@������IdV���5�L�:+�W(�_���)q6��Jc����_vP�&�yt�u����GqR�I*P��&��D�6M?�
���0�z���`�6��t���T����>�t�r�� ��k��E��+d5�P���yuNS���)���!D\#�v���0>�w��y�?$�r�%�a������ճ�$Tx�ڃ'p|�Q�L���N�R�o꼛*�`�q(��#�@��!�(�-)��
����[+�Pij'������{R�[S�W�Y�������o�k���H���lZ�1��VTǔ�4N>z�e� ��D%�Ϧ9k.��VA�	@[�'t��=O���{D#d�eC�`�i��?�Rfì�ȮY���I�Wsa�ʶ&'^ﾐg���˴^��:�D�>���~?���,�Z0���Q�����T���cF�}$dE��.I��?�'Idk�~QR/gz�ߏPoe�|�M��BaĎ������I�\��t2%|��46� �wA>3���/
#�8m���o����%u��a�Mp��)#���i�I���?��Q&3FDC�2r��e?0�GE��b*�@���1��f�V�����b=W�����wu��ޏTV}��uU�ll�L"!l"$�q%��6YJY(���W���!�|� � bǫ��B�Tq7<@]G0O�#C���~�KG6����"U�d���aS�S<� �������6�ŝ�_�O��u�c%�L���Nը}����F��<�x�.�Y)��#A׻=�J��Y�e��,����b�ɮ�!�[��L^��9DÉ���h힦a3������t6"ZULG���=�O�b���mM\��8��?�I��1��	c$�l��y����`D�##V`��+���/v���&g�x�rO�׎�c���;d�N6@ط�/v�1e\
��NU�e��M�ԛA̬��g�oi�gʛ���e���`o��=�K��оP�$�x:#���%�o0�������ч�z�ߺ-��Y��:�ƹ�B��HSX�P�= /!�K��e�����9��z�߀�'٩�⡤��F}<|��e-ɤ����M��e a�&��r'��LAf�Z��Ј����=����������j������we�WY�v�o0"˓����å��$%�����o���r�������#�
U���{X�~�q }Tq-d�[���vڳ�3w6G]m��tpd�Jl�:]���s�dD�g�B~hM>�u%�k���ջ.�\;�W_�K�Sb�
�9#'^��\@z�W08%�r8�Zɶv-'A^p��7N�*J¡���]�x��<[E=ɯ{2��u��R�:�bX�v��,�	����֯����k$�|���K�=�����	`Q�EB4�/GЗ�������{���զe�4!����:O��WlV�I +�f@���,�r*��߶`��F�,m������m��5r�#B�ap��5/뫁�`�����90��nH��_�ܙ�σFI������t'�R	_���bk��0��rv�
��l"����Ř�<�^[8��i��G6�><�u��x��� ��сX��d�vO�M&��|{�B����|;�w%�ty[��	��@H�nG�[&��`h���s��"����J��y��9^���n���v9N�a�*����z��+�v�#��S�Ĕ1���k���x�kP�@�"Sew�s�1o`-�p�c���fԝrG�H�R��)�ԓ����q&����W�~�D)>�5\h�ef�Za�S�g$)�U�_��F g�A�i.nOW�����	�̡��dD>�7^�YLD�`� D`��v�����\PN��"���U���S�K�����G��'�lGX[�1J���mF�~�@�̵��y����<�.dԍ����P�l����)���',{ ɇ/�c�=�����8����7�c�.ѣq���� 6�s_�
Q4��*s�aY��Dj[1�r^-�0��wj,�=�+b�DF�)̶(ˆ��7h�ɴ�垑�J��B���9#�>S�!v�ɲ�ߔh����R�|C�F?����z7,�T��."�j{���.��ڂ6ܳx���p7dvハ�`@�x��E/ �%Q]f����쳶	�@"0<B�X�5���M��c��Dy����{x~���:�4�[���k%JȎ�rxr{�N�B�����o�@~LjcⲞehww\j�U"�2a��c�5�L����5�����r�kZ2,�A���B����(����n'Ww!|HD��X�J�� ]=!g�h?C̻�U�� �nQ?���W[vQ8�����ݻ{wh�N��4[� ��E�Q8LN�mO�F��6�|����Qy��W��i��f'K�ڂ(������֫���H��״��+zl�e7�(ׄ�׻�c�f��Ⱥ��~�'?C��(ߕ�W��Q
�Au��ƴ|�sm'F����QG�?̾׺�,Ս�GP�ɔ<�����I�ĹLE�^����MY��UpG, J���(��\~�����ϴ���3]P�e$G7j����ҭ�����)��K��z�@�M���U�܄��ђ�\}/|G��7�w�uNT��o%�S��b�"�$�&[�0G��݉�D����,T��1��E[?+c�A�岡�=FaE-��t�M��b�2�P��P2~d����R�Š��Ʀ�O��P��I��+���X�����l�T�55Y$�A�طn	���5]��n�ԡ��̆�W	�lD������]%��%�@hMq�J�f��,7ٌ�?��:&���c!���N�U$���O�~������0>�b���ʭ�^�M2�&q�g0���2\<�UϚ����q����j�p�Ln�nt\�jS�%0Qg�\��ԡ'�مS��GA%�:�޻��P�C������ DX��R6yŔ\łiD\]�/Y�o}�f�h��5".�Z�,`�v������1�&T������U6d�M�{���o#�C}P��Uq�����U�F|㪜#�Z��N����Ze�@8��!�y���1��,.�k�O���ʉ1�@	#�¬���R�\�8��/�f�����Z������繐���&c���'@8B"c_4n׵z(l,T}�.���0��n�Z$��A��CO�¹ՃPM�����R��U��ܻ�5C��D��Ғ�A�{.M���Jޫ��l�����x\ஐpr�)/��s Ywث�������mBM�5�Ē�n���g�J0,�ngM� FHVd:^nq�40��t�㕡�6�MX=��=�-gd���j��Qq��;/�2�w�%C�:�^y�t�=�eKo��gǶrh�'^g�(Q����L�����@��폀Yf������R]�<U�v!*79n��鱴Z'Ѡ�E�>��cSi�;#�]>���H���:n�KP�ys���6;�]��w�ܟ�njvth�/�:�'V�0��wgR���(��<�g�Tr'ѣF0� �_GE6�P�Y���-1��.Po�}���X ��b1����u߅��,$↰�aT��Xl�A�߽�NI2�Y秒�ף5f�փ�-��L�1��.���À0w,樠���!8J��J����$���Dg3��b�#mGcD�����%B��I��	}��	�h�^��4�v����W,�ч�k�8���K�����e�
|� "�b���+��7�-I�P������+	��bf�
@(�:c��M����{�*��v8�����)����2���|�^nn���r��!���%�M�l��pڬ��қ������2����H�j���4?J������oL(p���3��	T��$��R���Q��V�qOi��<����w��V�>���NT�R�����7v^!�Z|ovNۥD���T�1�g�6��2�	�
�d��gZ4SHP���ֹih��Z/�잋*֚@e�6y?�sQH!�|��O�;wr]B�h���� $��Yκ�L��f��i���+5��Yk5�v�I�`�ʑs]��Bo�YT49I��D��K�w�*�ϣ���r}�Q�^���c�g\l{�;�A��:;��/�qH��I%�$}�*7p��#�1-,ÿU�19�}�듬��oD��G-�sT;�[�&����I:����#��� ���z����`�m�H�x���%ܫ%�L]�"�#Ff�D��\z�c�m�V6h7��֫+*�}�MF��e#�zhlqJ�
{���n>�'2�����<�W��S���'��CG{k6�Jej�!�˂�4����q����&j��6�.�v���_ø3��~���B�O� �sb�{��W&��{U�r��~3u*���w�C_�0>��T��u�[F��$]��V�
-���y7��ay�b����ײW7b�E����|g���ٌjB0hHb��B��k�?�� M|*�;�,�0>L�9����y�,	];!]�p@�������S��v��9�"����c��|��A��O��7k_�λ?n�fZl��0�I��A�pZ4,�̴x3x|���:�y4�����q�m��d_F�p���c	�i��M��pӪg�����8~�˛8f��:w�^�d	�#�a+XVY5�넶Z�������mR�{|���d�� 6��T�����<d��.::b��n�6�s�YAx���j�fX�U�qBnI.�<��L��������˥��3���u^�+By�:u�Y�����E�:cCE����P��'}J�w��\2��f����@�e�N��n^�6'Sqdw��w���t.�n�d3��
����$���v�������X��{F�N��C���y"���9'�=��o�}��ͦ��(J�vz䊪�p�2����G�7J���J�E����E���q�Ȳ���������)Y���e� NĤ5$3�Hɮ-3�!)V�8�����*G�
�xp�<G���Ye}���F��l;+��"H,~=/�)��t~D��Z���C:��M�<��m�"�5ҳD/��'<D�Ն���d�0.=��n��6�8���k��~S<eY�_��� �`�{07�{�b����s�hW�=�\�3r\~4$��s�'����|~y�����!�z�w����n
��%}�����t����LB��~�%�U�[�%�L�z(�����~�4[��H���H��?J�[V�,�5�M7A�'����fĊ3}�E�N�T����9oFM�ݎY�U�=��W\8*a���IV�7��rY�o��|z�G��1ƣVt���]/\/�S@p=2Gs��ETN�\dT�폛o��!
Z6!ۍ�aZ<oX�K������^���b���?�(��u��,*��m�
���͊}�
�k���i
��C5�=I�?o�S�#4�Q.C{�U���]Ӹ@�̇8|��y��[l���H��>I0^�"��j�B��|��rJ+ߎv�"��g�?)c����;j���\7�����W���rf�������Og�_��pr$�y�V�{��8+�e��7/I-���5���v��1gEY�v�2�+-&��@/�Y�����1�,���Yo+����7�,G����ga#�@*	�Pf!�Bϒ��?`��ʷ�3���n~���"�2�9��4I���U����V�v�[2�f�O��Y����)�xP�5����VT��!��C�"�񿂛}K�;�M�����9�2��r�!o@nB��vm4��-��U�SQ��ڍ�I#����3�.̜��q�O�V\:Z#V��\�Zj(À��b`�MGnСN�!_GƸ� A>�<�t�Md��^�	�u@�}6�^d�waL������.�V��&��6�����Ԡ'��I�+w�@�,:�p���a�V�n@�l�C�?o�!�1��a�&�_�
׷v�ω������M��B =��1d��,ˑ`�6V����]q�� �a@�T��szv�Q�V�h6��p�����q|��r�W+��H|�O��F!A�l�,�"��̆�V�$q^�ԏ�cR7�� Q�XE��+?����M7X����X ��4r��[���@�e������������`	�#�Y��*o("R̈́���8O&m)o��'+��;��KS�����	���v��ITv�Ԯv��5����a��l��>���q��p~D�R��Iĕ� #+;$�1 �űTb��oD՟%�꺙l_���[��yO��ٙ[N����p���"#�	>���lMn�@���wn�ѣ����� �V۸��҇�?w�J23�k#`�н~�"|9囯
*42լF�*����~6�)&�����j�Qz�O�B���e��E�b^��ж&�썍����z�!��_R����;g~���C'��&��I!�/ox�L���?d�O��!_�I����E	����r��:�К&���Ɯ�m��*_O���1j��E�cρ.���1��v�p$��z(&yCt�@�!��m-��{D���N�6�!��`_"�l ��f��&������ʰ;�/�M��rF�W_UQ���V���A��Tq���jt8Ǯ:���4Y!s��U;�������	��/_薻����^:1Y�dQw]~�D���&��K��<P�/�$:~�<|p�1�f1�%謁%cbe�eWd5^�� ���v�D�y�k��ݎFZ}�
���^^r#�6Ӕ��~��u�B�G�Ί��)����,�0���R��"2�=��o<���0�Y�������Z2W$�T� KHMAuW>&�X��"��_S.hN�289�qd��c�PȠ�Qk�@��Bߧ4(>�y5'1^��x�Vgy��X�%84�n�'�Q��E�����������<&�ak�ITҰ��s�Ͳ:_�.�LD�\���0�ZS���5��'Ie7�F^
�5��0�	���&�\|,6��x�3�$I��htO�:���[=񽝜����j��ë A��?�}����2['tP��M�IT�Wo����T�����4:�������CϘ_�uݥ���1���C��ur��ΆAG���u"����Y���x0pu�3�`�"b&�g�s��Еh/s��#M��A�k�u��<��iV�蒃e�� 4���y�ȬR�L'a��e�p��߭��f��\�@��e�G_�Phpֲf���w��{x�[Vmh=��V���s�lF]m*hP6���cWC��de��o8�Hq�j+y�]ǀ6t*�);�y=n[�k�5�B��B~���ؕ���V��^��4�(�*M�2z��٤9%�+�.�;kzA���B����f��c�;�V���e�l�Y�韗�Y����A����j�KE��y<8��q��_l^��x��~��;��=	'-Y�_�Y���q�Gs.v����zA�>c��o(��ߩ�����NX̝˓���k(7�&9
b�
���(��ӣ��9�!�A��B_�z�s�?�H ��lsr<����9�[AT�<̖��R[�@����]�y(&���|�<��5����곯j�"+����8�{%�s$q�k�6��Ym�Fه�%2lwIW��	�!A�����f�c(�I�=�a�$ g��K��iSQ�	�~d�a���G��r\�(��M/3՛`��;��#�7�g�L�rk��RP��ad���f^��Q�tQ%D������z�?#\-��3�2Kܻ�T�[h� �Kᴽr0��h�(�I܀z��{P��iS� ��c�V����ö3�a�}� �:�ڡq��]�^G-*V?���!���&i-x����G)P)�I�μ�w�N����#�v�=�i�0�N8�i�������j��-�F��퉦���o]��O�<�2�$�HeQ�ڽ�0-����sӅREw�#.�f��ӄ�2���O�C�H/�*���Uq[��^I��M��5�Z�do�ϰY�)/���*�R�4�H��5A��6b$�5P*7��3�QX�&O��.[��#���X��=���W���˝�}�w���\_/i�����W�0��������j�>*��:��X�+�m(oGkʾx�D�\���xٗT?9y���S3����
MV��Z��b��f��V�J�g�U�p����{V���l���c���*^��m���;�x�t�5���3�O`�7�|0�nߩMo��y�G� `Ol�	I�_���[��5�5�%�����v�z� _^�P�ʆ�\i����hqnge��ZZ�}�j�0:`��}o��IPV��&R�I*	�0�9F���i�q<*�j�׽_fF��T&�b��@ɍȰ�<�#���b�3���q�=�Q����}�,\��@��X=�����d�o���[�����t�)w�	5z���ˎ�F����pՅ�_��P�9�5�pZ�R���jO��E؛��Ӛǘ�D��n����N��	�h%�i���v��<*�PX!Ov��$���a�6��Ǉ��V��{qV��!i�ʖ~N.�g�=�BT���)?���K�ڤڤ�i�<�bO;������_ʹ��I�2�Jɛ�����C*���ɓnP=$6w�����,#Qk������Q�t˒H��z�day���{h����m'jck~ ���%��tci-,�¤�96j�B����|8I�=�x���[���#U����\���3��-l���t-5�-�A ���0\V�,1RΧr>�]5_�!a�|b��R�d�i呮�Rr�%�@6��� a��,h2���`
!�H�L��h�q���D>n��t��A��w�&���:�a2������uy:�����m5�8vciԟ��D�$�Y�f��vO�	�S%`��5�� ��|`�f���1Ɵ
���tK{����-���G�[2�4�������2��Ks>�R!�;���Yli�gc�wŌ�Os�y�"-�3�$�DKs�9	����~���-L�r�H�VZ�L��d�(j���<��V���9,<��N��Ϗd^MC�> ����Z�0�2Z�i�ss[����r�-����*���"k�43ed��	��b��B�Ig����4�ݘ`7���1pޏ�Պ�x9T�9�w�:��;��=}�u�l���b����?��������#n*�/h1�J�v�	c�ֲxj���򃘃=z�|���Zپɠ�e#��\�E����ތ�h� )�!9�z�L_�*Agh��]�dM�ʱ{u��h�nnkXѳ��;ի�+���n�n���E�ƶ<胿'����o�)`���
��|�Ӎ�r�C�����4�D��D��r�!p#�%�o�T��d���:R��FI+�ݝ Go����]5�����%�Ɍq�����)�`�Wq�u�Z�pہ��5��7��j�����������(o�D��;�TTގ*�
�'�5�SE �������2��p���jD��J����-��?%0#���*��5����B�K�h���^��i�\�������7�)�cDıD:4X�tyJ������Π����U�ew�G菓��v�������k��H嫭�A��U�r�D�t�ģ��/19�r�����Ǳ�W��4�"���ԽgNǑ�X͠��J��a�ɪ(�L=�Ğ>$�R�[f?�N�nX��!�5X�H:�^�ג���ǖ	J8�1C��˚wj��;�- ��@'���q�����N��F�95f�Ph������i��h&��1���n{'������M8�y[)K�:�l���f|�����-�D�,ZM�>��D�h'feΆ1;C�����TH�Jjk;d��G��ݪ��k�pW�z��k���p�~�bFNDe���Üt��:5n�F�D��,�Πd
o��\��v��^jay�|���wD�k�?TC88>���P�O��	oVL���� ��[�����aF�#�A �(��#��A��1���K�,��~y�_!��Έ2b���k�V�R�E_��L@�����)غ�#���+e`�@E�+H�Oq9�p6scR5j��,�K��b��C)���?�eN�$�ރ8kcOv��-�c�A�0�.nŐ �254li˔�E#uo�@�bc1w٬|�ԓ�A�A��:e|�h�W⽻l_/'^���������� �
�K���d��ފ�扊�e����TI��\��4G�Mj6Q��tx��u�V-&��hk��#Xr+���V!8/4��H���§�����|����i":�:���H�:!���'�F)|<�3O��`F)�8AԘ��:k��]���/��&!6p�ÝIH��m�������ob�&�ض����d~M��T9�x����A�P�a�2|�s�kg.&��+N$� K_�0/	�"h��m�66h/
�w�e��L$�ڃ�Z���'�-�h0D�4w��Y�<�!N��L��X���Kv�>�K��rA#��Ӿ
?*����r���D���I��p�Txn(&��˾�d��4�S��4��
�<p10�1˥|�)����7e/:>F���f8X�J;�ky]Bߠ��q��"���-�w�gM~���/�B������(������@�˔Mt3[��Q�1��$���Gp�{}{���z)œA�Cߣ�� �2[�G��O�<��Q(NzF3�/�'�3TE�9q����@ �]�{��3uY!w`j���b�&p�6.gZ9��=�V�����T�� ]�?�Dnj4��������Q�&�����{:G�p�vi� �3+�S�����O&��h���Qi>4; $��t⇷��ґd ��Y���F���{\�ˉ�;�=�)?4�`�*@�O�����cAZAɝ@�4@�� �4%����X���Ѿè�)���aW�)����Hi�����59��u�4����GDSb��^0���.���W��)g��nZ���_�6ّ_|A�==q�8�T��6����K�F����t�k���K|�]���ۢ~w�gހ�]��im�Z�C���IQ��ҵ�ԅ�K�����(�T�P�[��	D��S��
nX��ߺ��X� ��X#͸�e�=>E�z^]Jh�j�9��b���67�F�������7S��;J9��еzwR�M"�͓̙���� J�W���L���D;�z�L֣�R�Q����q���D�b���]!m`]����C��!GPt�a9�Tͣ{�?$�w�~]�u	#���oDΩ����]�d��AiZv�2�M�X�v[��:���p#C����m�Z�+�؄q�^�=˔Z��4���'"D�����0�o����{"'������1{��t��������o(2���ŵ�G2Ń�BM*�Đ{ai�!��1��R�,DZ!g���.E��5�:�«��0���g��n����;���P�h
Eݒ���B�̕r�	RhD�����;���O��%ڿ%; W��tE�u+�-��a4q.�	�W��,�58���Mz2h��'�a��7�o4�g'�T��>�G~@��I3��I��;E�]@,�@sje���kc���Xa�������dߏ�:�ˣ��F��h�!��v��Tv�2�$� �:t,��[�1�y��p�6��Ms��Q�L3��O囼"{�v�C�-�uݬ���Jn�K�����ݥߴVox{���!����w�u��❝�&k��IZ��3 `b�� ���(��km*��Q�7�@�MS7����=�"Ԗ��!0�k^S��z71+D�ހ��Y���Y�?�?��J�H���0�y�M�뀱���!-�S�����R!^�����ӕ+��]x���PYI�⁮��hJ�>��.Y� ~��@,�I�۩}ͱ`��~z0k��R-y|9�!���
�6��ʏ9�k��R.S3���қFn�O��/��N+Z��q����;y��2���>_j�g��^��1)�>���/��󠂍�'��+B:��~ʏZ��.�}$�>��ȉ��� <�{:7�m �\m���:��2�c�.D�	�4�a�M�CWd���.� Ub_��Jq+�gl�T���/������/-�ܚi��-З /CB��%�mx��6_Ԣ�d��Ys��}8XT��n�T���V��(]Wŕ��˚�WwWA���!I%���n�T���Q&|�c�w̯m��)"��U�+	GX����7~F�����T�Ol�Uԉ�&�0@V�M�fЗ�uzk��l\�������|7b��9��z�F�~��{Fx���XC��b�b�8�m���M�nN�j^�_wK\�kt�j�zO=`�f4G?U���:H�3���Q��7R��������	3��塨b\j��B��N���"��t(�5kex��<l�+��9[��,�����ѧe����E��*u�/³y�2�ҍ�����z�h5�(�a��V�L��دẞi\�#�/���}�n2��������!8�!l�E����P���j���p3H�޿#\Ġ^���B	�HGl��8��*�*�O~\���.����������`&����bH��m�.!��M���"*�r���n>�3g� r�w�=�ǩIv����\]�>B�-fPA��6���O//�?m+ւJa�)Zw7%��#H��{kK�y4�,6���5���a�������
!��+�	��"(�6���TƑ� p%�*����/�m_���@t$"�S����������֖Q�Ű�:�Y`�G�:���.��賀p@J2���2���X뵧֟��Zk"���X��Ay�"MV |�M�z�����	�#S"=��EcC
3��1)�K��K?��� Mߥbc��0�$�� L��9���|AW�HLEr�l�d��Ѫ�
id��
b�U_�B�Q���nƾ���Z��>Ёj	�~)ꌞ��� DA�y"٘�[�{�fPe˖rB%��/�Z��������w�|7qu{Ξ�)�CXws�r?�`ؤa=Yf���`m[�n2V��v ��G���SJ�����(GF
(4� y}V��9��J�I��QԲ�v����;0{i]oZQ1�o8^aY����2y�vlCpJ��{Hz��_��<S`}�R�{G!��xT���e�X�>�U
b;Ӏ4�S���I���Ќժʹx������Wr�OQ�<W�B=(%40f���z�~F�c��$3*�[��	�ͅ�E�0��鉁��V��P[�v\�%�u��v�Drmr�d�\�\���v�9~��_of��{��Q��×����(�!j�w�}_�u������� >��.ր��G^�DD�rR��EÙȆb�1���=i��M��n�2F���7��K�_�������R�`�\с� �c�Iql��ie��I��-�~�2y�1w�őh/���P��q�`���%�(T�Igo��!U�𦺵kq��������Y_�@SnbI�Z3��E�Gw���;����:��<�����8D��b'����"j�xV�	�f���@�P5���������a�� :��H�] �̈�fHз�������Qz�c�:�A�^��
�^>`�m������t�V�?`
�S�oڞ�H�m�9�k����sà���E8��LK�ʷL���y��<�k�Q\�z/Tu���A���&��.�~Vy���@�#�ЙOd��r�%R�Ľ�j�(OCo�rPa���f����g��]���.}�=��_�3	#ԍ�K�ډ%Y�!��y=��d	�5�Q�WK�0^hzD
Y����B@laĘ�T�φʔє<X�\o=#��,DG�P��_"��
�{�͊Y�I����"����y{}�뚆S��O,��m����Z�!�ϋcܠB�+ WpVC����:f�����a��>$� C�qw"��P�����W$z�N�m�17�RM0��g����1��R�*�v�u�I�"�9��G��˃ƻpۓO�a�� ��+��_�-�1�-�V���!o�~U����7�ѸH6�cմR�t�^�+Wd.�7��5ŧc�t�A{c)���fF����#:b��0��u�J��q��P��6����S���2���h}h��_bY�2�,s�<��p�ha�gp���M�R��P��$nI�2!���i@�m#)\4N�{���L���u������9B?%NK��w���o��i�	�����G�JW�T��b�3���o�?�%gm�8
�g�VZ�����l�R�Jpb�,���-�K�=81)d}5���=�Z�|$Fb��f�./�xj��o���O>��a���!���ƴB�Kw�9O`"����r�����2]�3z�2�ˣĴ�ߢb���c��H��f��� ����%�`[t<!ad${iDcH��/���%�N�B=�m$��9Ƈ��=��%��[��$7���������߆�SJt�}��x�&����$@����<��#9��c"ۘ+6��hƙ�*���da
�wK�/.��Ph��㫊r�?�o���"�=
u���PQ���b�AR�������䎶;ª;��J�e�G�(����8��Z�&~����ƚ���8K*+=�mVA0�^�8��4q@O7QAb��`��V�C�J�Ʉ�Њo4�Y��z�7 :���3T
8G�Hőv�08>��L��y}�7*�	�d�?�����$�� ��HC��%Za�(	��le0H<H���b�ZL"El0�?v��@)x�[�u�S�z�!_�v���z~���}��2ܽ�6T뱢�J��`��*g�?d����8ǵT�=s� �Q0u딃��co���)�+��@�s�I��#.p<8��R6=L�ty��Aa�E�����p<4@�C�G�n	�?��̽9#���1�bD��ݖ�}٥:�=(�l���X�R5=�V�w�����F��A�
�x��~^�X����*y߀��\���?q`�g]XӗxO�E�l@�Yh0Hv3v�	ԙ�H�P�7�q�25_�f��X��'�Q�Sz�Q���? E����Â���q�I�;'g�Dy�C���E�] }w����m����
�*5x�v-����̴�5�#f.��r�jI�ܱ1����V
e!�Q���D�C��r�į3u|�ض��p��Z�[������B!�<H���Օ5PO=%�=~���1��׶�+�y�:HY^�h]��e��լt��骍��L��H�`���8��viɸ� �r�e�1��A���9� 9 �yY�bT�"7#���f-��yq�f�<�D�0��gs�j����EV�X
^�!���ɖ]E�� r���u��@\Jle��?	V���Tv�lP%N>t�C�������rHSK����
��L�7�^L�rl� ��2C�b�q�P�].�"����[W��q�����G��5I�x��)Eב�=1����j�y�{A�Hvi"��P�����83���߇����n欎Ե�V�m.�)�%࿪K�, �$X���z�<*�R"l2�`M>�v�l%����|�)ƛiU��4�t�R��5/��&i�B��ȉ��\|��$؏ "��o��s��1C�퓩5��_{IL W��ԗ�Pp%;�a�43�_z�ɳ���:�w�����l�#�V�\՟����ƃ�j&�������%��@����Q�E��6�N ��(捧�͹ ĭ<�i�#�d����~Ҥ.�~ԇ�
;C�'���d�د)�����Px����o2�i6լr��_u�'1�4:�U�T�gK���7��6�y�ֵ�z�����ʋ���BI�U�������H�V��&ٴb-�	���������PlSi�L���O�������#��
�,�n\�t�1��0mt�Y�j�I9�T~��ZW9�7G�0�ǉ)�j��Gޮv������j�#����J���I�7�&�H�!N���O�Yj9ps/a���}�7Ț�iwc�>!��r�ō� ��x�w���I�"heN(y(hm;����sJ+��!&j��q��]�b!�ک��s���@�[i�IH~ڕ%��! ��/�K3�\m�����K�g*|��v�<@-���G/X���b����+���y�|+�u�*
}�b����"�>k�?9��)���2�|�f�(���>�JZ�^X%��Jへ�m�	%)/��Ƭ����J�ۥԁū�-b��O�:�� �[9��^b�N�y�:��ȯi�^�*v7�M_���.�������.oEL�	������Q�@f�_�ܺvtW�G�f��E���F������ȇ͡c&Z8J�>,�v//�C|��T�7S��P��I8ȾH�|��Fϛ�W3�y����D*���N�&ϒ�|.���iT���_��� o�� ʻ��}�s�'Sپ��2�$U�ps�����b�}��^U�Q�Xw@��ѵS�l��!�Rߨ�C���,v �9vl$宾���s��۷|I� ��3��В�>y��2�i�g�ȧ��x�q{�s�������N/�[.h����'I��bŻ�"5��\lM�G���ӡd����榮�ɞ�14p�ԩ�Z_14�� �㵫Z�3�%k��D�\w�ݓ5D.�A��V!sxB�ClrV�l�4�u7��Sn��T��ǯ�8ӷG�z@n�R�F�?���,M���7QY�%�`�f8�˰*cKl�(�l�)���ԙk�3O�Q�{��v+R��!�n~�ߙq����/��j&�%��o�]�p�:�h�И�����H�#�=ub(*�`I��_��/�~�(Q�-��WqH{Pa�
hu<�ce:���P�i�^��KvUU>do�A�=	�@�O��S@��_ƆDg�a�B��U����$������#�6ʩ�h�j����,��T�s��X�V+�[�H������[_p�y"�G��DyC�}N��5$%��ȑõruѢ8l�:�0��:dǨXS&� Ke��v�ZÏ�D_��]�;�~4�S̀s&��R�$xE�ځ(82~��bJ�o��N����������"7!O@#\v�utЂ�[��O�t��P�<�ً� ���R�5�� �͸��lMH�P�H���b^%S��;��o�H�v�M��O/"�V�4�>�L�E1����P=·Ƹ���w@L3��Dʘ��D�*�����X�y��/�4ja�ik��;�T �-��Ňր�'�Ѐ�����:	0�k�ɿ�0/��5f���ܞ��`��^+(C��"šHڤ����� `�-��OO�͇��V4�X��CE��Z��,�����2T8�!��i�G�9��-б�x�8X���`t*�׶h߉6�4W�ӳj4�X�Wߣ���x�2�{
����Ŏe˹�S�Tݘ7bP����I����3�M�醐��g�b��9���Z�y:_��=5%�L1��+��0)�*��i��
��)5��z�]N�i�JA� ��z�F7��Q�-3����T��B|4��=�r]�r�i��" -���y���"[��T��u�����Cc��¯us�[rl�>�Z��d�zA����� �@$`5/¹ޗ5�h��Q��� �D*)��Q���V�3��8�g�0��{cXU�Q����_JX�Z��_�vv>��/6�"����.��_�^oL��J�\v� �4$�Gt�̟��+g��["S�Ŀ\QY�Wq��j����x�B)�O�E�8V�|�:<y%*�2Lx1����gk����啬�O�9�)��x�?�Vb�T�ǬS�������bP/؄���ȼQ�Z��i>Z>NL9:9��	����j+�B� � *�)J�3r�L�uǸ�� [���i�Դ�:�k�8��goW`�\m��%f�E~���{���,L�/�덫�6���sn��xrx�����b �id�Ü�'�ͫ�k�x?g	[H# �]e�&|�#���	�[O����7a�\�Ԡg:��^Z���gK`c|���zga�׍���ru4*�w&���E����>x�2��U��pF�-����H� �`Z�-/-?B��8tQ�+U2ˈH�|쎳���t�T�f���܇��(˱�U�����3Ǉ�5]"x��2�����sЦtL�P�6w�[��N6�]��g_��4m���B�z�H�5}�ϡ��h��M�� ۬�yg����*ѧR�jtȽ_J)�3
o�oM5hZ�����_L]go�e�Y��b*�?0n�Rlb*?�+���S�@;�e�L����ݔ�h���{&s��>���I�t�54�הyݍ3���m�^�f����m�P�t��:(�8{�9:�v7�m�c�(�h�v���G�7�/K��\_�b�Lމ�� 0�kӀ]�R�H�f,�\=?:m�-8�ݒx��U$͎���E)��];��4T��B����]�"}PesSD�Y"*�h���7��<��]�`$[)�^mr1h9<7XW��\��	��v�Ow
���4y����hmI�8�,���Lg�]e��\�}n	�v����l�M|��>oK7�:��t��t��UB��g[�`Gy⾙d�y0�H�yd@j�o���Zܮ �Z��?�-�S+����d��$+��	����bGۘ�e�k��b��8x�ٗ�x�ܷ�]�!(� Ӈ�GF�A��ץ3�Y%[?&�X�M��{����� B�Di��iu���='��XE!L�W'o7̡P	|�� �~L��誦���/80����Awiy���������kVz�?q�.�|M~ ��8�ε-��˻9v�~�ވ�Z���\�a����"_j�򯓀CO�,^:�����њFAL'�Z�Ѿ��_ژ��Vi��++�ŏW�B���j�Q��+PS~�Iw�qm�|�.G���2%��@;ŭ����d�:V��SNlw�m]|��<Q�jO*e��u4!AK'���紣�-���0�N�r��	n�-!�/�c~\c�7�C|���$I�0q�m��'��B�#R� �c�������o=��I����;` xZ��t��'�O�Z���S��R\����l��r3i��f�#�-GQ��%�`���;�2�0 `�jF*ΛU��d����3~���~�~~���ɧ�(�m�z��;H~\:^\"�,����Rǽ���ۀ�Dw�]���� ���Ue3�l�n��^>@����5\���2ZD��w�q��!+ΒL����)�c�$�?����jZ�T�O�m/���A9G��ßgA��X̀��ϧ���-�?�w�R���P�h�Ȑ�G���_܀���,]�_n�� @�!(�������6���� � Vɥ��P�T�j�����#��^�g1\��F��F^�0qR�K�\����o�TuQ!�^ݼ��	��x��Y1���h��b7旰�����D���?��S��m�p�)�g���)Y��<q�P�u:���o���bM�va�?A3�å��S]M?��j���iY�:�Y����/�J!�߬�Y�(�Z���ɇ1w��t6S�bWw�*���a�s| �dF��ǅ�	��o,�TH��y�E��� �$.T������8���H�����j�	2`��*=�B��+�Woj���f][�M����+Ir�ʏAG��8�Q;/�^���.	G��Z /�^�����d>�C}~�{`!��E~����*�`"fS�و�["I��1�ܷX�b��-��,2�K(t��.�~I�e�Ɓ`0�ǥ'1�h�Y��K�ym���i������O�����$A ���ًM�w;� ���?JJ�R��E����m���NdFG��Q��wI����~x�P��h���M��Y�:�����C1pɵ
�(�ԡ��Y��]R�� �2j�)�0��{(�ݘ�;]���O�߽�^��7��v泝�z��։��]+&����s�"H�}��<~�"r�����ٹ�J��&�MT�0��	0�Qwå��s�l��$ύo�v���c�ΰ���SRxb�R(�
<nᲹP�`�x'����r5"^�k��_�I�KlJ��^Oo�����~[F�_���Z����
h���fɒ�|j���� ь�����WC���+���yٖ'��#�����@o~�:y�����k�%�d(u��A�t]��I�f�Y�W$�N�D�x�ߥ|QI:��Z�3��>w�ly�)|���8Ro���Z�m��^���ä��<��{z y���>x����4���R�3���8�^�o���P&b��բ�MTeG�̸��3�J�[[w _��j�W�5���%�q��p��x�,�,#��$#Fs�r�N|�_fq�$e�Ej��KK[2�ڈ�R�EDl���
��_�����>dtI����3P6T��H�{�pe�^��"��W0�_�`	8w�v���F2]�;�( p�۵/\��$y���6*�����l��"���=G#�Qu"װ��*���N)��ϘT�Ņz�ր���0�ֲ"����[Y���#u+�)s�()ؾ=\6,��$Cǭ�#�]Ԉ�3��:�Р�k�'g��5�16�O��t��	4^��6��1Ɗ�5 1�P��=�r�N|��ʊ)|�P���4_G�^��n�gQi���$��d���䬯mv�$�������P�u/�}�IA��_�f����|�A�v��o���jr��Z~h;Of!E;�I�	�7�_�B�KI6�YTKaN�;.��=<�1�C?Fe8��B���FO�įg)p�_��]��n}c���p��#�U΋ %cs4��Z�n� _���ś�1��p��"ȸ4^�#��G�9�'QKҤHFY�4뷌1���|nF���\�79D����1іx¶I�qyG���0.OGP��PJ�Შ�x�LQ�~I��{��?��O:�Te12�����Oa�Of_�\�g_��Ȳ�C��OV�-
=�|e�Z̰���4�������L[�*�`3�͜���/J�d��99�1�ի��%�H������p��Ro�B������O���i�;��v�?�[��ǵ�<j���-�ED�$d���`(_�<ٲ�R
@�cc{M}��kj^0n��wG��G�e�^�T��y ���8,�.�6�o�=Nz�s�Ԓ)L:��^~���4����煣qV)���)Ɲ^�U��Pe$����=�"m6[�IBE�
P!ڠ\�S�^_y�7ț�d�{q���<����}�m�h㇫y1c��X*�0#XϾ����%d~���l��u/)-��?���K^�~��B\�ԏ<�Ójp�+kfv�R�uv�>pYs{P3�#!f����;�xE�Z���F}թ�T�J9,��Du2.Q]br����}N��L�H��"�����^N��PLei���O��$bi)׫����+�:��-oM�֤����� �>�<�ח�ʡi
eʱ��c���l74�������%�dW��y1|?����z����r~�չ2�Xi�����mY\�-��(Z�h"�� Ky_�ȩø|����K`l�������8D'��|�����%�z��.PV#�=�?�:�(��Xy��L�:[��r�鲮�.S����/�#�����m��w�7� ��.��>o�g:��	��.��0�(������Y&�����+��D�V���vZ'��7c~0�st�RW��;t��?�+ R:!yڴ�@1�;��Gs�s�$B$uW.D�8�Z/~�B��W�x{xhpk�>��/�$�D��H��A�%��N:���Y^2��-��(}�9��W��_}���ֻ���xЯ�����a�)�o�&�Jy�dwKY����Ns��wϾK�Kui)��
JF��7e������XH�
�e��o���%%���%y���%D\��P���д6�]E�
8!��N�
�w@�R<��,XF<��K�4������]�W:��
5* ��|y$�{)�'��x�EE ��fJ���r)s�=gJ�H��2@m�%��8���k!�.�mU	H��<�����IdE��rC�.U8��Qv�݁�$��R��QL�B�ّ���C+�����5��`�5o���T��V��9���l᯦G6RM���m
��l%���ж��Q�#��e���温MBϔ�!}�[��^�����6���i�5��>!3d0m���-3iIC�!�P��bg��$�xh���� L���:n9���O����w�=3R~�L͐~�LA��^�Ӂ�Zē0U�g��Rn�H�a��C�������OFTJ9��Fn�����K� Ns��=]ɲӟ�,0D���qP[[���4Q'f[���k�	��R� �)���Y���o�������
+�+ތ��|���I���%Q���BC���pV� ������eّ�%H���p�8e��JÒ�����o�qކ-Jvʜ�Iv�T�7�m���3Pu�m푭M5%�ZO#�h�J�x{�qӣ�����i��2i�*�Mݯf���$��)RgE[%��:�	¥�&���y�"�nx^M�EiyKq��V�x�ݑ"����kx�͖����1�n�(8�gMX��33N���A�U�Ǿ�c2<cƏ����t��:�7s�-q�w�eI�����U��n=3��ǒ��(�{P.g�ȉaѯ�h��r����Jm���ݖ�d�O�/�@@dj{����$��I"n�I�q+S_mWC)��Y(�Ц#Ց�[����fu��e�l�#[��U�h:W�%P~���4
��F�g7n��B��j>1$�}+�[�5R�@�P�N>E[�n'߃��9�c
|j���)�P����@��u_B�!�v�W۞������������w��a�ߔ96M�)�Q���gi;�{s��� �_re��fx�9jMk�J� 928e�}s�N�����i�E Ҍ�c{�D���ߦꄔ7�a0� f7M��	��w����%�|5�!���!g���J֩� ��T8$����y?�yk �[�^#	�h�ܬվd��b!�e�Ҿs����t��ٱn�@{�C��/�i{�v��'s "G�uԒ����b �[��+����7*|�;�/X�4ƒ�I�p/�W=[2�Q�����`+��C/��*�O�~�!��7��MEN%��"|$84�&:W"`�X��g�UZıH�xk̊�愐��ޏē��Y,0�p��du$�7�����k#y�RЉ��n�_^m%�H����+����ܭ�U����v�| �,��n��?tI����s `��5���s��5yZP���^��*Su����཰�1M��s�w�)+�a��J��Ӯ$�A�az�O/~rF����2�j�K�1��u�1��Ю�\��ڦN��%�:܁����c�nr�;��!�I�������U1��x8n�n������Í�y\\����G�G����{&�P�PB�����)`�6����=�كͿ���cL�o�zL��}��3��]KGS���Z;	�p4��>.0(�vV�Kx�����4���88#�#�0�)���"��&߬�ȓ8�4!�����fQ[�Kt*2�o�Μ�~�Ӕe6��#\�J��u<�.�;<:���i�j}n�j�
2�Z8��Z���8�;*6�q$ ��qu��B��5U�j� Z�Ï�X��k��^�EW�DtHfNW�ʤ0�r��1�^o~~k�~а����-[�Sa�f�8�
Y>�}�Y�������wr�������#x|��X�f��^�9D�cD��?/N"{��	�c�A*���H٣T��;sY�K��q��l�T�z�Z��u�Or42�G��S�|��z�����o$�r��%h���}|�;�dܟ2��'�U!����[Nƍ������L5�UzR��w�yz�'��7�� �o�+���ф8�����zO�����!ΰ%G[Sf�Ʊ�:l���dc(����0d<.��	TP��LQHJ��6�o+�'�:�]/+w~�ڭ=y�h8���) �E��g�FQ���D�����H�Jne4�JCcJe�� ����1'��
�5%.�|�Z��A|ENټ6��!��4O��wqd�ڃ��.-U�E�������8q>.)�^T�1^1wo��g7D�ۮ}n%�nW[����|4+N����\XШǭn0��"���ݗ7���p�/�H���[Q^���w��&rm,VI.g����f��g�nA Ն��K)�����y^�����E��i�:#
���vVg�+�f�nB�]]2/Z<)$��t�I�WDػ�z�.Az��V��V3��	�� �[R��5� ��*bᑋ!L`,qV�S���Vp�4ˉ",�'��{t &!GD�g�]u˻P�=��Ќ���_�LiqRH�r�M�w4��c����u���fv�x�ǈ�`-;%�`�	1���{lT�h$�p�t;Y�:O^���e������%��>�Yz�F�,�rr^J�!nW�^aqX6���F�-۳�~��m��j��15�Ze��PIs��8���zF���>�m�0V(��6�Rb�5ؔ����sB������Q2�f�}��L4c٪��ƨQ�xP����P�!�<gI�P���ay�XN*P	րT�4v�}�!��.%+
k� ��?���lpV԰(�EJFI�t+�s6�{������̉s�0��&�E7Ǖ�i/A�	��|V7��EU�y�|����U��>'82O[dE>�/|`L#/���i7�t�s#������.s�K3�V:��BH�` �[��U��N>��4�rsbe��Y�C�B��?����rzV���R0��ҾK��l\���E-<bR�]҄[���[5Y��>�
�ĕ��<�5��k�?&���e�����q&:h���wT8J=�,<	�0�׼�|��}:K��#�H+��;�}���:��+�?���.p�U{�+���_z��Wt-#|Ky�����F�fCqb�f�Ǎ��BP}��� ��f��"Z���J��� �&�Y���l��2�W����F !�Y��^R�>�}���U $\�ql�	���%y�����ğ���%�*Ѣ=wD��,T�|�^;���g/}4q0C3���NRa�4���)�`�${��>��Ⱦ�X�w�J�����Xu�q�^Z�Nd,ͯ�}V<�{#��V!�����Bՙ|�5�j\�z���(1��Ч��e���1$2���Zk�D
���B�"�>*����3�_m���3W|I�}O�g�Q-��;6Leͻ<��e�1(��y@TP?�������aRq����'�ހf�\N��^��lԮ?]le���I��@��n��˃���$�I]�a �ڶ�+o�O�ެ���h�= �L	��NJ�����!oML<�]i�0cY��-4> �@ӭ�%��()j���9g)����T�*A��th$���>T��7+�<������ zX�2��G�\I�F1Z8�D�h�b���H�C1t���
���FB����aL���jft\w��Ŋ��Jᰨ(=�|EXd�¢C g� ��̟����uB�3R�k�!}{\���*��r�i�t��F�rvr�NF1(И�7!�ӊ�)O���|��:p�A��#JT�-������.kQ~�n�P�t[�.�P`$R>VN���Z��6Ɵ0Zn/�9�,�K<��e�fmGK�S��Y}�P��9�|�!�;��,Fh�yt�H^(���:�9N�t��A���.��Q�X\��{��V��w�ǋ��zټSv^��gi2�K�O�����mQ��ki=� ��(�FvP9�%z�(иl��/u<I��%��c�f��tDV:�.W�#�願�Dn��w;��w5z��P�P��F=�|�>�����w��Kh��@J����;�W�rx/6�
=_+#���G����w�?�kC��������Wo�����ί�B� t�jh����C���P�K�X�	u"��E��j�!�av@pu�������2��o���rT�VE�{�Jy�����7�\c-b�k�jvl6�lQՇ��҉��,�u5�~���6�K��S�M|8ɳ�!`��
_�J+���\�`���YoRd��_��ܞ�d�!�)���xR����4��_=P���pq
�GF���$�c}�X�b�a��]�z��3S������zh�C�w/���9�	�&v˛|��aƽ�)e?A�o�n�f�x�7rD-���h�_z���*h���ג��k�a۷�Ҍ <��ˋ���\��.�D:N���ǂ.��^L�>���+"rU6���B���'5%��
G��x�a�*��Sd��W�$Hc��ڮ8�|ڀ���}�m���?���g���΁�9��C��O��\�Fi��s���u +�MC���8�V�
��Y��&�Y�C��υ�tMy��33w�^�"��9�Y4�=n(?�)Y�4�Șt����o͜A��w��t�R�:; ��{W^m�큾���Tut���A��둍�˵�EJSE>aWJ~.c�pZf�[�+�������WV�gV�, ���X�5{A����	�;Z�oP[�:w���T�E݃k۸x	�AM����Y����٘��b8@Ï����9|������4��D���ha�p��f�7Hul:�Ϣ���'*����Ki�I�z�:���9"!�ř�m���h*��U�����۲e�#�0�΁�!:F�:� �A�����:;���4�#��>�Z�6~/�=F_ƒk��rǪ>���dE7�>�L)�K��#�8~��2}�����ة64��0M�q�z-��q6��Ѣϴ���N��'�Nz�z� ��I�}$���CG'{]��o��<�����2~��2�~�W�w��7�-�e�t�������,�-�J�=c�@����r��!!
�nD	���$Z�sG2cđB����~���h{�)�^��^�RB^�I�G<�E����7���P��?� �y�H���c�Ζ㪬5�L�d�8��q._�!D"�!4�D�a b�Q>�~!d���&�'&�y��iU�->�\�ň�k��ؙ��EJu)@�I���#�ٵ�i��g�J}�A 	TJ�z��T,Ҩ ���s����v�R��s���6�^g߁��~[g^á����Q��k�N{�>�>#��삝�$�y��C���A!�K���tb������\pz⤠z�XR�c��]��!qm������\	96Q�!h_\&���E��|�9��L�c4T�?҆�\@��,'�%���,ԕ�����Q;���
˾9���\3q���6���Е汪2kbq�Ca
a4u%��)�p+�FC#��nXf�����D_$u!�&Ԋ߶��gC�cפ7�Aq��@�p�3�z�b�aN��T,�[m{��{ �(�!T˝��	;�	��H��2=C�!�<s�񠻙n��E0����!�69*��:9R�"�Ƽ�ԿfJ��R~���:M�4]��L�1ڑA�@[�,HO�q_�!��_�MnЋ��.A��F�H�����Z?�1k�u���]�O�� 8�-j���mR5)"�l�p�L]J�L�"b��I�jpkv?���j�gW�N�&�J���}-y���� �[FQ�1��8���R$� ���!�ME�~�m4�Wh�.�ۆ�� cSk	]�����|a�C^�o$攪�U�o&ب=������P���1#���Ȣ��	O�U�t��0�\��܋�4}���W<J5��N�u�rY��B56�
��ꃣ�r[u�e9��U���h�K��3|�'�i�0�o����l�|��\��oz������+��J;2�)�ʦvI!���8#Բ��'8m��X,7��{��2rq]l�/��~�qu̫X-Y�����째m���Cl�[�iJ�Nc���9����^9YW�7������Q}�'#�
��
gb'��ח��m�וq
�,'ؚ��1��#�/X��;|b�6�yS������U�4�>�C+f쬟V��0���n>$X ���$���W=5�M�W�1`5���B�*f{�B��U�!<浦.K�����0���;�@�L�\	����Z��x��8L-P`(R�:���ई|-��
]I��c���|�_�j�*���Ś?��'f�T�A�c��w.��g"Y������RG|�1��������
��=��q���E�P�nz���S�������]�B�B���'rܓ�P,ƾ;���:��B�� �B�\���M'o����Q:e(i���6h�r�%璭���d>����E���8�9��w�@P2`�1A�A�wN�
��ˆ���*!1V�(^��֭����?$�qT�[���ֵ�������g��I�=z�V���IG�l����ur�MU�>�k�v�m9��-�ؾ�������Y��%,�����-��>�ؘ�%i�d���Ć`CV$���閒��u�68�������dM��>6���Ɲ�����3�c%{VX���H<AY0�Zɷo��q�Rv֋t_(2r�'�t��z�k�� �eL��x�:J9��8:�8� <@�����Q&�lq��d��h#�d��Հ`��tD�-�̈́L��h'7�`h �;����jU�P�v�z9t���;�ț������l�~��y_A��	ڒ��eP���O\WCpM-�Z�muW���q�]�N҇���Ǆ*�>����ӷ�k�a��9}��X��,d]V��1�xl��m�N���7 _�1c�$���u]f<��_	j8�g䡐��:�K��[�i�18d=��y�x�W�R�z�Y4�6��a ���Jj�ei�}�G��|���^N�c=�VH��7��U��?i�����-����l�p�!���aE��cP-X�7A^S��u4��nb;����>'}���Dt����w�x�j���QNJ֙�����Z	����ۅ��q���{v97�Ԁ���~<p&�^1>@y�U��{�T'���Z���n!�#� �=d--(�A���Y�e؏�%+�8�^�!��/��^�A�Y!s�|��,�oǜ���ۯ<|����Z�7�M��H����wA��g�W;���	k$pq��bcW���<�=-�V��U��_�X��
k�C�����+3R��qO*�c��o�,��ٳ6O��7CU�Hj�� �(9���w������a6iYF�����!"Z�Ƅ~��O�^��Y��<x�����m�e�ɴP;u�&]ے5�x���ѻ�����h����Jy�KŞ�Q5�ؓg�c?�e9?�"�`y�:
�*��μ�F�++M4^PypOƝq��Cv�
@���6������`���w�
�Q	�y��&�UB�0x����u�@˫���O��y�g�ݸ�̨�tB��G֤�T�ً5-��si駉���IvpdxR��|v�p2�Ė������A*���,��{�,g@r��`'��/�� a�u7q����7�:�τ��t��µ[�lF:a#� �g"�%�G��$�P��-@�/�3w��M��6k�%�T��	_��h��u�yb�������¢�����6��x����0�X#�� '����R*E+�ރCۼ�:��Oë�KC�n�Ύ?�d5�gR�0�O�y8�x�����%@�P!�0����>�����"}��^�� V|��L-���~.�B!�y��� � @��,}�P�=�g5�ڥq�T&8v1���z� ��Ԙ2C����n�������ޅh�u�0�E�� ��y���r|j�4{c�)D���H��Ix �]��X���6ڱ��Ż;O!��J��?Ff��6i��<C�/`���ո��+q���菆��ʴ�U�$�/��{�kټեEpC�hW����)�|QX3�7��c0Y>�a"ПM�y�̯�nF1����	��G����l�u�b��H��sqFq:����ǎ�M����G�b���92'�W(�S�:Ø�8��t0:'7j�(�Ք���~��g�~F�sj�8r*;�����%�����;Qe�r��`�e�|.�q���M��"���E] !ZP(�����}5Ț��a��tB-�a%�L��*�0Jȷ��Sf��Ð�Ә^/��G����Fp�=��GC��c�}
�<E�a�мґ��%ĕ���K1՗S������������sq�l��C��)�xx֌���IY��95(���]�t9�#6П�\�����e�e��vFe�����iQ�}�Ϳ#�5N�X�N /��H��jF�Ȇ�a�]я&�W�i������l��`7�Z�yQĹMb2o-N&T ��g�W�Kc5�u���"��;O�m	��L��7�=^���v�������i�
�m(Ȗ�ɧ2yK�8V��@�MH�eA�%�90Y��#�.C��M-�[��60���Ы���%H��;�]s.s@^��D�<"Jل�p���v]]��~�`̴�����/E�S,^��z�bCE�0{�|����Rڶ���f���v9������r��E�˂v�/��d�!F	F#E1��T`�����e����#�Q��C
�)z~Q�4uv�HOLɱK~ކ�����[PM_�ڜ�=��Y�]2���Rfc�
è�`�Q5h��K���>GĒ�rJ�%������'��G/gљ�����X7p`|��-����;��`�=�Am:�8���$1=F��}�N]�Ѫ�)�5���>&�#L�'ti���n���˥��1���|7��*��>�er5rjx+�8�Ag$��뽧���-;IU�$G��u鯏�t'�^���ƹ�-6��j�a��c�bd_P�\�)�!̽�������� {���ڷ�F�K"��)��ou�v��<t&���M:�h��k�r���օסqS�={�0UڗӸ�KfC%���9��˟W�S�|5m�:τƛP�+�BOz��L9��xH��iN�+Rj�OY���{UA�K��!�I?�EЄ�^��[(H��+�y�q^� B��S�J�ni��7!~O�L���9����O���ז'8��*sP�Ӝ���y�^vW�B苲T�ǦB�K�뗫��@�r���XWa�"��i��Σ�S�P{6%r'm}t0�xq�����8����E�g������	7�6� tނh�m0��Ȧ}�{�a�������Q�~ž�T���t�/ �O:��bsw��}�w�3�z�h��~|&�v+y�y� ���2�߫R�	UI������:�w ¢�枒�y@�L=�^ڧZ�k�o�z��(�3��@�p���-��t/���d�]bEtP+ +Ĵ�"o�L����:"(����.1"��EM}�����J�R������B
�%#ڽxe&zNW�ٺ�U�}�&�V��Dy8���.6��Hu�P�xd��5���7u���q3+OdiN�p�_a�K7�����H���1{�S�ɚ|����`a/��^���DRڏ���#gʫN�����Lc��C`��늂�e��¬���_%�5'ѣͅ�.�w���mpD�����l	��xmo�+e�)��g����Ҳi�@���-��֬MU���:����Q��r�����)�b�Pd�?�g�%r�8+dqc��^Bx�G��xu)�r£�A:����Ӽ������S����2:���@XKOv�4�鄸!I�E	�������\p�f�$t��,ot,sE��x�T���� tv��dO�ϲ������C��Y݃s�� ���Z�zݝ��8Vs�����`u<�.h���Y���.K��{C��I
�Yu���|ֈD88$��S)��<T!�&�y��]=O�=#X�M/I���m��.����O���Y[�<�E'͒���(�P=��i�B4^��Ē,�߷����4A��
���K
{� b=b��n�f��T;����ޔՅ��� ŏ�~��(1B̰��g�E�6�L�Aˠh���Rn� ��K��pd`j$����3UH^*t>��#���= ��l��d$0���l�m�f$l}hiS�����v�`��gY��~�i9�׏�k��@��&��L���)\��:�6=��֝����
���U9�.��=�/������(�9ǱRr��v�;/����62�r�o|��g��j���m>�?��.�Sȑ<G����&�ր'��M#a�@�5u�S6��L-?^��
�QԜ�EgO[��p����͍A��S�0���O���^^C�;��kO\��}E�8��8��v��L�{�%|�.��s�#Θ��6s��Tg?�}W���X�"Zk�\TJ��� 4c�?��Zb"�����"k�'Ũx n�.Ō.����K:���	�����J�Ѣ�*\������S\�V9�ұ%j?���[�h���6�fmdD��4��o�Ygt�l���_ނR��R, � ϻ��c2X!�U�`̫Z��#�b����T��o��p!�Zk�bd�;+h�D����]^9�AHSgֶyr-�e
��� <;Io_��σ���PL����`�m�^"Iu�'A�����7����r��{��3�)-��B¦Hؿ�$��!a"U�w#� Z�Rd��8����b��uz��>l�Ӣ�lĨ��9R����[>���-��xq�z�
��C[�� \������I��J/�^-�m�|��A߀�wp���\e�%��bh�f��UC���s�g�˺ �@�\������΃�8?NV���i�	(f�;�)�6�y/!��@�{�։��IC��љ��Ny�8�UB����u��5B��d���N�œ�/N���@v]ʦ�s�؃3)��^V^�7H��ѽ�ș�����8<nq�~1�j`�u��e$ S�hqq��z�}4�3�;" Gٚg��k�P=�}ءj�W����n��n����t�Đ4�	ĭ�q������Cs�ۢ���b�wM��pآ)(|E��ډu=,B�ѭ��X1A�ͬ��P vu=��]�iÓ���i�+��!�
q|��Z��G���a�\�ۥ��L��Jx��K��o�� ��!�OXÏ�ji�l��H^z��D
��WgD������#��/��U\0�����Y��P�����%�V�˶F��x"�C�uY�P6�_k�{(R,�u��jT/8���4|�b4��
%�HW�����r�'� �Bq���a �W1�e%���,M=5B��>o�����ȽKq���}~O�*���oS�r���g{�Ö��*�D77C���c����������6�JU��~%��Z��H���l�B����\�CcS������~��$}�.ѷdP�RĽzkk҄a�;i��5���K=���	(���둽���Oɹ��7T���
�%�t�
-id'��^zT��x�qC	�h�-�7?a��rܞ	�����Xx�M�7����ڂ�m�ypo��K�Y��z���p���:F��$�&H���da��7f������F�҄��7�)��� ���b��;-���[�s*Ӻ��^����,��v͞V퐎֖	n�16���:I��4w:փ���c��i?)��"�+U�/��l~���VFHX�" L�ſ�A{���z�5';%r���[p�C�=�lrG-��w{�k���N����<R݈M�B�~�/,87X��r�������ZY#?o�y4'����-5�JN5�X72�����$>D]a�]��^蘆���yLkRk�]� a�k�P�VI��g����\T!�f���Yl�H"h�Q�Z�t:<^�4�u�b�-��Nfz۵	��J �����Z�Mѫ��LKRSl��&��36+ d�v������<ծP<�&���K�O�V&�Gji�Y 3k�����U�g�Ⱥ:��f���11�N 	v���C�6J�\S*�N83�@X�:�1����,���fS���<#�g}�w�5�������w,�m����<�-�i^2�L���T@ONۜ�����	7�ޝ�J��D�+�bW�� MC��(�-l��?![�!��\#�(^�*���0� C�ړ�z\u@T�F�B�`<й�/.}�	Ha=�[�� 64�U�%��ԫ���q��=�5����)n�IT�����w��`�6�x�#�DXXSπ��u�NU����;;�4l��8�-P��9C��Z/乊�J���=
�0�ug���_��{��j~�,[�n������yU��v���j΄��U��9��L)D��!+^������BnC�������]ܯ�%掂kw���������q"?�	Wپ$��ϰ��MR�󙡧Ɯ�s��&q#N����D�_|�b;E:��������%Ɂ]��]Ry�z"��R`����T�r}?�S6�\�!�Tn7?�& �\����Rz9F2� ��h^�[��� q����۵J�J,]�5@����~�����Wx��������o����fjN�����o@l�k�ϩ�$^g=�*�p}G@%�	�he�ƑmX���XWB�|�:�a�bQ��\ߡwfg�'��6�o��3�"{��c��]�{��M��ـ	�,ۇSJ.� PR�{҅�����>�O�l��P��,81F�ͅ�?b��oP�ThMo�(l*7���$��Bv�̠��k$��	$	X��������߾iu�4F�c��S�|�զ��=�w�ILr�^��M;.���
;�@���n�wb�M�V*rd�\-�cv�i�wNy��Úa���12-9��|E�6;�u�*���I�v
`1����㮢u1�2V�h=���נA4�+� 2 ټ����,�"�y�@�`Eb�u�զc�#�r�w��*%մ�cH��PQ�&t�i���4���.��g�NQ�T���5-�AE}��%  ﺛ�ϾE.�{sW��=3G	d�&A�^�
�M#���IE�ޭ���3>�6�?!s�&V�C�Q��q(���*��[�ۙ�s��*m+����0���$���Ͱ��+3��|��J�]��;��4A���燳�<�:`hTȤ�f���{x��l�~s�K�f�+p+�'���M���0���w�|���������홅np1�^�m���-�c���b��C�K*2�4�%��ML�}r�T8�?������~ڐ=��h�xS���
ZP�1�	���t*�������0'����=��d��n�	��,�G�W�8)���!��^���F��0��lK��x������̝v��
T�^���N-�=��RƊr�@Gt�\��%N�����:Ǎ���i��]�WY~�i�\���P@
p^�+*����)^�ڬ�kÏ�}j_��Io��C\%���h�?��U�g��w�9�k�b%AQR��B<���#[�їi��:�Ғ@�Q����G��"�@c�rDS����oN������xO�_�� �ʚ�B}�e���|nw����j��M���*[W�0�̢]urD���VD)�k��݆�֎�9H!�%Ƥm��1�^F�7�is��oIt��\�ณ�����z���!z?(׌��~�v�7Y�"����7+��'P<��l����1��}�!�/!�a�&��&����_�='�����Z�}�OD����c���$�פ̖s�ȆT���!��R���u��å�@+<�c"Q�q�Z{BP�kN�$>���i[9�n�����`���^K�U�����"ٽ�ЖI٫��Ot��@=��䋔�X�.�{�~�qP�^��p��w޻e8x��=�CA���� 
|�<h*�T��ֻ��g �)��iᬲvX�p�-���f,׭���6�'t��!�^+�J��e�����VI��6�s�F�����D���MQ�V'n(^)��"/�-s���Yn;�߬�6� �a�8>bAW��CO#�M(��^f�ZE����b�^���kv*�mtwM��o���s�����|?�x.�t������ ��U�sc��1sKJ��^����i<��F��@�ZT��\^�OBp�����:P���iA�2���(B�zi��.���h�l��J���gl)�C�-�ȉ��e:�nD,%�W��D~�|�e����\v�>�- ޼�n\_�]�%�ϝo$:���8�(8�����x��'�$y#�d�D�'v���_��y� ��)�J/�Oz.D-����U���Po��3�Ι���"$PS3Z�߁����A�E �&���gђiq�W`]�����Oiy"������B�)g�O	�W"w�D#ᜑ��p�R6��'���:��@���z��V{��e�P|�g�h����u�ʛ���
/�:�G>}���FG*���u8�p��@�dWT�}�e2"��6im2z�|v�obM��o���(��C7�vfg�������2JW;�Cfe@܄�ç!�v��kH�Ȁ�ݡ�\����߸����x]��<:�^}��3���{���S^�o5j<'s�_������qYJ�}���q�9��]�L{�,Nk`!�x��jb$�!@
����?V��)�_�G��Vjw:,���M4�A@�Z(Ip��cs��g{�#c�W䍸��m�� g\q�V��e��(��l�"�>���H:����/`/��ff�̭_�p�ȓ��7V;��⁶���a�h��a�����Z$X�@�\�:� ��#���z��W���
͋b�<Gu��Ӂ���V���Hɺ�jdǎ}�"�lkE�䠛�lx�+�g$���/{� �U�is�	�9������Ǭ�-��n������6h��k�eL���q6Y�m�Rz6�ӕb�M�g��ۀ��|3�����ˁ�8B�@c�1���?كa_|�d�ϐ��L=<�?a���N���� /����L�;z��Z��Z�2ԁ�h_k�0�a۩㎫��8h��>Q>�rE�;)FX����GO}�3�C����=��T�`�U���l0gH+U|["KL��u���2�M��rbҡN�zB��SR@��]�I������B��|Z��HL��̪�/.�ßv����b(յ՜a!�{h��u+Z3D�<�a��8f�^������ZH���oW��nP\�`��)�<%'�&�7X&�6;�VJ�uI��N��H�}�E����iI؊��̢A��� ���7<��U��];��x1��Y��qr��|�<z-�+sTs�,Y��G�K�S�"�aj��r��}+�'L|�{:��������	��q������5%�>�ּ���������Ma�n�m�o^Pt-�B>���s��5�HW7+.؋K��V��|.2�&���HckH=�`����0��DA@��a�D(���:&�gEU-YV�� ��5̄�ABs~ +W�N3Ҹ�� ���nAAX~+�g +����+��2`��ȏm�k�A�@�?t*���n�K7�Qf��6_�����4�B���^hY�'�����[B�Foνs����]�q+h�ЫwMi�ل�d��,[Z{�Å7�������`d�q���GF�Q�����s��D�ip��vvNh��CA�ǈ+�;�e+}���(��S��jv�G|�հ�!G��(�D�֌6��%2))��i!a����"�8��H����tH��C�O�����Y��H��|���Sƿ?` ����6d����5�~CZ?��8��-��W,�oM�KFp�K��N_pi�ֽ&OY���.�^J�sl��n�6�3k���%i��燄�X�R������u�U�Z�P��gڞ��:��2��<W�k�v	~.۬P~~�@���tK��_��1�=b��!����I��SW^R#eU�$�m��ebӨ[��(Ƿ�aG�`�$>k辶�"�M��г"V��:
�p9��V�W|N�|$�ȀzY�j����Q)E��6�Ѽ�{��hT�Ny���@*�e_����L��8�^.�<�J^vE�G�(�����9G:��� <U m>2�;4�s��5G�-L���	�������O\j�	�p��
�cх,uP��O����o��	�~d�����F��m1�C�&��oU����f�K(���N�	�������G:C���Պ���w}���q#a΁P��z��k/ϲ�ԹoF��P���:	d�r*&M���� wꙹ �T�ss����V���g�W��(z(Fh�O�X~=���U�I �b ̶O����Hs�R�+�A������c�������'��� ��":��P�W�+��߷����/iP�Q�/sSpq���;^��(*4I����)B��Ψ�����{����Z�,9ML���=��L�������պ�i����'~��$m�&�]���4��#
uD�w�[�'�JfMq�Z"�H[R�Z����"�|�ͭ���GvI'���JDO>,�!2G�H���}�i ��\�W�<���S����f9���+wa(����N3/���~�W�楎ՖY/��E���-(�ti��c�����H�ϲq�?�=�����O���eo�p̑4"gyX�ۘ�G�����'j��?m��F�6���*�0Ѥ��ku@Y��hJ疗bU���z�'�(S��Nm��ũe�-�)�<�4�&8tY�b���'���sT�~Q�x�����b��DPz�-w����t��k�����A�Ď�=;h	����n\"����6��3�T��9"5�gd��Y`�/��mz�(.�'�Zm��h�E+�s�_]��y25*(z�(I�%��Z���eZ���:�Êѵ���W�,�x3����4y�5z�����G�&<4��Q�l�;�n�K�g��ob6Q��HT@��ˆ��O�f�!�{q$m��vЬ�g�B<3i�-9U��;�E�S1���"K�H��!Ě>kId���\ϡ���lJ0��߆��
[�R���lkH�=�U��������G��ų��C����Qh}YV�����i�������È50���LO!����>��%���M;�6= m�R�t�N�8���O��>�2�гSB����5���~DR�m<����s���'� ��w�Z�tr���_��"3a6a�%��K�;�Jn%��Z�(�I������w\*v|YT��lCw����r�*��jEci�\�����[�f���{�Ke0�Y�����s$Ud����2ۏ3��*����5�MJt��y�p���#\ڝ�6���5�S~��bb� �F�����g��z��5���6oa�8%}�L�ڷ�*7<$�e�q�O9o}�zO�4���%Ep}�F}/��/��[�8�,����:����/H,&�/6����k��=m�IV��"�*m	��3L4'U�k�\Nw��vXM^�?س`�kߎ�#z6��'蚱zD��1�թ��>��	+��N�����t�[��S���p	/â�9;���|��dx�t 
�дk^�Uq�(� F��Z���%�3j�O:o	���3v��O2������+���Wc��^�����q��ϛ���lŢ]@F�KFӞ�WH��	��[4{�\ɶ[G9q���&��\!��*��k޾̻i�S]�!���V�,4��> �3ˊ]�s��T��i�����?���2���c�q}�j?	J+:��k��cU���;ybۨȓ�.c�"ĝ'������!3A���s�.;�b@�t�a�:�v��g����nl���լ�^�o��^�_iW�D$PP{��J��3g��r ����٭V�_��7	��U5\�\v_*��#c�ڂ��z��������f:��X^FҾ���a�!��qf�ց���.%,MՒ�x�̄/�S�IS�f��@��-���/apt1B���ȁZ(�M�&1��
TЇ�_
(O�H����d��z�5���͎O��Jz������8|}l(���k�����y�E�Y�ͅ�w�7/��ypE��j9�CP��a�@9>�1���
�P����ý�X�0����"L`9�W�8
݈���bp��kD����*p,!��cK��sʜ2aAy��V�M+��M�q
��=�,�#Df��Π�<?e!�S�-��'[����-��k~�~��E
3��J��tU�e�ʹ}�>q�0���]E}[�r������{��-R�b(�h�Ǌ���$7��^O���7KN{[{�1c�]n���=����Y|��I_*�Ѐ��\2�����m4���2ˡ&8�W�Css�������(��pȿآT�nnHl��~a�ۇ��u�^�G/�鯸�����H�v��,���t�P��������XDS(t���x*(uM��GͼB���87ϯ������6\̅����a6,�$MZ�D7��M;f}�S�G�1r��'�Xl]�̵�viϽN�\����Y1U��V	EJ����_㠤�-�֦֥��WS+��I:҃P�o'�y �G���)����7�i-CXO,x����|��� ��fN��~~Z�t�B k�q��>jfT?�WV�q��ʙ ��a��zP�ىaD�]��u������+@z)��=p�N��k�r���'�p�Cߌ��L�&���%G���Ҏ�Xqg��y�=���QT{���_V�"խ��Ƙ�C<��e�5QT�8�KB���޻R!" � �)�R�L3G��'e4�ȪO�w_��r{���[� ��ǆ���4Lr���b��_��|8�b_���'����J�����hd��B�MR0�q��J��z�X����=�
j{/*>d�J�-�9��$�(��`~+	��[��H�Q|5��,u��̋�Ð�NQ�QF9lZ{�eb��B��'�%w��J��ΐ�!����Vas%��u~%vL��.��_��e��=r�66��j%Z��FPG�G������[�A��E�+�f�����?Փ��,�����Wv>�����\�V'd��c��	�gi;+��<B+��-���4OY �.݋�q!�&��eܗ�r��h��F�0� �Y���L���[
HK�m�F��&�%���B�W�̀�����{�ͮ)+���7lD!^o)Jc-���=�X�v|$�y FZ����[�ϥ?Q!E
�#3�bAl��>l�i�eZ��+� �/{�4���Va�A��h�>R�+e'��������� �����f9ݧ��v�k蟑1�����=�]4���S�a�|b-�I���/g5���%�c��P򜺩�o����˂��n�M8~�W5����Љ[5�8��~cI;��,73�.�޼&����s�o�G�ڡ{���0Y�2�O�[��|�w�8c�{M���U>�0��4����d�S\O���>�ɍ��;(��l�r�S��xi.}:h��3��YBC�X�H���qţ�<� �zfrmTG�zw"��/�*$L�K����u�Lih�Lv.K����[8}�ħu�4O�.������~��w�츸��͇l�a��Zb$�7�z� c~��^%�ӻ�N"�� # E�+/6��-
m����C�* 2H�R��8-����=�ܾjf��䩺���$:AjԒV��N(�3����>�݌3@�.2b��7L�X��2�E�-=XҊj4R�sD���qv��>?��]�'�Y�-�<X�֘S��-@�]�X���9t>3��ww2�a.��&��v��d�6��n}��/��ORU���ߦ]u�K�t�û�ƌ�x��ĸ��[�Ͷ޵a���N������q��j��,�@�Y)���<��|��7+����,��$d+]䋌C�G�
��r1�c2l�5~��8P�lL,rn���Oy�I���2ۻ��	����ZpCZ~�KQ��};��u���T�bn!VI�D������ gBH�LZr��h4B��wH�9�}@;	eI�)��x,��v�:?���Jnr���.%�ܵ����W�0�{G����s��Z���D����6�IH��g%����2.1��A�B�MeGG���}� Y�tx"�}��ȶ��	�A�"��f�����5�z,�\ή��S �n�V��5PS�ԝ�<;�;��fwE�.�e�h�rKgtO���R��ܫ��ٮ� 塉X�Q�[��ˀ��d���),�6A����8�7I9��.�a=l����@����26yZ��Y�z�2f�[ߔ�]u\��{�Ҏ� s�k	�xl�R���h������E���({�]��&,Sv������ƪ��	�6'9�=aZΗ���ˌ���.��&��XM�'`C���	Gf�+\I�y�H?�u? ��k~u�;gW*� ;�x�2 ��BF���Ė�Ԥf�O˄3��
)N���i�G��0c�ntW�T�J�� �p�C�Ȋ`5Oa�dų���镚���Ѳ�V��-�4)6ò���M)r���0ǁ��wy<�N��l���[:Z�L��>yb*�Xs9�C�FQ<��6r�P͒��E|6Wb00�Ϯ t46�e�z;SO��q�f��]WD������4�<� skS0̩�5������S��jK��;��fȈ���Rb�M�Ό�W��k�6����+�W2�k����D�E+��_+���E~���w�y׃�R���k�"ԲR��՞_%ƺ�b�>�5s��mVW�'���K��IM�y�|�� ؓ4/�x��U������6/����)(O�:��US�u�`�"V @3y�A5�K�fi&"�U�W܂�'R������(�&�ˈ�^v�fZ'~�V	�8�2�Д hĮD�<%���CP�x�|	c�%��ή��G�ޓ�y�'E=xu�4���I�$�щ�L$'�蚫~��6'S��Ǯ{�'�*��%os���c�k�w�t=×>�*��h���{��!��"��[��D��<��JנyDd�X��o�鄁�&n�lkYT�{�7f���j
�ly �s	��W�5(����Z��\~�v�ߋR54���2���.Y9�#�h�_Rm��kH�]��V?,�ue@c�B��� �f�����#�[hkQ�` )M�T����Z���,9!��t��!m�[J/l��n5/B�5�E��&1D����P�Zo�Is�c2���4��~.�qhR}eM��C��*��	��dq�_�C�*�$r�v��֮N��7�g�Ab7��~,��$f�O�_��[�
�{�l����S���yt����3����8�v��DY��~=M��Cÿ0!��E'e�S���k�)M�l��[�l��Y�%��!M���3���0Dåsa:�삫���=��K�X��g�2uH�s�#s����y-eu/\�3�`�p���!AN�3�-�S��a(Ѧ�t��Y�8U�l�n�ᥝ��o�9������]��M,�i�>�b^
��i�f��@j��Ai!	��z�C�vz�Yh��.������ N';E�O㉭n"T1�q�8��q���IJ�x#Ki� s�9�.!���BTc�<=�*���l:>��.�=J�_N��mK��e�=V$��T�������:�[yD����H���Q���	���� �2?�2����B�#���Nə�Yͭc�'��1i_"|�9x[�m�s��
�K��>� ԗ8#W#6 P�	}���?4J��um��à���`D���6:6Ɛ�B�d-oﲮ��*e��Kg�zL`4�SHs�ٔ��m$*ͭ�[��݈�F�v�!�GK�\��䃖6�ꗭ(�/��{�.,#,�F��ܪu$������4qQ����>��@�yg��}��gк��$Q$&�%�����|"g�!�Ʒ�BeK�;��k52��\����:�$1Zg��	<&Uz�
����g����yQ:܅��܉h�Y Gd�d�����e�;���D�`*�>���)�o��0o
�%�������i�ST\��k҄f ?�I�X(���~����T��cd��r^��
������n�Esf+�����nR��ߦ����u���'�|T��r$y�;Ŷ�N��`�jR����S�-���	Ւ8Wp)�y�yސRS-�� >˜�}��[<b�bG#�?��t�2�*���7���7�Z]Z��0���d�|��.��N�!v't㗁�5ơK�M9����Z��⮒�2��}2���ܬS��m���8/*��$�ň�OM�H��꒫*+j/a=�,M��G�N>�mSY6u �EFa��Q�6P�_l9�oQQ!�ݩO��@`V:���ge�4051�<4���ˍ��e�4L��ޥ;~��=� ė�5_a�(>�;A��D���iҫKGa�x/�ՠRI_��<d�)���E���<J~뀄sYMs��voK��l�:�Cey��>���j�$X߮Q2t�(�X6��C9Vl�T��.ಣ�r!��pY��H�� a5Y�f��(;T��P8�{�V��,uvDp�HT���.�i�dfR-�O�0�W�mѷ=���=�b4D�'�~2*ƖO�bC�ӧ.��7���O����0�q��_��~"��M*C6-�u)��E7��`ٍs�7���y,σŒm&Z~�dY:k�i|�#m�CDqeg�;V��XW0�����ɔI�R�_}��+V��f\�[VY�����PG�����"=����e���("R)�^P��PKUs���;5�B��*��Y����T$��|:y�$���#��pC^$�aQ������Y�IR���y�hP1
���1��?D�c���k�C��9m�у9���D��b
5!h�(]�9��?Zu��Y�p��x�\��/%+�$�<�J�)/�]�iɣL}۹�IĘ���Pv&~q����1 )i(F��\����A^[�4��)�>�0D��M��q�O�& �nR�A��b�x�Rs�z�8�t�k y��Ԧ�S��We����Kiw8�x�ٗ+ M��V��{z����cXc�W�dRS�����8 �Bb����R�c5����� I�V�>�s~��V>Y��<�q�a9[9����SBe[��r/~H�����wJ2?{��0���"�������++���p�g������V�;��.4cJ����I$:�_&����&�J�HŤ�r ����C�I��Рw���`�B��T�'�&�a���J��T�����h?f3k�L��i�#Y��ZR^�-��!�����S��/���l|݁�Za�]�'�ѿ�p�B4ͦ�W��IK���T�Oi���?Dy�l�b���h%V2�
�����	��u�u�B����BC��Bp��+��5{��n�YĬ�T�bڈ[��t}����-�Ԋ/�� ?�;�(&@��|2AL�3F�y��<)�X�S�"f�cy��\u�q��x(%ԱMO<�5c}�ڎhOR�Ԙ3��R��9�V�Y� `%�k��5���ck�W#ǛF�Eي�����,�+���&��`��}H��yS8�� �K���`2ɒ��:Ϣ�*��|��x�I�kf8o[���p�xȔ���LF�$bY�^f�5A�s6|-=R��7�"�`	9���o�Qv�_J+�A
:��܎*�%�wz�cѕ�����:�7L�-��B�ʗ�B������K|W�U�0q��(,:\m��w�UE[y�jq�@bU@!C��y�b�`/I��*s�;��Y"s�^Sk��a~��g�po![I%��B?)�VPAsQ��J�U�b�8�{�`���|�7���zR�9��O����%e�������ʆCB_'	�v���C���^ɉ-up�/��=��!��7u�T��ţ���>C<���pL]OI}�=L��(X_����v�6�yȿ�e�n���_�f��f��b�Q/��\rc�ۼ�R����}$�NY����0����.�K~��	�+Ť�����1l�����0�R�z�GEnY%!���좭WA�46�N�k/i�3��H˨{YP��T�U��ݜ|RE�ʢ��L���Df�e?�D�Q��/dX�`�h9~�HeS��OttXI�|me��D� �2T���x{%X��+:�d>*�g�@C,���dJx.��!���Vc��,4��h(����Ve"?X�*�g���C��'�\%5:�B�k�^��rN�YL�A�ȁ�c����{x�����j��!��-�g�j��&��'���s����6�<�־�E�}��G���(��.�nѶ^�t���'W 1�5���	%�R�79�v2����x�%��O�G����q�m���7�"��6Sn�t�jG���%y@R� ��Ɖyg-˕�7��ꍚ� ���-/��qkI�djh���2i��އ�_ڸŒ1gx�Y,S���#^)x̍��sЋ���5cM��e���;K�x�r�Zt��E%��D�7�0�#+ ҡB�����@��Ζ�f[�o��跞��+87F�ݥ��=��y�*��p�L�M�U�k"�u��}�~�����b;���ҙ��i Y���gll��&��c��C��X�1"�ź�K&����7s�����?d>����b�;v4m���$@ y\+��ˠrȥi�^R�hj(��=��H�c��}��D!�%��u[��ų:z��+�vd��:+������ m��eYt��0��[��X��1�5T�bQ�X���2�?�K0�cTݷo�!
��Km�3���3o���,�ɾ��;.s��Uq��m�e`�`z�����:�YH*����X�p6�{%h�"d�8��-�2a`L��G=�����Uj��sy� � �y�JV&�����T�h�ym@ƈN%J�C6[�\�*�ep���=�D�z����~�[�����G�v��|T��]����A��V&�G�����w`s9�m���T{��u\�9�=�_�{��b��
��(d��.���Eߋ;���1��Zx�n,�}|�MƘ����!�o�x�O��*q��B�R���&$���zj+���ƅ����?B$�=�9 �%��~�R����<sw2f;��@=�y�;~��וl&�+������`������X N�,�Z[K������0��FȴUy�� �]���_�8���k8���\�K��g����Ō5?P�i�Nȉ�G�I�v���B6���/������`U��T���T[8�my����n
��av}RYR�,�:����x'���J�,Z��Z��_7��u3�L��#�v�y�B u3?Zj�d�[�͋7����D�R����,���r,����}�+� �n�nj�X�5	��߂�Rf��I��?�H�\����W՚��0�87N��v�k�,�H�T�"��~���}	����Bo���e��׊�/r+=h83��Y9�x�Ÿ{q�? �c���"܁\	]��GB��VG�����l��IX� ���oS���Vi��p�l�ƙ�ˤ��n�8�ȹ��aK�3���Sc�X�!p⡀�H$n_a/��Fru��\�ik������Ö!�i�˃�^�Y#���(�]v�~q��X	`}�^��a1
Xm��f��.^5���;L����rc+U���z�����G,���.K��[,���l6�O>T�T�=��N|P�9�W�'*.wZ�@�@"�� �cy�?��R��q�*��h�Yv#���jW���9-$9
v�7G��	L=S���U��N#�/5�]vK���:'.&�MV�>�CE��4�����îlp�4RQ�'���-�׭bϧO�օ�5��X�3��˯�b�h���S�;���µw#9୹~n�6�I�F��E��Z�)�AygE:sXT:�?k�\ɕ~L:?y}�h��9*l��zЃ���A�Q���.���u�02�pW�%����*�b���Ȧp�"'͇�<��X���0�-�{�V~)w�9�*p`,��o؞@��pb�7W�����?�L�k���I�����޳�9���_�������--����1W��i|�M��ކj�o�j�P?p0�u�6Y����tϓ@�x
\e-�C)��;����8zS��KG�^�ƹ@���.�!�v*�ܻ��Ld2�6���Y�flm~���ɀ�V�.��8Բ�e��Ԟ�@��>�K��@��Pȃ��3 ~fCl|}p5hhXkc\yJ�
�P4�~'���[Z� �P��}�?9���Ƿ�Bm[�ӊ����k�/�����R�9/۫�.6y%�v��r�FvmJ=����xT�S�w�1�Ur�@�ՔD�(]����4���U���fH�Q��Xԩ�z>���`oL]�!�6�$S
	��X���[��<LV�KMLC"���qv8����.�.�Y��@d��ȕ�5�EP�m�ǽ�Q1��f��s�0�S1i��O2;�$�S[����!�<D��d��߁2��6��"��[������_�>hc[hN�rM�jzSld9"��4�Y��$��鼀/�b�pf�}�K��I~5V��K�s�Q��w>ǂ)�,�q�ι6�o��+׆a���K�o���1�u�g?vc҆P���ct��-U��W0�"{�?��a'��`)���8\
:���6�W��ޣM��	�G�d�h(��]e���p���s�#�M���ѣ��r�/y��6�1U�R�aTǥcҺ�9��ġ��������sP�y]O�v^��|��1�d���O�nh*�c�<�GC6�t�W�jUz�gՃ������B/Q�P��r�JH�����
1n+F��{�Q��eAw0��&nB�ZJӁ��W�s|p"M]Bz��r��f������I�8Z��\',��1�������RT{Q<U�t^��$:����{��0LG#����^�����o�]M�n��[W��K]���C�VG���w^�?�L^sd�bF9��Ϲb����;O�z�E8i.8y��_)�ME1X��4�gR���Hrb��3�V�4����9$)����7�}�)��'���Љ���k�d�F��ߔ��ǙU�S���o������T�ͩ�ۡ8`�� ��»꿞%��3��C�i�6LI*�h1���>��Q����5�:����0�2͙%!>���(�r�-���7��:��cϦ���u��������,��b��J'�=����N9n���n�,�q���.�)�V�5�ׄ�k͌�cG��G�,�"��h�"P�`�0���J(�B����NR�	t~�U���q�!v�9n|-f�f�: 8bQ  �9�ڑ�b<������]�ҞG<���1�s9^�u���T�J}��m_�s�؀��	�W�`phE
@'�qi"��x�Z���~h��e��6�O�bH ��WJ�ax��J�"��Lp�P��`zAV��&��on�1K���E��m�`�2���=�E���a����m�f`d�Z�V�����#w�7/ݸ��
P�J���c:^9�[6u���N�bȮ���y�6$�f�/��;���2�~�V@5�*�%P��&��x�1��k�x��N�uc�nW�V%$�`ʈ���r�z�%�iy�Bk���y+b+�!�*��V���x)�2�==.(0ӝ����E8�9����~E�R�_naT�o}��Kf �WCbz��]j�'�Ǖ�:{P����n�m��������B�5B4��Yyk�/j�~S�(_�fۍ�e��Б�).<��h��:�J����Jz�m"�dor�2o8������0�v��eGp��"���p~��2�9���-�-�K��P�@ٜ��'�09x	D�M�oh�|�*B-ON�6_��sA���S��~�
�D��;ܠ6f�T��Ί��{�i���,��)���=w
_K���s.�M��5O���@nΖ4Cڬ�� G[�1�#����q���6sIW'a�մ�>|J�ڗsG�q��jI�0�4��Ł�����!�����'����/m2�� �$� ��e����;�C)���$n �1�h�S��cy{�����-�?Whq.�3�qv����z���   �hN�����:�th��/���ę!#B�o�҅|EfTp$�g�`c,��T1�D��5ܿ�G��<�It��h���oe��s��jyDږ>;�L	��۹%C*kq�}rHB�K.� lua븭h�8�0ol�1�X15׭I��Q.P<���1'6Sٽ���/��ަ"Z�q�p��&2���@uɂ�qð&�s� �����w������N��H^�k'Q�Y���9��|�V�O�k��qB΄\�F�����X�Hx�E��:�"����h 2w�euZ��S�o#͍�w]�tX٧=��A F�R:"�^EJ��"�T�Ué{ɺX�d��O�R�$�6�#R��\�����C���w�u/�y�����&S�\�ߔ:�Y	h������6��uv���I���-�'EGj��«�=�p�sa�oH�Yg��O4*�����"��6Af����i��ƪ��c��x��o��3�o��Kk?	�C�m���)5�"��P�,p{A'��L�h%�ư�y"�s+���BK�o�rH��m���J����ȳ�`���B	�{�S��3�=S��=<h: ��3�)��qU����>��`E���P��}?�,x��&����ұR�^r�}�ʪ�Ҁ\1�5�~2���D`�����Ye��fJ�����5�ՑM2���;�1��o��㧥
��
=#�Y�h~Q֩�H�K��ܞ�a��"�}>�)T��'�n���$��R'F����m	\��k2�3�X������~7�bH��G���7�`�l1��_H���Ҝ�ؤGqi�P:���g(��87Ҝ?��\I	�&s��?��ު��>I�^\${;F����P6hޒs�������v���]	�a�a�&�����^Wc�=�pD8�~
�������1��r J}׫\���)V1�=���f��E �	����c,�'#Gl:�%TQ"�:w�6(�w
��
����buV�~���h��H�k�Ӄ��V��S�o���.��R��P�H�"�'�"�EÝ�d����p��"K���{�c�ِ�~����I�h�v��T��{�r+�([��W.�<˺,8.�$�]h7�Y��|�I�?�y4gZ�s
���[z)��8H�pK_��� L}k��Ã��s�(�i����|�
+�1��Ӥ?�W��r�A̡�j����5%�N�m	�[����C''V��	�.��2���G�=^6!���3�zi�P0A=LqY�}]�Ȗ.�����xth��7�I1��D���S��t��B;T�i��&]�	2<��ØQxRw����-�����n�D��a��ΛK��PS���s����f�i�ES��m�P<���|]�b�S��\���&���z��c���������Z��c��#o&z��w'OP�����+DW����=�Ch��`}�^�f�Rn ��{ַ0�B�����=����B[������'����B?�_H+���a�#fZ@�$◻�_2HQ�K	�f��S�ث_����Xl
�㊬�H�Ҧ&��7�y�4pҎu��=�aA�(}�5v[�ϗD�;��w<O���'8�v:E�Ȼ�f���Z�^iѽ"�����Jh������b�zs��$G�79�5S����h��	0 �&x�����x=��0��	�U�s��*gР��㟼r#���	|�n��B�4����?rop�Ek_������NG@2Z�����_���B�����������8�p+C�ն���A_�Z�"�}�5����x�{v�s膐ǔS�=�HM��Nh���.{���Uw  _tj��]f;�ͩ�ݙ',�o5�x��xq
qɳa����G�F+�E�ze��)	�[v�>�5��y�&}(�z	����-1��D.�Jɀe	v�>�7s^}��~[o|��r/~/��!Hݖ����{x,D����������Y����pل��<w�,�W��ϴB�$_ٮ�%)~�y�}�`�9��!=��Jf�.�3xɷD�H��2��P����´�ș��F��"v /�%�j߆�H�lx�sӹ�HR�܏ae������Ԑ�S=�&�J�P�!����PV;��qZظih
�&R0�`���cY�J,
7��{ӾQ����2b���+{�d��� N���dZt�ou�MF��l��}�6 �	�>i[�2o�n�ތ�〕E�4U���[l�5�^��(ٙ4gp�EP�f��9�� �`�B���fe7!V��{3_`��.jߕ4��vw��Rႝ�_��=�GU��ST�Լ&𺦐�?����T�K���5|��.w�ͪ���-��
WD��Uֵa\��M��2B�xH��|���u]S�aT����#	�lj�����6V�$�ī4�x(��=�a��#lZmK�xGT�O�&�	����zrN`�_#야bj_i�60��_4���ЛZN4�]U�ꍆ���c� �}C�B0V�Z�J�e:��it
&�N�J�-0\(�՛@I}��b���P��Y!:Ν $Ѓᰚ?�q"�ycUNMj�&��b�FEg����E��D�X/k�`����z(!����4[��ډ����!A1�)��u����N�<AnA���_V�[����kx��x%�7q�*���s���0?5�ES@=�;I�X��F�#%q���z��.�̲͗*�:������mT����&1*�k��>v��U��F%�\�1v��6�9=�q���� �Ǚ��+��!�s9"d1�e�Y���p��u�1g{@F��{t�/]�9���x�Ϲxo�.�v���d�TSV]7�4T���L%����~;d�������\�wPHp�?���݅jE�/|�����f��-�Y�(9���x�U�ῶt͎p��~
��`[m��UͼF�d$�:��v���$�2ws��j��~�=Ԡɳ���Buo�kf��Dor�=�U�7<(��O�-]F]�ZT�;Ǔ{��OK��P��q�K��x��5dKy�0�Z#VE�$�Iv�*�,Di�r녺����6�7O]}���<D�`�W�G���d�Y���� �ڸ�~D�JE�Z�i�D�~���w���mIܼG���?��I�95�95��^U.�ј�8�_9�*٬��3'�mpE�aXQ2~���Tq�hO6���p���J�n�����!牼���M��O���@[K��D\oa�j�����[kN���o���+��j��bz1���I��f�Q��AqS�TE���O�a��ͼ���������7����_���	Ǡ�#Yq7"�s=�@:��bbi�\$q�Xҷ����AC��k�-+mIXY�y-%=�ߙX���Q�W��	�8��/�g�/��9���#[��c��Y�S�ǋgY� |�����:8T����PA�@���"H�fC�D��Ǻ����Ηɣ���F&��ǐkH��Z7�߮E��)d���2��!�\7��?��
�P��@::<�"���y[] ��"%�(κ�P�����/.�~��0�2�t��F��.����uh���������W�̰c2�ak��t�4�pa3���?Xe8,�ڸ�}�u�MQe��E�H-J,B-C�w$UX�O���Q�?F�D9 l��"�hC>a$�H���2|��+;Q���Cd]���q�guMz�G�+^��o�N���M���e��~H��@\��͝aг�$��Cy�����o��H��W��Z�87)E���}�Ѧ�V��fI��,c���q�mY�$��]����[#�O<:��,w��y�2?����p#?4���Q:���g�e0�ôI���a7��\��5=���Zo�@ � \��[EA������u��[��Ȇ��4e�r��XjY�])��e#Gh��� ���_��q�-ԡfh˥(�:��3�����W/ C�H��+�]��E���������ѭl��X��j��Ç���P���`[��pk-�^�>��V�I1'�ߋ%����
0b��'�O!Hzx�@3��a1ɜ�.�aF�ת���;�9�g3Ĕ���)���h�F�兑���g�� .�X��P��+�F"�O�L_Hb�"�}�3H���g�]n?�ܤ< P�5���48��g�u����7c����n�{%����:�Ϝ����}�,703��?Y��HV�l B��T�D���U$��'��/<u��R����L4c��X�T4�$�=�p���5��`�v�!-ݡ�DN|�u������pJ'��~�� C�N%�LZ'� 4�s�\i��<�x͌K6g�ڈ�I4c��Hw�5q��A(z��YĮ���wh ��� bF����O⚗H�2&���h�,�T���64��R�X�0K����=����F|�%è��xD{6�7��t䨋�o�2�n�'^�WME~�0��yX�v��.v�.�_/�t8q��T��t�O{��<f��!:�d`R *���Y���$\�v�e��p>��(��h���#ϑE��<|�C�W��t}5^o兗��9�ڕ[�5޷���}҆mQ��^h"T}��8t9lvעj�W(O��C?ՊLE�DӠ ��#E�rq"^�m�>�*�sJ8XiS��N>elR:d@��U�=2��B����Y��S�sJ�91�Z�u��9E� �x����Zr�+R���o�i�AAn/_�>a0c0a�L��QF����]͑�@�O2Z0�F�����]S�˭�����7�"T���'�)��^����~����>�s}�>@�KiosH63��@Z�.���;�"�W�8Z�35����n�FI���UXM���Xٟh�WĶU{�r10�Z?�{|sƣno�q3" 7���?��4�A���)���!_%�IU�����(	w�N�D�a'Nb�K�W97�SXH�.⒳�-3皒� �8^`�m�)Ϭ5�Ӗ��k��8	�j�F[D�c?��uO`F��@Qe�%׿�fG�Ŏ(�rBA�uܼ.Y<��[Ct�~jF���Y[�F	]�W���W盆�)Uemf��l~焹n�:	GD�Ii~l����S���qa�)�w��,�ټ[�B�+����\�4ec���ۚ��K� �F{)�p��c�:���\3��̛� Ck8�`��Mt���%汢v���l4���A��0�sB �L�(/��h�����7�>{{�$]Z�D��00W�/�Km}��a06T���ł�B�bd��Q�аSw.�A#3_B_��Aߌ3��@:�]a��� �=�R4fZ�>��v|�q��\=��L*ԭ���+"���w���Y�xv�x�3ag�'��:��Y�R���6���#��t=�ī��� ��1(�_�y�����mW�9��s*���6�y���P��Dcj�� ��٣�V�?��e��~�� Cf�FFG� ���K7iWȨ�=o�j��L�kq��Dk�r� 
h��*�����]Ůj'�����kX/Y�qyor�~&	|�� o!jŇً?�6P�MA# ��렬X�d��Iw^a7���LP۪��p^������__�+l"�F+�~��]/�(C�7���+�8�oAt�.TS����a �z?�]�x�.F��{55����R �Z̶Q�~�Ɇ��xœW8������ڸ��>d�;�[8]�1G�e�7r߫zFv2�������^}�B�5����m�7���l���#߯���S!�w�d~�V����.�8J�6����R�xԚ{c�|6H��p��34P7��h��t��Wgw�r��
�m��-F�\��I��u��ςo�z$���%�x�"�V��ט�Nρ�/�E�	s^�؝��#`R���f�-��T��������d�(IW�3J���q�^�Æoy�"�=�+X���s�[b�z8J�:ڣw��Q��+�<N)�lJ(ٸ�R�p\=I�mH�T1�
9���S��t�{��t����[�T%��U΁C�(϶u�/��}�ګ���ل	Sgh�c��ߚ(��u
)�s��ue�3gN�&7���k	�:��\��E���t�T$��Fs3��Ϸ�WF_�qA��9�2����T�:u�>6��Od�}�)�nD�VoΓ�� �p��
�͒��9���k�,/�(T��,���
8�!���=k�[8�Y��?�����4�q�;2�����r��s��g��~'׽�~�"/ʿ[�od9
ɸ��Ө�[&�!v����6s��B���#�H�a���NY���O>2QY�4����x�S��sE5Y�'L�\c�_$h�,��jm�<���Eh�T*�j�h��ӏ2�j���<�w���c6V�c���?Rb����ۯ���~�F�c_u�����:�"�cu�{������f|���ۮ���Qڌe[��ąة�[أYWK���U�d8@�m�0�w��R���&حQ��U��x�;ˡ�J�c��g�L���;ur�ҍ���/���Zhoq��$�OhR�\��1�	�
Ye���n��J��5	v�C�f��.L#�}��pN{ڜT�S����R7��shM�0�����xgM���h�(����/������?f]J[���5-�����G�7w�ҩ�% �q��-,/���3��TA=%P͚F��b�]�����+�ê���-�4fIQm�5��$��D��dqk��r^b�O�Z�"F�>�d;N����c�>=��l�|[=$9��YA�a��N��UA��WxGw6��*�9 n�L�`9A���S>�������@�f�49l;0c��@�X�`�ؕ�F�'��y k��5*R��y��x����IQE����l�I�Z|�f���i7���tA.��%�M1�Տ�Ņw�)�n	R��ٓ{�Ȧ_#M�߬�?q���Yj�,��-�g�]qn>�<��l�0t�4g��J� �*kf��04К��RyI��I�ﷻnw��8MY�ݿD��)�h��y��]�����#
�.NE���Zl;�i�4��p��E$�D�W��H�������I��:�5���[�W���G�0A�f��?c�J8�7Cn �w6�t?i)u,'miF�_�Y�37}�w{6{���l��e���=�Vb]]�(�=5���� 4쓧,��,CwV)@����'B��5�oxX���L`& v���{q+�vF����<%��В�u�6dW�m�S{+7������K����V���&F5��STh�W�F-������R��1[�W��I_t|P��F�i���䮢��y��eE��A�5<���_����ј,?���!���ǌ�.�)�6�n{Ie�b�� t�i��D;W=��N��"N�.��2M����0��d�\�f�gj�B���2��4�M�-���fʄ.�:�7��*C����ձ�J��Qw,&�9DC��u���H� ��#�;	�s1��K	��+Z䜩_|�V�4��AQ��~T����IJ0]0�����V��q�Ǣ�f�+7#��Nz�WR$� aG�)�wKЦ/#�Y������e(�0O��
?���q����Y#\���"s,�������4.ܾ2w֌���iB1�{QI�h���-���B7�tY�tJ�O�˙��zf����3-φ��؛e�@�	�4's�/B�J����6��7$62����18�����)�2sxF�ȘI�nE ���"#�V������~&���- l"�)�/��	W�Хu����a
�T�m��#�p���%�p9r�D�%� �@g���jTur����V�T�2���-�̖��!۹rRk�:8��M>����i�I�Թ=�F��؏�q�g��r|��b?��N����~E߄��p��{��s����)��,�����v���a2��oڦ/K�q:�hW�O7�HQ�D��؍~<>;V#���s�u��[a�����I�#�ٯGB��,�y^�r�-:�s_^�m��m�(���P��|*s�e�L;�:�y��{�a*���/GcYt#ձ>z_R�&D�/��b��F1с�����{ٵxi&�D��JO�O�fGk�J`�x��c��tQ��IhĐ�݉�ZR��ß�d{Pu�_��.��hcFճ�y�Os,�@Ӝ���2��gzC���kMJ���HZ
,�X�I�h\}z���~�XwYe+	v8���pV�ܩ(� ��0.C%�����h�^��c ����d�� R��&�t����F:K��e�r���eh��e=���0�:�.�.31^sɀO�E�jB�������b|��3����V�w��T� 4�� �cE�;i��@��/*��T�bn�6�[B��ik�]�[��i��[�W,T5+��<(�"���˖L��5a���Ku��g�w��jn| ��ƒ���r� �^�����ٕ�`O/�,�%��2����JE�z��8��%OA0���p�����(nn��>����а��c�y����mR�T�glTt�W����˝�x�V�PfLM��MD�Q �QD$�&�&�ډ�3`����F�D�)���O'.�S��ZdSr�d3�L���-�v�J�@���t�4�.���J�(-Y��G�B��0͠9G6�����J�������t:܂���*�߭8!������xan��L�0����|wݐ��e-�1Gm@�7z�!Q?�-&�׽���< �9�?4�-��G��j�L\�7/^�4�' uX<(��[vAs6v������IG@�{�����;ռ]����u���.�P�Uݵ7�4")�c���n�?���ѿZ ��A��T�$�~(> ����)VManE.=bm�������g(�nf�t���!d��`�=�o��S��@O��ҋ��bV�ګq��f�$Ӊ���{d������\k'g�*��j:��듩�e�
;c�Zl��\2�ߪ�Ѯ��w*cFRwZ_�Ԥ��^�9���]ٜ[f�X����&�Yz�/��#���c݀��N2�M[/Wʋ�لw�5�8��	�ڪ;�{R�	پ��i<v�7w�w{��l�����6����w�8�nd��O���%[��BF>�ŉF�{8g�^ 7I�ǭ�	��9h�s/	�R�u)Y��!Ќ]����0
������0�Ő�{�}'��@�FM�I���&v�A�(Y�I݁l�2��L����>��ǰ- ���<D���X��7���i�P��rn�}��)��]I2��O����@K׬o��a��PR��	�O�<3�uV.&��m,н�I�+�CMZ��.�4[��� g,��j��!� �ɪ���\�8��$[K�8u�On: ��݃ǲd��HVL(�L���Z{�	7����-�=ϾB�@��w8�?+����ȲaZ�O)���V�����\�n��Yin�Ӵ:rC��!�!�l#��\�OD������l���q���f6�l�_KXONYʑ����MTy�D�0�n?�10AD���J89�������s!���.�B&�h�(�g����u�,��>n�+;VpP(�-_����.&�W�)6Y��D����v�tv7�#���(�$��'�=6͎m�R�8�ބ��q�q:,k)��j�Ϋ&Sk��i�Q�:"�AN�{��_�A怗#W��HJ��,̞`zx�Nb6�M��֪X�]��g뚁~lt3xŐt@�_�H�;Z`�ʔ�V�f����T�G!�F�Gr�7��U����g�Qz�4��qf�A6��zU���Ae�㙃C�<��M���DhO�)��ˁ4f�D��	�����Za7�gN�D��O�jz	V��Ɲ&t�s��lr8��?�+a�M��j������|�E���R�ߩ�N&Ӳ��J��A�6��D`R�oN�G{��1c3�u��	�	�>��O�٨:��F���%\혮7�<I��qj_4��-�!�Yp�=m!�X{o1�֐���vԩp�P�s?�����~vf��,c���K��yC4?��n$#EmS�_���9$6��r��t`C�,Ý,Tk��"�c�w�D�����ခGԛ�W
7���Wш����q��Ɂ�Ic�D�d���F��a�$�o�g��"�j�|��5��걏�����D��z�ΰ�������p�[B����dY����TA���m��D��;��u,���!�c�ݟ*�u�"�`^��!�����QK:E�ɇI�����f>��%��[�L+F���wq���ߴ�%*��:o�o����6��<�={�W�+z���p"d���Î�������]��`���Z�i�xV4�ˑ��_[����2���|7:�{l�q����v�n��o���C&?��Q�h >�&�E}̃�L	�FR3�Q�k�#c1f>U^��p��;n�39�b�۪1JD鈧5��t����d�iIQ+����	����?k�sp���"���A7��DQ ���)q�8��
��oM��Y��;�G1�%�QM�\�OJ"�s��B�'���t1��}�>�A["9yL7H�I)��AL�o��]I�N��t����߶� ����bAԫ��,�}�"�k�&��NT���W��|�"����� ��p�W�0��O�d�D��Q �L�} u�;ӧ�Z�9�ѵYp�t�)�Lx���x�{S
��|i}Z)�Q���'��c(�2�K����қ��e�S	.�f6�����o@����Q���0�"�1�,��R��6O�����[����NU@��e�iK���H�^�8��	�k{.㘭�b���jѦ,88sV[���U3az��Y7��h�'����?��(`��� %��ˢJ�4�γ���s���r	Tf͔�lz�S��}G��0$>O���Q=����#@�Q����ι�	�$��WF@9���*d8&	�E@Yu���¦�I(�P�+�sYH0G��Tvz߷�Z����\Y6a�s.�pэ 	P���ɫ�)�#7��a�՞���' ��\g��C�Tr��U$�̈d#Ȓi����M��j�
����k���b�����-��l��p*(G��>�j�|��`�������t��ު�A�|���W�����Hpe}�Κ��61�� Fe>����1&�D~�y��d}��`��ˆû�v׹%��B���A�R�:�XoK��yAN@{�1���~(5S��qY9�4W��fƤ�̫���.�b�>���I`�t���zU5ǎxuo�� D���M��>���}�`��V%�Y��ǧ$ ��l��z�(޺�Y�_q谧@ޡ�~��,��G��'���l�K',��tB5�ى�?L�,�~\g�N����� C�N�k��j{�:o�:���pq��1n_�,ZD��,�'�-Y�h�-��T��z�B"��i��N�PT�]p�MƩ�毎����!���
ri���ݰ'3o�tϰ�/L8���'yt�.J	ӵ11���������^��xJ�-��iv��.Z
e��+��
*���8P�C�Up��f����{5ʀ���9{��q3��Z� 0,��e;qU�W��ХW�٬�|�?�R��bاQI�r���K;��#�*��]F覫rݞM�+����4l6�|7(����g�� U9v$q��-	1�V(>'2%�$���m��,E��l}���զ��UO�O�ώ{��{Y��yi�r�B���ZP�6�CR7�B��������Ѻ�VT�r(SZ#���N�X����O�y6D��<�k9�7W?[�45�0�0e�9|`m�I{[������+�I̹�T��ӕ��|�&3�m���|��N��,�����=�πR�\�`����b�L�� Q�\^�\�9��_|E�:>ܿ>݊}&�����W�Aߠ	���V���z� �i�6��/I��}�T�w��;�
�FU x3�9�)ul�m���kŒo�@��ny>�H���5/�#�ҏ�~�k�u�?'�[{�Ăb\h���'P�4F��0V�#ىl\R/7�`��Z���[-K�<==��E��J,Ex4,v�И΂����,K��#�t�/�#�w����.-�ו�q�=�A��`d\�8�n�p�j\yV!���Ћ�}#iŹ!.Xt��gW1E0"#MއZW�[��Ts� ����"Q�*f����U��������uh�= ��	��	�}��m[����n%5��y[�J[�$<�r��@�#*�����B!|��L5��\G�r)�'���Ѝ*EΔ��<�)-�^ %�3��NEhڨ�	�Du�fN� ɞ�}�p�Yjl��>�h�z���9c���68�r��n�n����U[�u<�s4O�E���ɫ3�ȫ�s��ꡑ�!���R�l����\_N�q����(����\�W�m��z�������7.�8+���D�P{/��Y���ނb�{ ��Ǫi%iH�C��q��J�:��{E�U��\(��k�74��J���oN��f��z��+?!G���;�������!M�ֶn"L�M�;%��>�7��SB�o ���Ө��"+���������t*��|z��"��c�&]�~l(�?5,pm!�J;f^�䭽ק���i��K��A����F�|x���I�x��&ؽ5��(�kx���zX��IR#G��m�¬D�t'^8�������������k6���b����O�tq���s|��C�B���.�[��)�������5������d�xΦN�'|h�u��&��������'��^V��e��7	9��wՊ�E�gT�G0~���GYdg 恹�!4"��.��j����X���
�}m��B������_S��~�,͗jA, ��޸Ɠ��M����ò�V#��$��뫃z�Bf|Y;�����;�G�@�c{���� T���)�0�L�1v>�E�tlC�����_~URlk�}$J�����m�~Y'�k�ʣ�����Q&�7��
�����bm�I�-�֔JmѠ-���&uҷL��/����\�|T����3�K �CZ����J�B�.�����2	t�rK۬��uv�<��$�6K1�/w��u U�[���N���cv>=yL����q�Ҧ�#��Nh�!�� W�^��bX�СF>��Ut�"v@�ە�S#ї�E'ރ�,�����z���>B��J?ũ|��%�'��y�N6�-��1�����ׯ����'��%Q����XϽJ����ڒ��6����ͽ��q�ݎ��H���д� S	#[5�;���T�1�$�v[h�	�)%�쏹N���R�5;���2�0�X��^M`�R5�ļY����j��$勀���x�^�ߴOGɒ�
'���Q*�VN��1*!�ʡ���*Je��Ӛ��(��ȟ"ǹe�r{`^$�^��T��4�3V����{ՄW�C�K꼦7���v�Z����Ȓ[D�6o^� �I�H�Bw����ޔf�D�	%��'���"as���Y>����=I�DW�8���HG��Y���� X1�+�]>�#����E�<)�t�I�/�s�;K���|��#����ܵ�o�4�[I�_�%��վ�a�Dr���3VػC�D����^����N����/�P}p� ���](۳R?�_@�h���ZJ�ё��RY3��;��0N��2b��4���=8s�����(�� wJ����J	�sz5��Q.5����]WF��B}�ߘH�@wľ��g�� ����Q�X_"�]ֹ����
���,�uD�։]��d���f������T��i.b��;�`���i� .�yOZ�aI[B��4����P;c���X����01�LG�>Uyp�l��3�c�D�Xa#�}�ߟ��;[���%��၁�]<鿋��֑�3�y�ǹ�r��yj��%�`�i{0����R�'˝�r�z%b��������(6��V�t����1E�&l"%�Y���l	)w��������@aK�\F��Q�~K�Uo��U�Y捍��,���K�Q�:
8b���S$\
���M�u���8�~r�E���d$��SO_ ���<}�NpE}���>�c���g�����X�HА~t;�we݈�sކ�"\�T�L�����q(��G� ���%?#�J`F	*�a۾h����,�ē��;e�ӽÞ�^f|ى�sЙ
{豕�3nzv,��^�	���A�Z�����Lʗ�>�j���3 ?���IA�W$��
�#����=-`O=BY��8Y�hb��Sf�
22sV՛���M�-�#Z�V���P��"k'�C��G��F�12�w��wU\���-$?���(�ffShw��Bp��ơ����Lp�#�8�Ҽ�PbV'�d�����|p\�ÿ���)}�M�O�ʁ�y�{2��;�F^�U>㓱����2�w�5���{B��CO1�nտ_ʋ�XУ�sS����y�b\�}&*l�"Ѧ>q��7٦G2� Jgj=Nq��8BИh�Z�=ll��&��gX�i�*P��2�<�E/BlO|4̞�J�q��Z֤�8@��P"�mj)_��jN�:\x'*��Ù�R)Ya�o���u�+j��h�7/U��w��.����V�P��2DgS)�������?�l��w��/�&����u�}(�8tpU���,�,��l��;;!�"8�j��7���tⱵQ���͍����I��Ҳ%�|��&n`a�ގba�F?#�D�XJ^9�q�+Դ��2��á�5��"Nٸ��=:n�u:����ZϠ��(�մ�m��AqD��r_[�}�r,?��l�&��:�Lc��Q �U�J����jry���.A�F��Ȩ����~t���D�wsu������l��,o�X%%AcU9<�+��ٙs�p�(3�J�r2M��ײ.֤�l����S`M��2�M�rC&�պ5ZDW�I=���WM��dާM�;��ɊOX嵌u�tꤧ 
n�I�����_V�I&=U~��,����1j�:�,�fo�zԇz�n��d�ê�&G���G.���d��6��X��Z��3���@��*�e����5i���^���Q.�S�a����noޝ%;'&1<"�M�w�u�H4&kW��4(�_|=7�1gN�֤��ag�E�X2���SY~
c�W�h/�}�AČ�hxRc/UH5����w�x��@�z�f����xa�K8�St��#}	F�W~+����Ł6Oq�{E�D7^@�i�un����[},�<	R����`�k5�5�)�(w��D���E:�H��O��o$�!�vX�g��
��|;�4G���H�{t��n;l�kIP�n��X���01�����5T��/���eڰ�P��|��-Pb@z���=���j,��Z݀4�V'��O����׷��g3+�*d)"S�y\Nd�I�	�>7������~�kukCg�/4-G��5��({��������Z��`rަ9]�[�ЙVi�\^jڵ������=g,L�l�x����HlF*��(�h�e��f�i82g2��)P�(X�U=��o�<N�:�4.nXI|2����+�(s�u>��"!es�Nis�ک�9����z!����{ٙ$ CH��,�M�p�ʒ$ V�h2K��߮0CA
�e���RA�Y8\�(���t9⊗�ۖ��� k=��B���P6�#�U��"� .��M��Cbc �i.���ĭqn�ý��b�'I�mmdB��B���}���iƀ�NVF+1�Ŗ�݌K�"��[s�"��9�����y�t(	F�sBј���|�ϴ#$��,��/Y��_����ص{Y���z��'��WNQ����1j]�M�J��"��:����`?�:�^��TDp�e�Y�u�����
n�Ӡ��C�H1��@e]A=uJ�{�M�P�?c��z]�F��I!v!X���]bSq�W3��h�L�� ��  ����l�D��%΀���a62�.���؄�.꿚�#hC���h|�*i��d&�~6���h��P������k�m�_<�_!D`����~p�՚^��ō�
���bԗ�5!��F`|�������ļ������ډ��T
:��	�\o�������(Z����F�$+	@(�O�*�ЍO�KP�fm����l��4z�3Ԑ�������S�{aoGB� ���X�K�@;�B��/�k�­&6r����X�H�"���Z
ik�{�v���MQAL���xￛ�+K��P�}tM�dUh�ԙ�Ty�5���Y��^S�I�>�TD�	iԙ���0/" ν�����K����0��֕��{�GpZ �E_Ne���檘\�	�nH�8՟r����u�Mh�Z}� �M\ C��:��{�A*ַ���Hurm�A�c�q�t��R;�����
���6��9%˳��$�`��c3Be���m�_U�PW��]�|��|2J��L���73�O����5���;�i������yH>6Mw��ǲ��X6���t��W���ω� �ց(�̝�SO`�\�p��i��à��R|0+6(�
#v��i$��Qj����;��E ��$�P�R?N�|fav;x�뿍�������J�J芖�D@��hQ�w%_���C0��<.ћcOg�b�}I�9T$÷\@e��'�f����/�YM��?�<1\ά�1��u���؆�a�\���(�,/6����9����z~eR�W�{�5�	%7b�y]�4��莩>3�=�ڜ_�-�$
�'��j��!�8�\�����h�����v jkt����`Bv�"v�tc�|����t�S>��Z��])N=�3�q����:h���V��F��.eG'�u���Ud��� �L�Tڶ-�G�ٞ��O�m�'K sx���9����˳�����j�{i����!��1�i��1ŏT�׆��`;���^Z�χ{��(;H��F4��sF��ݔ10.4�݇#]�&h�d5�蔲o6��7&�M�T4-c�01�5��>����c��	G"��8iƲ���� {]U�ѧ����ce�J�Ť7���aߎ�Z��$�F�g��PT�<uLHs�_�Yh8��"�f��v�|5M]aXtņ*o���~��5�%���O:&o�༢�]�(���Z��J �8���W0�.��V�x}@(�JK�0�9�E��@ؖ���ח�-v��G���1�2T\��"������E���Gǳ&�&�L@�����T���	�9�qڛ-�-/�)e���chp�ݗ�q9<f�<=Yv��j����lv�x���ӆ�g3`&�=�	�L���r�sC`5Y�F���m��o�/�{o%!�˯�򵸉���$"�g_���D+s�ɒ�J6�;K��d�g@�Ķ��I��r���WE+ܳ�:NdÌz)�Q�"[
�5'A�kOhr,y4o.p��+�����o�j"�Y����Ƞ"F5�ݨ��hm��0)��ymJ����&�^���#��^�k�s�X�8�@�B��2��(<f�a���O�
�D~ (��&��A�?����nJ1�Ō((�+� ��k6
��W5,'�1ł��2�
,Q97��v�Sї�$Ab/6'�xiz6�I��e��I�U.���{�H�A�����<��7�#h�,��P�g�����:5i�0�sQ��8�UgcP��Y��.%�����V����V�`F�Y
�}�����B��4��.08hT�L�rvƵ��0[��dUP�.4f~���m�u�a~�P.��_j��\����i+� %c���?(@�EU��R"'=BJ�V=�!#UF7aF�V�^Ѽ�N���פ���as �U�	�Ex>)���<y%�Y� ��Q���9��ޢj��%
�b��������Qo��K�*]��V���W�G��v7���,�q�oVr��1���*�A����JlUZ��N�׳��A�c^c�4�3뮛<`�|�QAz�J��DD����1KK���0���9����� �T��č����%�l
����
�����0����i{���G3yXٹ*=gC��dՓ���q�����j�b��Z1��K�}eV�ɀ���:��������ەU�P*��v�"�`J�ɓ��<޻Kהvi+HJI�n�TTo`:`g:�=�h1����&�����*�.N8b�@2�[=�C6�ԯ�0�Us�^�g������.��<�Xd;gÜc��m��QBp��-���\_�.����k��v1G�ĕ����/n@��8�p�_�|�BQ\�+9t��};&w����+v'���6�V4U\�rp3�61��4�v���T���K? f^�������eO�=��]��Y*_�V��9�7���
}k�*f#�0�J�bJ��Kų<ݻj/�F�C���Oci����9P�ᰢ����[«j���S@]*}� p��G��D��J��X!����p��"Z��j�Ӻ�2~��+F{�j̫���i�5�,����%O��A��EC��w�A�3	�a�!؅��)����jl���^�p�0�!��1��`u�;�^���OHZ�#e�z��Q���6o��8\�;>�+湺u͹Z1!����8�,撑�Y���ڧ����\<�{�B�ު�1G޺�'�`k��SaVծH����� �@.�A�C�p(k�UvL��_���
����fT�$G�"��zC,I/6ef�n^>}���mu�䠫q��,ec�<Wa���]-
?�?�fc5gOl_�z�K���,��I�\�I��!-;U}o�0�JuЩ?lBt�k2�A�5_=>2�W��tXi=KA]+��j����*�f����g(�?��}�ې!3z��͞����A��!5���
��9թ�;�R��y�%j�m���8XP]��.�p[<i�<N��NG����!��_�d����~�g�Gb�m����y6`Wp,5����v��CK���q�@��M�ݪ:,�u�s�q�ATG��i8���dw|OW�^J�)��Tz)	�@D7$;�
��,P���*K�.�,���`}�B�փ��������9�� 6�:Ԟ��>wo�ONq���a���[��԰1�~��I�M��Q�b�
��Ij�jS�8�C,�o�J����Y8=oõ�tw:NZ*$x�X,����l��s�7����rxԎ3'�²9u�]�ߍ�92��g��q�@Bs��A~Y�FKŇ�� �=ݟ<�3�-t@PpM5�m;ؙu4rL���8H�.8�Qͺ g�Nq�࢈�g�Q��w�m��O9l!C��Y���p� �Ͱ?��|Ⱦ�#e/c�� ���-�b�WG(w^4B�0���L��>�N��Q��c�� P�H�A�Whi��`9�8Ivh��y�Ұ��9�}eh��9���Y�}�Dt���Z`��-�+�-�K���ٮ��/G[���$�gE0� Г�r�'�׆��ED���.V�����6��}�@A�_�(N��}Q�[���D8���4�o�HĈ���P��l۾�8�%��5��ы"@��aYÂ�G�!�lD�L^���(g�g寮R�ps dlwL���<�E

�4}A��}�.N�����>�G��Fò�����*|�-��ټvX�S���!X�"*(�VYؗ`ܠ���6f�o������+`���=T�3�l�u�?�}�޷�y�#�-��g�Y��m�^��7@9>zoj�n�h����V54H���
�BQ���y*0�Ƃ���M��&��f����b�ڂ�~�)���f���.��6���گ����(���t���B�5^'+]��}O��h� B�O['j��֢7OH|��>�����n5x~;o���� �͡��&ou�x��u���"�����MOs��ھ���9EX!������T�?�NA��n�t��T#���Bqm1�?��Rk�>�3�:��Wpg�=��R���A^��1ڨ��:��V���{f)��<!)sO�����<�K��&�	Jܙ��v�Ӛ���6EoN=�I��]ŉ��
>��2���4߂�p8��� &��ir��=�*Ƥ�60l:��R�Ԁ�e_Pؼ�QE�*��f18�}�ڂ.Φ�9�_�=Thf�f�;4�|��S�h����5���T����,v��?Mt��>�u�K���h&W��`�7V �N���+��fq�㒲�D�K�X��s@{�u!-'�jM�ؽ�,=i�U:��'e�x�*�g���ljP��I[����-�p3��o�=�F�@SVީ8n]("��5�r=�@��>c��?����p>5Ғ�f���3H6-���&Im�(�+�	�t}�C� ���p��Ѐ*#�wp�eb�4�+��؊���ղ'l�7�8 3����Շj梭lӶI7o�Io9��b�ݍ:��[���:"~Q���Z!�MHmB����z��\M���	E}#]���iU���'�]?�`CÂ�� K��8���k�z�՚{$���w'X����K�5(�dk�9D�~L���M�8�l�M卤�RI=G#&j��=��YYZ"̠1Zu,b6��N�N���b/X�&��U_B��}K�*o$H %���0'��R�Bo<��r;
/[N�S$��,1d�멡���Jr�u>�̶�;������Ex��چ��Km���SH�I���)��R���7��h+�=���v'����f�����^�	�m�Ư��|�����_��h�G�����e�c��N��r�)�h��Z�0"pR�i��]�B��ÊO;�j�8$�}븶'UR�s�|�ܴ��d����[�Ke��n��	r���63���X����N�OڈO�n����C�v���֝Bq�Z�*����,G�{'r$%}�v��5�+���f�;�B�N+@g����_
s�|
��qT�q�ޱz9�Y9#ݚ��۸$I^�l���<5(WL����n�_�v��s����2%m{=W�'r�'�|9�n�㰔ܹ�,XxG1
ܖ�����	R~~�m`x=�w�o7~�3��{fI�A���%_Ʋ����Y-�� ��#�O]�өX9� ߙ��<����_�٠\w|%��"_j�4�h� �n7ԵMM�u�]31,��[�H-W�SS}	�l�0�8�eI�V�j�M���خ���̎���z���!a���_W7�A�A`�SP��Q�{_-�s	Т��C�qRE�g�ǣ��!F<��7�
���̋A�B�޺�1E��L�$gQvk���^���P�%e'������&&����J��m��V�M�j���!ݗgQ]�`���O�+���7@�ȅ,��ɠ�o�?�M�jj�x�w��ОO
�1B]����])��w��%R��H:�"�|��y��e+j�����0^G�1\2��=�Խ���'S~�Rlʮ���sk�[��D��(��Z��J#Xn�Z���?�S�u�E�@օ���7���]V���+J�+d����8��s�{�6�Vɫj�0 &w� �Ԝ�t�����Å���-��l'0W�5����RAr�0b��DF�ީ��<h1��zƒue�Y�?�F�.}�)(
��?�iڠ�I��S&l J����
�}�����ݼ^k�E�	�s������QS�w�8��<KT�ZqB���y�t\�J�!���׃@�]���*_;���K0��k@m�wOx�16��͂0�A5Q�F���9f14Ұ� �8��4���yvO9�R�EL�1�ӺLO�7����(Gm��Á3�2�X1���{�	 �K"!O�r�|�w{�0�K������ĭ/�T���TY���R��%8$.SM�n�Z�����J�X*E��0q�S3�v����Q�ֽ`23f��P���gĊONY޷W�r���btL�2S��[m���٫{�P�7���B�S�L��,��`�]AoJD�����y�q�~5ل�wD�m#���Z�@�$�qH&��D�$����eu�w�|D�iòʯ��.���n�Zm�7��R^�[���8e���6��B�0�u[�������aA�Y���Ǹ����3k �''BM�	��3���(���p�T`��Y�":*�ꓳk׫#(m@heE\l/%-͚��a/��ሙOo���h�C�`Hܑm �Kͭ��o��ْ52�3���i��d��u��#γ����z�6�f���¦�?[��r��lC��C�g��Z�v�E,[�Տ�\��H�o�h��U-ϘE<X�R\/ �7������Sg��� 57��y]��2Ը>�x�Gu�
y?��*֞!k�S�%w�<H�[��X���~_d��J����\f������7�$�0��Ytx	�H����Y��F]|�O�ƺ4�+��A����kwx��1i!?Z��o��ѳT��:$�Ϫi��BL%U��]�a��^�g�1��a�1m���6o2��R+����P��N��k��mP��Ǹe��V��t�C�4�nȨ�hD�:D���:�B�S�~O���.G_X�ϠY�edP3�������3�0�Y�V�@�.?}晋[�^q2܋���j����_4��A���&U�E	�ѿ�B��L�00�ᩆ�T�8�jg��(E�@ v��5q��kw��e�o�_�sć;w:�Rg>넧A*4\6�XIO��D��3"��N?��Nx�|�w���c�&�E���%H�s��{��`�uE�:~�K���#��ڀ��5צh�
�3����խ��y��Ԩ��5᣷���~�1��ݟӦ��1k!��K��>O�Vĸ��������<h6C�O�coq���BQ���	��c�y_�6YV��,�C�I=�m�p}�d���H��H�����}ĉ��M_=��em$mP�oS^q~o��k���r��yH���+�੉{ 1���wz@�^:Ȟ�'��4ܧ��/,��,	��ml����Uc�� �����S�D8�g>E�j��5y9z �LQ!P��|Cܔ"i�*�t������#CС�N��x��+�� �OB��w���=(?mCN���/��|Gi���Ց�w9c�����Oƈ�Y�����}�JZ���A+L�Hh��4��ܴ壄(�,����WY�1U:�μ$n�^@ʞ�Ա�d��5'aM�V:�ÐX4������F7w�E�_J"[�s�u��e�<l�����Ę��k2�ơXOM�ژl�d]���Ќ5o�����}�י�&l��Ыr'_֮�AQʊ���H%��q�,LlT�M�GJ:��<u�L\����W��#���ɔ���F쫻��D���}b�d�*^�\�����҄33�v�������aL�s�2b�<zG$��IH�Z�+d;�ST^�\�_fՇT�n�����<�݊3��m����g�MR��őM=��szTn���a�R��;�2���ܠ$C#�j� W�)���BtOb��oz�|�b+T�15f�dF�������	w�7ш��iv�)�4���7E�aa���.,'�1y:�;����B���#b�c����A��&3ژWߤ�¡6sA"�y{�E9�8�
�ç��_	��D�(�V���Z����UI�>�oQE�zƬA�y<u2�K���ߔ��`��s���tF�}�=�uLB�n�L�.��t�s�;Ұ �r��m�ħ��暄aܞ�-�0)��m>���\�@*�%�qEƝ��Rs@h�,����X���E�:\�@�}��K��箣�*pTʬ1�P��u(�Yd^#]��7����p�j�.��)"�Ρ�y2^l
Nd��IZX��xA��d<����ME�#"5A����C�����/�kvcrxݛ�����f���"�ϾVe��B���p��|�
~��L��𼝱�����Gu$��QM�k�n��<(rhj�,��B��B89�p6E��2{ �)�VP�ӆְ��o��9�����~Fj�}жypO;��z.�^('G���e�����:�+t_ԫBk���{r�Η��Eob�8񓪻4�����}��_���q����<�v�b�cm��+��P�5:P~��ᅊ-G��I4��f�7S�_� nz�qq�
 3�ڸ��	iX�7u���o�L�f�S[�1�}&�����5�"oEKJ�Eo���$�Z鮏70�������f�j����8so��b\�c�L��ǽ�,�Ah�����]��4�\y��,�D8D2~��}��4��0��;��$������G,�JP�Y"���pt�VI���`��z�-F�D8g(��(�F O���H��g���)L�.v��Ó���fRG:y�^�_�I��C=^R= ���^�`������8��&��6�� ��ޑ�V����QPi9RM o	Z� ����O��V�PX���A'J!�8�p�7��W0�������]�*��>���S��nP���zU�R�?ײL�pCƆǡǓ:�W�� !��MM�Q�{32�~VGC��4�X�C����y������W�AM��O�:�0A)C���/�zm��c�S�v��n�)*!����Htnd@���$ؙ��2��5&����X*bad'�|�� ��ƺ���V�u��ԑ�gx_����3��e? � �4��<�O\��o��R�g#��X�����i�u�\>�gϣ9�4h�Z�"��&��AK����!6\�|bf
���/��&b�gס
��%»�t����nx��v��T���n�<�<��\�ݧb+��������l@g�k�_@��=����M�{��U~�X�����'l�G���Af ȋ3�}K�1�wo�]9�"�W�Wv�u�v���Ī�ͅK��O>�N��YP!9 \V�Zg��Q�PY�;�#ӫ|�u��x'�>Wn��%��]��巋!A,t��:^:�<�Qrs �y3��p�f1�o��@�s{�2�^\�.�����m�@�����M"��^¨ݥ)��� ��+��F:n	݋|��JDc)6��ob�O�,�q�t���e��Fx(vg���\�>���@���s�!�ħ̈́����֓Uny\H�n��E::lls\�!2)M:�L�%�}��g�ux��-����he��xB����'m����!b�n�h��6�]I�Iwv$��$��9�Ԍ��JP+3�&�Y�LXl���}��ũ_�N��� 是��|�'x��Y��Ux|ᰮeS�S5)-���q>��G D�4s���W�։bS����O6�q{��P��	�tIV������EC?��3'������aC�ȑc��,.ޘ]�
���;J�E�	��t.)�;4�G<@L�H��4>*�g��f�t����;��Q<�$���$�E�k���n�����}�a��?�_>yMk�7�,.�����}^� �}J�	ֆ,��(9�5����B�٭�K!U4p�k����l�HAi�ӡ�Ru�SZ���?0ck��9w\�+�͌���<�U4�Y��ZK�R���L%&|�ˤ�֏X0�05oaF�1��r[�P�����GFao����5�����l3ˈЀ�L�Vĥ��"���s�vo�%�J�K�I��
� �.�4��,]�M�	��P�����o�"�#��2.#:X��S�����-��\j���F>�u�C��&sUxZ���)|Dm�E�ޯ���Qv�U���K��t�tThy��|�F]�>ei �zE,RuC�� >Y\37�������@�A� v���������
�T�'⦐q��X�GqyN2�mO�etW�rSƳDj����Thد�[W#�*v���MϱK����p;}O��V0�D@�i)�È�⻋@�cV��Z%X�>+K�Ц���[H(�it��c��~?�5��
N�n���<���Jg��._�|��Wɨr���Kpz*�h#��Л�m]su��������<��2|m�x/`��޿�����YQú�Z��fΟ�A��C�Ds��t�MM��o]JԀ��,���ءQJ�0&!Gj�0}�xii)9��^��j&7�5�p�w�r�&mXF�V<�%����GϷ�^ȥ��j��r*�vB&m�hDZ&CM42:M���4q./��䛏ga�6�`;�ōY<1�5��O��|M�JG�����	jLt�8�w�7�v���N-&�O�9֝wuOU���K )ߡ	x�*S���XI1/D>P���ݛ��XNK���Iz��E2�>O��Ig��D�_��B��� ?r���L�2�Hؔ�b�4��<�tZL)Et�S��~����r�d8I ��N'ݻvږ�us#!�u/mK`�)�^X�+���S[HB��W�AV�OV.��H���՞y?��bv��ِ������"��������P�J6�{�����2���a2
�����nl�
���ǩ���P����2SK)J@L���6XS��tA!k�hn�w�=?Z�nJ@�@H\f���p��^Yf68��������	'��&�J�G��W��
�%�o�&Ⱦ�:�� ����{�4pQ��v�?&8�?n����/'6QJS�����T^_tk��6ٗ�O`���!���_c�K���q�$d��|�9+�d��MCe3����C���Ч� CiAE��=��#j�Rh���5�v��=A�H*L��|����J��0�4G?�a���җ�!�+�v����	��
�J(eתz�Jq�ؔpP\����M�����3t Yx�:?A.�.���Nh�-"|A���a�KO�J8�@�Ċ �h�g�ڛ_F�����2�Lz�(�jFo�,����=�,�,i�
'p��3�ܬ3:f:o���Wh:���#�lF��g�D^D4�d�+\�{'fBW��S���z��y� iPb�d��I�V�K_�+kD�Ѱ�>I!?��sݷcB�56a�t$$.d�tQ1GF������_���Kc�dh����ԿNDq�~@�^�ƴ��0�/� x�,�MSz�]w�U��Ņ��51��)��R���q���[% �}�*:�s�&�5�׀�}�����Iإ�Ԥ|s�fI4Q,�O���-,~�לM@"�Ƽ��\�鐛R$���RY��[n��'��_�_6]B#�
��A�k�<1"�A��PJ:���w��%N��3=).���os�]��fe�x�NR��*/>��HJ�WYGQ}i.IcN���QWd��w���q�J�ʦ<��U�(�?�a`l��4m8%T�6�gw�r�d�y =�;?�)��t���(���Û@�w��(P��L�����C ��U'D�;�ܰGsJ��D����w��@�}N`+G���$�x��rL�*ܔקH�f�<�^㻀�s�� ;sV2����.��:���u]�.�?"�|��D](����1;v��.�[�a6�0�m ��~��7-����{�������k��BG���QFKq�P��g��/�e��j�����d/y� �Y���W�D�o5|�;���pTٍ����(���@�+��a_��Ǽ|W5 eh�Qw���U�N�X#�(f��M���v��|q*nv0�����p�C/����W	�ٝ�E�A���;���(rz�U9A�0%��}z�dԆ���XS�����k˭�)4�H�U�nۺ;Iޛ��-]�,EUd"@�"��2a��C�"iY���Aߵ#���.?K�X�o��;H�'���W]�'�S�fE�.����H���^��(�m����dMV�o؝f�.�bJ>?����%�}�!�gpO%�IiG����ť�e��u����)~��jjgj魔E�i���n��iz0����9�0�p�9'�W��U�s"���Dj����=H�V=Vr/@�O��ɭ2�]g0ͥ�}��8��~�ITo���P��0BR�����Hd�œ1�iSF|���T�&��2:���#����]1;�����y*Z/���q\���*0z�d��S�*�ْT��2e�o�Bɇ��E�]�2A��dEZ=��;�B�"�$���X7U��d6^{LV�܄8d
�Ǜ�h�Q/)#
 }�`V�`a�Ҽ��0m����@�� ފ�K����&b��ȍ��2��:6�U7n���c`5����Di�Hv��;�U:r��[���He�3��p�b�2&�-�lA���rs���5�����L8�3N��:�F�%�YN�"�8�@��Ӏ��JaEc�,�GH���&4L��q`.Wɽ4Oa������G�/}8��<H��&ߜ�(0��k��k�f�\HJ���úzoG��g͏5⢕�et#��Ҩ�p�6�e5xY��G��i��6J�gգ7*��c�KDZ�:�T���A�(W�Ѥȹ�`��甚xLN����(���8BQ�.
cƶ���R~�N���!�/;��)ܹ����Bw��k��a_��
�#����+Ν��z!���$8X%�����M��O�����y%�l.����A��K�'��ܷ�V8͹�=O���\Z@�퍮հ����Yeƍ������ �����o�=�Hm��%��mK?"*�kB,��O��/�3<!`�rU�俕Ј+o�����3�,���Rz�+�k���Q`��8\��i<���c�ӽ��ڴKH���A��G���,�
��G����%�=�&�P��H#�c�%4�?*qf7���\�� e�?�ԭXC�ܫ4���>0{̋�_�ꅚ�i���@Q�P���\�R�c�<�i�\�Z����Jݧ�i�>H�2��WO�Y��kv��U�I9wW�N��t�k�=�Z�Gs�`�s>b ��r?�jGI��o�x9!��dT�E�#�O`)?ݝ�=�~sFX�ۘlF쨹���{u�S|<`�w+yCꂣHZ7ID:<�����^Y�e�/��	���x
�y�����C�瀥?��>�NR��$2;帯�x�5�:���jM��u�R�atF�0hF�O�5��|�a �VT����'I0�f�{����/s����'��I�6���Ӣ̈p!���W.�Nx��'��`���Kyw���;�k�X���&�$+�ex1c�:�:nէ������EW
d!�9ތ��y�-&�䩒�PS���EsEY[a�N}'}l��0O?�F��5s�k'�d&2j+"�$��v��_����Mљ��3���J2�obCY��Hl�[���݆6{���\"��u%DN�=נo��,c:`p��׾J�j�eF�/(z�<�w�F ٍ�=�ن��=&`o<�d�3�&�":�����2Hq�{S�|Y=�%�ھn�沇찢-Z ����̥��A��G���#�/rjsd����]��s�q�e5i�-��� \��O��ӭ�M��x"'Z�L�g��'�ݔ��p��{���T����] Ӑ}����O�xƧ�ʨ�N�t��mTm�ОZ:�u��ƪ��<���ŤU�&��6��v������и ��'_�z���d���+���g?��Q��R�W�Hp�����7��V X}̣�p�i:U�A���e��\���~��r6�:��C����8�XG�/����jCä��þ�/*!��z��p�I�O�A_����C�@�{��">��e��wr�j�+�!�&7`	������ዦY��C�힃����W(��9mf��Q�#�+@����ܶ}V\'rP޶t����(k�1�e����(U����0v���S���Z��(��z�>�j��-�
��?��,��S����5�^�%h9R`�Ҁ�W�,�O۲y���*�_ K�'kF�<Y��!�U�L�d	�Ī��mm��eٛD���0@����J�D��LM�{��f�ĸ.��	�:p��ys��Y`�;�T����c�J��������4a�g�7{A���������B��Hg�E��	���(k�[��(K��W/ͭ�O׊~/jհNR��6$C�D�l�ͣ��B-�\��=��7��	,�0kց+/��:/�U΁�Ad0���,d�b�T�����G+�-�~E6�$�_+��/8��kFjIv�#1b���w�Oۗ#�]���Ƅ��h�� ��A�:�Ģ��u�_�����P����̓�H3����v2��6�����?a�ʇ2?$� [����	 �� �=�1ԬzG�C��:��D��-��TlF�Rej���eVhF?ru��	�"D�a:n1��O���ٹ���LF� ėovpp3�x3��K[($r���F�8���X����п���ϱ�p�+oj��nޖ&�v��*^Cֲ/��6�M5	[��/!9V�	�:g��R��D��+�R�"=I��8��.��V8�e�y�s��^@��{ai�k?u�D��s9�;�p@�����	�?xx���pt̴��3���+/�JǼK�k��L�bܒ�����:�U��1�Bя�p���~����v~��(�Bf��R���d(���%����۽3S7���o�HY�v@����)�3����S;+i짔8�C%E��&��]��4�4t2��By�UGJ��;�p+����d�x9������b�L�&/Bhɶ�u��[�1 ;!�.�޴�$����D|���2Sr�@s
��r�Gu�^q��B�O�u��1s9��=��Z�D������\ d���VfX��C�Z�'z�r�s*�~���z���;���
.2E��t���D�Eu�!����&E��H|��2�����V��2w�?��=ʨ۸݇*o�F	��P�m�]q�� w@tqOc��եcbu�˱���P�v,��k88ba�]]2��T�	aa�J�D˕�Q�?J�)�|��	���X�f�&��&���W��G4��+:v�_������ƒwK����^ܸa�z7�X]+���&�1�����]��8*$��+��`����nܾ[�46�����z�J5�>i7/�h>g�-�D>4�����]���KR��O��P��w]�=��q\�fN���u���;3��$�u�:�/�̄���˟����	E۟^E��|v����tq����K+�-����mQ�O��7�􃖕5��Q�y;���8�;D�h�M�6d�	�ZUy0�/'�i {s�����d2T���T\��@�q�c����C$'��e�Ҕ�C��fj1�����6o�����GLta�w(�C�Sykq�H=���B:K��ː$N��_�t�]������h!K̺6�9W�m��!�xk��↬���	���q��?���{�=����J�\3R3k�G�o��n{��Do���o���&(�#�(�߂���o3K^[O3@��u�=V|�+���Fz�)�,?.+K	/�N��h���l�fX*P�m1��+�V6���r���h�}�4�J[96v�-7�������j�����[<�画�aD��N�N����EnO��	��]��c�-�w���_�����82�Xv������e!�X]���H~�SF�6��UN�"W�*zb9�)m��N���ңc
a�Oi"[��k�ݛ��Z��~��Ddl��+p(��B��:�t��,f��S�~���)R�,�m�e����� �%�M&u���W�ֻɴ*w��I�4�n��/2R��°8xd�FP�U�t;n��z�P{�ٕ���d�%w!j��NL�%Qcy>Y+�d�V�����g��r������6���L�o�G��U�t�6��� �����>6rC[���Z�}$���,ژݱ=ˍ���ˆ���r�.b�t�H���	�D=@����� �\��(qj^9=���kq|t&��=�"R;)�T���hv�Q�P-���ƣa��5\�N݋>[Aj`��༏��r�k�O�a
�+�Қ�&ăC����-��z�\�T��s���m5$>�[訜	G��-i�"�KҰB��h�"��NeCn���s�?z*4r�b�w-�V�X]uk[�#��VA�(������jO�q�@_�v�ݶU���$O`&���nvn(�ep�æ����(�}�؀W�o�(.�m��J��J�=G���Kf�^?Xz����W�Rl�f��z���J�?G����D*����T�Q����=��s�-w�"$[�ZIA��-7���c<t���)M�s��z�X�܇��+�����f3vI���
�Mۂ&!�E����^�Z�?!?�gʃU6$��6�"z{X~M��̷4��HvK,��ؒ�)�Dd�_�,�n�%7���\�.�y�;�*��0�e�SYI0^�p��\z�E��k1������w겾52@���j�!Jӿ�	O�مG`j��\��HpR�=�`���1���	c���/'	\a���y�0��ÖZ���?a�}o��#��y�f������\�e��QZ�3��⹃ޥ�X��Jh��fr��^&�OǼD�<����SN�?RVU��K1�j �P��V���Q;��D��-�机TE]�)k{C@m����T!���J�B��i��;�B�*��I��jL�Nr���4R��GX��z/�s;a�B�ړ��Q;�L����N3�yy(�m������T�P	>K	�i����C���"	ӆ�d��;��S*u��@woɌ�.�*�8g�qV!�9D	�[ߦh�	#�=5�x��T(��0_|l��J��ٟƠ ���� 	2��A7�^�=x���ipn�g���~"�8�h@���T��}wek@��}+���iz+zدN����D����5o�h���7��N�sz7P¿�	
�iuv!����� zs'k�O��,����	Q�4\쨛C?T4���T%і�'��J"�����j����~�T�Sn[�)�&��(F<<Bq>��tK��#�af��!�l|P�V%�Zq0*x�Hiad����/�Pj��lz����<c	�[{��<�#� [���Vhn����	ק�@���1od*�J.^�-6qd焉?�/O_����⭒26հ��t��!hW�+���mCJo��h�:�
B�Pո8�X�6�3T������x�<Z�j��)�����7�t��t�2��%��kn�\��u�*���W�t�2�̑s�'&ft�D5�B,��Ŭ\>���[��_�@��Bxj8ϊ��t����D�~6�I�S�2����4h
�k�gV�9�j����E��J_?:q��p.'����^8�h<��2�#�Wė�lP��;�⁐�fxRbbf������m�e���W�6��nk���=�/��!�X�c�=�ҳM	$��9�d�>�H����9�f�.U��e]LA)�DU�M�M��)�W^D�ڒ�rR�L���]�^�����^��$�P&��Z��`OC��3��k_�@JXdoX����1 s�vL3qr�[l�c�@��I�pTbH�Ֆ�dK�0C��r mxt��&��@��6��Y(�?�Xlnb���\�$�2p� �g��W�H��dϧO*~ *S�)�.*="k=+�s�Y�:�����
����*Kjٛx�����@ʻ��o��n�$��Z+z��4TԌ�o�8���`�uZԏ��*ӵ���F���O�K�����7%<�&�� �ߒ�ZT��ڹ��br+ޜO��-�ө���l=��ϻ*I���6�p����L�1�mP`��gߩ��!����A��	G��`�G
��p W�H����l���D��\M>�(��N���Ē`��X l�e�#��<�ra2�;�1�����~j%<��	����ߋ*��$�sH�9�[����.���.Z(}�H2��E0���^��Ψ|Q�ӹ��� =�}Ov���0mYmsAp5d�=�R^�+�
r)�� �.�k�vD˧�JYox����c�Z7��L�:P��'�t�n?�oX|A%Z�A3ˎ��o����vn<K��°�$��})����l;��.�%�jR0�;�$ն5�A���}��i7t�0�W&ߦ�6����f�b���Q�e�yr��P�T�I%��!�d�����wr�6/X����ƁA0�|�8D�y���Ӧ�4�N�@�l@ ��v�Y>&� y�f�_��<C��<��d��R��Gv�ʴ���4j���u,����M\2�jf�S����:�T}��@g�:Y��Nϓ�3��� ͵�1
��zG��*�5F�B�#�W��Ɗ���"��Ǔ�����9��;�t�V��xr�>�DE��>Rl���R����M��~^��q�<w��)~*���Ӷ��ȡ��tT �k�&�Cv�������2� ��?&c� u����a��~�=#?��8��𧷶hX�0�lA�D�[E/f3�{ojs�m�~�l�1�P N'�?Ѣ�?�ݱIzlnr�yk��1���Ҋ��~ܵ'}��E(�ݣ�����Q�@3/� #i�t6��  ϝ��0���i;쳌�1}�uaPY)�&��}+�p#?�=N�Q�Z��%&�l���0�x8�Y�A�y��>��b�	L��m��:�(�%D��� Jo]��׾Py���v듥��"a(U`q��<0d�-FÒ�3.Э�Hߊ�Vp��j���!���wZ߷����s+����e\�H�w�\����D
���yɼ�n ��b?݃�a�����>O��6�[�U������ů��H�T�� �"Q�_�h�Q�N��S�-�7L��ǹ���k������w�m�0Kx�
1'OBe0'�t��0X�2���^��}�]4�(=9�����ٙn��@@mL���ǋoC�c� Y����[~Hk�T&���x�k�f��o��kǽr��faH�'I�����v�>mK��'	g�P�O�2��C����tW+�
�}��a5�$B!W`�~=�������ґ����Y�B��w8\QO�dg�s9�T)�����79�M��?��	(����i�������y*zX�	%���%�Ƀ��&��I ��3������e��o5��9����K���i�h��XI��4t[����1��-u��=B�:�أװ�\QJ��9�>�l}���W)�O!�wmYN<2�U9��!�s�':M�r�.`C���Vt�����V�JŒ9���ѹXl|3�e�$t���6s�ps(�'o	��~i-������1XG9�# �e�m�}�g�x1���qт�O�5j��?�>��Ǭy#���!B���=W�k%�(�u���X\l�zty���7�e�E��L;����l�S�����T_���~���.h�����ɁyuSw�M�ʯ�P���%��v#%E5 ���q��i��^�ߗ���������O�\ě�%��s#�.-BV���B@:����>"��T�����)؈&b@Bс4�<���[� ���q<�"՗~�SXܠ���hJظ�s4�|�/[�?�K�+��(f���y�j"U2�'P��D�ޗ�!�J"q=,]�
����./����)�Ռ��M��{�$��h�vǠO��$�� ��A�TW��(� n��& ��!�~C��/���m��3$ˍ�~/'~t�g��ޝ�j��v�C�iɽ�i���^���U����W�Ѧ B�T6k��r�Ph��y�@ڲ�����W����(r�P��].���_�}�����f��n� ��c��g�VX!�l�7/@���j��c]�-B=bn? `��T�o��Dᔁ�-b�}u����[�;�W�i�{�:�YG�����6�o��R�%���%,�J^��Lyy���9+�Wj�)J[��׋�����x�h�yO��B �`NO����E8����?�2-��������*\JM����PH��镯XwIt���j��n�y��G�\�͐��M?��]]nM�p���'�d���#��F���6$.y�Դ*-�{,��l�HIL��z`|ݻ+�1�c�V�p�a�q>ϛ��h\�O��:�$!a'KdsWvLF�WOǽ���)�݃��伒�)#�^'.$v:��"�������hS�y|Ŷ����ס��?_��aƀ��]�mjq��+�1�Ad
hd�������-�d����,�5���ۨ��E��&_�n¼�V�u�TA�!�M7�{�I�E�:6x�Zi=���톈��A�x>e�,LU2��H����AFeB� �����h[Ā�@���U�RVb#��]�cH���O��w�((�~�� .�����M]2Z�_�(�t;�!����±�3X��r�7l�����9��!�
���UAPCp�_?N�^��4 d��lj!�$�I
.vf��e��rQ�<#������k%���@�ή���@������>A��|9C��ۮ�:)�����5~� ���$����N�;���sϜ��lNӋ;G��1_6x���J�U�P�7��1�h�nl��4x�S0#�ϰ-#���p�r�xP>�!d1���WyC�g��<h�Fʀ��i�[v3<�#��:6��O����.b_��,�U	>K�V�m�N`�bgJ1�S���[_YX�Vaf�B�DUK;�r�Ƙ����xf?��oVU���?��;�.e�T��?���G�$
��R�(*���ѽ~�[
�Փ�d���vi/S��SS;������&/y���F>s!�G=%c��Q@�9| ��� 5���>\H�f*Ď�%��1��(� ��)Bv�$ƫh �x�7�ι/3d.��@� ;
����I�����{��۸�QJ St��o��^���.@Ǣ�?G���Pf�~�P��-�#�w�?w������	�v�q���`M����6��v�:ZZ��E�����%+裾4���H�=�
<�G�5�F��o����cHH�I �c�P�>n���a�8J�\#�!�����c��&@IX(��|�(j�6˱L�J������t£MT��-����b;}�bb��7t��ߑpX=$�e����(��j�3��o�*";�Ӡ��[�R�\�/�xp=�Dh�]P����^���}�^I����3�8���I!�a�ӷ���y7 �.B�`�G�\d-�K�9|>j�B�~��	�a��y.�촕�w?5�7���t�n�� /#��T�.����z�|J��,p*��Ǔ9w.7�K��%�4��d�x9؄׳���l��/A�Ǎ׬ə[	� =i����Ċ�d�ޖtlҥ�]�w�P�'X�d��o��
��!ey��\�����n���g�g�ӵ����R�>D��Z������XO(��t\�r�k���I���I�����2r��&*�4!6]Ȣ���Bz7]�Pr��7j�q��Z�r�6)�k� U�tB
\Z��or��m5�;5W�Y:-+���`�Nu�)�ٚVے�86����?M�%�T������J�VP��-6#�n�� t40 ρvWl-}�HH�p�����0[C>*�&M�+�_�����5�8�ǧ�cP�#R&t�!�����z��M�憍�j\"�Hڣ��=��l�Y5��B�w�	��r �џ��{3�7��2��إ�0<�c&"�h\A<�`�K��l%�Ո����"��#:�uK�+r�,`&g�?�� ?�xp�X�����ENho�} /�#|M����)v�'	s��Uzj�(b8�bu�uah�7"O�*[Ì��}�L M�D�C<$���'�-�+�`�H�QǬ�?2p;�+��<jM��ft&:/{8S:���87_���s�Q�*N��
߁���5��5�Q�xB&�	�d���o&�g�;������)��VW ���[���~qcڌ�$&����
��2�{-D����cq������+ ��/�b �k��Uޞ���{�H��3 ��:��Fњ0��)��0 �E�[x�V����^�=R�1��7Ab�w�~X�0z�9�#���<>��V��r��8�%��x�,Ɖ�d�d��S��~��e3�c��ڍ=�=oi���je `��?yM���F��ڸ(@@f1�4$�e[J{�0X���h�P�-�/έ��G]I�1楿���������8Ew&Yy.-$]�8:�5D6C�9ۅ���.��J\�X�(t��8�6�zG(`vD������怠v�lL<��&yX��cZ�1�j���؃�5]2}���o�w&��%��5���n���:�������1�2���	X��
���ނMb���<�:�������ߑ?�R;�e��K栞��("ӁI������˝D.���d�>iE���y3H�0$�ί�� ��Q]�|��R����.i23�`�)t�10��PAw7�M��M=sd��o����xr"8.��JW�}OE��V���E,B��w��^�<�(��M���k��T_0�σ����f]U�<y��R�Y�I|�l��
����;�R�S[�Y�Ļ	
ҵh�����3:�����d�M��'��?ʜ/4Y
�}3�ڣ��R68��)�!=���Fl���wx��WW��?���lJ(x��O�ǉ�����C����2;Jo��A�֚�D��D����ģ�n�m�i���;W�F�K�o��0�(R��_�m�yj�2�6А�{1�M(s����K�1v����։$�ϫ��#U��Y��(�E$"�u˄IX��O/_�T�̼tׅ�>�q�0�6��j���<�5+������ ��f����-�A�2��bj����'r�������U�Ѧ��@��n�q�@��8��C/����;�S2�+�_�8�Ȅ�F/��I�e@/1:�ni?�7�f��d�^Ɍ	�wo��ű��Y&����:�j�,�HĀ��󚞂���c���4--Ĝ�Lk�{\a6o�Ӈ�w�@�4�i*3���lB���s)����MZ�DM2��EA]�Jt��O�`��|�.�^U�3u��oLT��݊U&�_�M%Y�98��	�e��AiS��)$q3Ӫ�9<}�K�I�~d���8l�7$�5��������2�n���;��>��O<���
��s ���keE�ȕ'���'�c���Gy�<i)H2��z��[�B�d�ٳ������U0ߐ;��'e�K"�,�b<���;�bۅ�9)���I�7ȶ#�GA���@/�q�W����8���$�SZ�Ӹ8|,B$�P�fb�ó���R%��&�^Dg�����N�ss�X`�`�{6"�af���"y�5�(�$�P1�ğ6��J��̭�U�9��p������
�TcE��xo:M5�K2Ð�i�=c
�wh����L"�˜0�-5�Ϻ$bT"F��KC7`D�y�0��¿��v*C=Ь����	���_0�|�Ԃ�מ._4壪G)�p1�����|XRHW/Mt^�~���Z�/R��y2�>��4��\B7�;�}l'�W���@m21Ʀ���<��8��sӼ���ㆳ��QF�p�oTX����A2�~AM%�ֺ} �`U�m,���~��X�]����uhQJwR�@R�o����d�'zEaϘ�����_"��m�y�i�����t��y2��zح�?�e�2��"iy5f�G!U�R-�N��Œ�inx�
 �����%��Xe�H�s�Z��
�J�F�4�:�lUy�?��і�6|�����0�o$�UI>Bp�/%Ċ�$��4���̜�܉��z%Ȍ�lw\�\�uQϚ�V)�wo�C�i�o����C��ծpstl\z;���밗'�l2���~�Z���W�ok�^oJ�bȷ>�]!eL�k�r���*�~�JS��b���������@�;rӑfIyjHy`Z��v�_�İ 9n��5�+v��Ʀ�����J�����ɍO#7j�S ��0=��%�6�HM�� �mh�f\��)�׳����f���EC�ػ����(F�H�%4�h7j��H��M�hL�p�k��"l	��1���l`p�􃌍�l{�$�}�xj��N�����%�*ЦE�O�7���L��<Ο9s���d��#��i���7Tį
@��i�.{��i�돎W�z�E�;y�n������P�C%�#�d6ɻ�(i�@�R�w�� CN�10�qW(�2P	/јJ��ZI�4��;ͮ��@u�AƜ/�����H�;�`$b���[[�P�����̞p@J9u5�dJ�e�:��{z�n��iU�@?b�86�(��N2��'4��q�:����D,HH�QU���y�AΓ��#���/��=��H��ם��7�ݠ�:2*���Y��C����pj�j~c�qd�%o�d,#�ڔ9Lg��e���4s����?��e.�N*����{�|�î�^XVa-q�_���H��Q��N̚LԼ(fo�
�,)g'�+�ĥ�n\�4f��S�R5o�[w��k�,��7�d���v��'��Bz^>�I�Ό�$��P��:n�I�3�2r������O��TC��V�K�_��8�D�Le�NTax���Y�R"�P, �.5vH<�F6�	�����ܰx�ǴT��397�����G!ۻ/ˤ�Lq�l���pwoEOͮ����c�8vΉ�hu�q}�92��È��Xү4d�|'C�+�2t�\�#ڔ�3�S�}�Ӊ�� f��;v����W&�?	Ǌ���y�܋,sO��`{�ٻ����>����YP�n���m��FLGʬ���V��ys�@?�Ƽ;��)��$��b��/�-[&'�L>���])dd凧)c����.9����1�+�,�G��o1���+�g��̣��c��� �ok��&C�a��s�5q��0)����o⡱h�qf�#+s諿8E\�^���q[+
|���-�6}*-G� �Sn��N�k��*>��q2�]o�(��eCR)m�\M}5.ٺ�OG�,���j��4�:���~{�d.��z��<��B=F�N(x�+�o��ۿ���Z�DE���hq���Ga��v~���2���X���
�AW�fF0G�4Z_Hw'm>,rVif��׺w�M���u_�� #�1�v'}� +UZ0�.b��Dz�V�lm�@j��v�:�]��g&�T��(��}������h*H�۳�=��n��å��H��;�	�ZC�8�Q�[���}&�z��V��W'������_'�`*�3�E�U5��A.3�T{� ���4������0y��0���'�갚�P��D�k؊ebh�$4�����<N�.�vB��@&�|�U�S��.�>��f��9Kqy_l�����u���\Y�69�y�~�����@��׵W�7 E�YyA�]��6;Sx��g��3�I�7���a�[{O(9�����(:BuvR��q�Ւ�yr���\l��BU.<�<�Q8����_�F����mO�ˢ,���_
Ӿ�{��.�r��
5�*��E�"4�_a��)�"�^~�����_e��� /\5�h���d�-fk�!�N�}Mv��)�c�5	w�ɗ�����n��E@%��]m����W�:�?&*>ser�(T�x;݈�?�6�i �z���_׍��iw�4f�ok���t��aS{ ���=`����Ċ���@(+yP �L)����ڨ�f]m,Q����:� ^_��Y�&A/�yV��=� Zq�y��S P����_[ي!�I�~�Y|8T�3�ޥj�V��P-G~aI�S��dӥ���M�/�g&��ե@��C�4�% q�3-p���7as��O ,����ױ��6���U���������N o!N�y~��{�)��`���;��C1��F���ω(�Q�����;�w7��,<A�B�G¿������Q?��BHΌ�s� ���3��LR9i�7�}�d�����\]^,ߧbO��ut'��-��Ugݽ~厦D�`q�FC�+���i��*I�IC�|�1b6���oMM����k�j�o��������)H1�Y�<M)���8x����t��(K&��6$(�XV��G�m����yЬ��_FA䦘�����'�N�Ho�!�+d�m.G�(�Mk�:>��_$�u�4:;�D�#CY�29�������_��^���	P�F�NX/֛�p��JurS5���m��϶��Er,�m�V�����!��)2���Y�ʏk�Cp�^���%�z`�V���߀t-����G���;ލG���_z���	����p�A���\C(3�#�ЂrA��{g�p����X��+�� �.��֯!X��E�������%�A��+�zM���\�T}���܆ f��}�4��:������� ����6��d�7Qi@�F���.ؿ22���9����Mn��G���׍�c����\��G��r�p��8��p���+�l[D: ��V
}����t����*��[H-ς�j:j��y�/<;�̅��Yo��|O/COH���;���_�i��-�v��g7�r��b�p�C-^@w�ި-��N���ٵW?̮W�Z��]I߁3ǝ���0Ƹ�sGx��wt�s,�렲>��\��3�5i�e�H{{*H�+�%�eG";�%��~�57���.�fQܯF��
H�R��������Ȟ&�-��E�x�^���:�cO0`*�ƿ�/JĲ�j�zK���t��	����i+4�k -��V����w��h�yOx�uO�Fh�<X�~v����sIY�U%��s��*��4�ɳ0�(΄� k~r?q��4R�Ӈ�,GXYV��I���@|�D��'���vv�޿�C�û�\*�N�kUk��Z���h�:)��o};��<��b,"�/~W/VQ��t��Z!�`�;�y�Z���չa.5S�gN[���!1�i��&��#���Am����ɘD���C�OPh��bH��C��i1�w��o`��*�6;�sL
/K���Q��e8�_�X幓=�?%\�\�hH�f_�I���a&-�k�������F�?�H��E��'����9cR9O2�ό��6��]�!�iz(��:��m�v��"/��
���������N������|���Q,"4A��D�f�,uln'v)�;H�2v���T���v�:m+cq��kڋ�S^�; � �c̀m�=J���.�������C�7(2�f�u������~/�gj �/ד�}j&�=�_�'�W4B��o�_��u���{ ��F(u�iS�I���X�+Fe����ȫ��L��L����:үU�4	���F�-�x����t$�	���t��	�#���@_"6M��t"0d8�n��h!.��+O�-co��M%���Rp�z8ڀ{�c> 3��P��]�TXC���혱�2#��?��"0�`�F�]C{ev!H��h�//ē7T��k�dU����8T�d��`ͺގ-�X��`J�!2��֔�C'S�~��`�?��c��ݠ�wO�	n~�0jڧ3K�d{��3ܸ5�A�0*|@3��%"Yup�cX���hT��+�awP(T0�-	99�Pw��-�;aR��$���g*�S����W]C9���uh7�T>����*nDc�c� 1�ud�Ҳ㰊,%�	,9Q��
��-9�_R�q�/am�Q�#�i�D�GxA���Qg��䶉RXGG�b51&T$ڤe�1��S�p�<*���Y�E46?���b����/�������ݯ�?�B���H䫱6�B���2i���c�&�'�!J${ߺ�@��!Q%a=
M�*x���?�>���(��G�/�v֮�/Fu�e���j��X2��IW3�/?�6����5_���f�H,74��~ֲp�sq�Ŋ�Ii��<��R�0K@�������˱2`�!Gu0�T���~Z�㟬y�E8�d��@7}rd��M��k?�ܣ�*M�Z��l�s�v8��c0Q�V��vX@d��䈦(�M�Qmqn�/���N�rŭ��Hx��sD&�Y�\����#��}����^��$�~�"������F{l��9�+\eCIk����`2�@�B@۲|�E]P�	�����5�>������q#��#kq9B�ŕa~1�i���o�h%��HF��aAHBr��� ;�x��3�x�x��Ӵ���H� ��/��jk�u6H&�]�P뽾�a�վ|�,ĭ���;�	��/GĲ��w ����.�z�j��ZG��]
ڧ����8$e��~�ߡ��F�tΕ��fc���ȧ�wb#P�Vδ�ڿVW�:7�#���W����-G���B^!��'D)2�8Ɩ��������1a�+k=<l��4�s
}կ@�,��
�ѿ�I��e��X��tJ5�wE3����Zp�z�A|�P�� ��T��t��+m5����<��C��-��]ɥ����e�vr����T��1�9����Ƀ^�D�̴���_!6�F.9L����S�/֗D�E�N�3�'�ׯUA&�+�_ۃ��.������C�&S��7��~1֘����N���(��m�)d�4���%�1��PI�]4iQ�?�Z?��IJuD���ra~*�Cs�Wf��_��)�����(��S��̜.fjXb� 4�9A9J��K��H8��w�%��R��	�o��ݚh]��n�g$v\��M���Rٗ�4������.&$Y�*c�i��7��;b�].����
��S�+�F�~ �[.af~N�8�HQ0"`��~�,k�Tk=x�;����X��x���� �+A�P�x���.KU4�9��S����3	�.���B48���n82�ψ]�Q5mVcb�HR[:hm���EAF�������Z�~ο��UT��W�ש/F�YB�X4�v�����PXi����G35+_��$,3�f>+��$���WF��!��D�+��g����i3	�����L�ɏ?n�o����ݤ����I��t�3�QSz�C���)�}Ԋ�D���:��*���@�Z�0�6K���� �P���������[L�I&a�)ۋy/�EO1�o"���z҆�1;���0T��W��E���WSa�,�Ì���9"e*�����E5V���a�����p�.�a�簱�,@A���W���]��<�"/��R
�(�+�h��$n��Ty�ݧ|�y"� �J�}�7*5Lf����H���Tz^�;����\b3�.�QR���iӿ��7���/@ۨ<��j�ɖ���H�d�w��Z�?�� �ą��Q1��g�(����O䊕b�ڶ	���\|�þVv�2k��gG��rĀ���I�H�+�W��o�jԽ.O#�0�n������"�JɒT{s�:!����3�W1T�����}�>]��_?U0�n�[P�T'fW�o̷V^�)���S�3���`��h�a}�,}$�����Ba݇�#|�Gm��ù��}�9�/����e7��w"p_��V�'�l����-�O�W]@�����	�������*�^��0����]����!V9��K�A~8���]��P �+��NoWu����o-���R�F�G���H��I@��'�)Ƨ60�5z�޵[���~������iO��Ep�ϔ�0��=4o��vĀ�t�	_��)J$��t� s8
��G�\���gDK�Z�6wzx��58�UY�miN^̛�U�-Jd���]���������5~�ѿ[HzcPLjk^�/A�[�q�	\Z���@e���Gi�F�u�M���'¶�T���CS�r�B���=s��яbM�K{ѭ���䆈���Y0��Ȧ)(��ɐ�*F�S�P��`Ҥj�ĺ����K�C��/(��~���]�<;{�;��~So��qel���gIh��4��A:[���l����|����y۬Bg̹���6د#��ڟՓՉ\�s��z�|t�a�`E�.jR��r��c��J�o��X��E��a�'.d?�7))���ǆ�7�b�U�,���C\���ZO/U�G����y)ڇD=_��@���k�{�qP�`�Z��,�:Wc]ޞ��ǁ�ѣ�3�::�r _���b��=ZD�����-,��Z���.a��`��*,6�4 ��t�P�61�3���ؠ�.�&��#���%��lAp8
�s�
7m1">s��׽N�9x��0�9�G�E��d,�_|b���ːs���Kڈ;�R���# G���M+���c���� ^%C�������Y�y`>����*���&=y��Ո}�&H�������Z�YYW�{�K����ޯ�������|Me%Y����я�t@�\�n�\/��k�k��J�,�Ѱ���̈�s����+Z��Ț+�*��+��@��D�/�����d��%]D"᧵ģy�v��a�"��ł)y3��f/L�?����1>i�6�l#20�59_omB�W�8�(}[� �y՘���19X"[��]?{�ܮ,0�|B�V�Z8uR�X�r�7ĺ끆�Ps	�A�zy�׀��p#�߀q[�R'�	�q�Z��0��|Wvl� ��,��Sݕ�ǳ�싗i6ǽ���Ab���F�tנS;�c�CDN;�� <_z����X�p�� �bU)UK�:���`�%��{���σ��x�Q|k;��)U��|%3����_�ɚ�V@����|�D|�Վ�����E*,yJ�b�)<�:�[D1\
]����|<6�;ig��3Rjǧ�o,�y#���]f,4�w���۬���~�y�|��`�_�����2��b�v� vc�n�,יִ6�P��3_ܡu	�͍��Ƴp|�V A,��e���Sw�Y	;�+}GP'�+�o���%�DĄ@c��P�C�Z�I�ț 
�
�D?^�?/�K����S�~L�6�D;?����*g��5��Mɐ��n�u���5�>x�y���୶������+=@u�����q��2�z����"��<�z����"pH�-B;�J����q{��F�K^��=��w���
�y���|�'��,(�}\����`���}��VJ�dH
Is�����s�?�٨~:2����L �A��0�����K�K�C  ��i8jv	�t
ۢ�;�Fb��C�{܌�F��E�@����������˭����r���f�*��t�<aU1FYg�.s>G����}1�ʼ���\��O7C���w�[��9DM�}��V�Qs�vޞ�B�wm�[j_%����kn���;ɖ�Ch�@�y�4a5M֗Ė��39��10zلC���������3^G`fʊ%�VW6��ɭ��}�!H1 ��m�U���GR��ei9m�
��R4�;ؿJ�����D8�8P��y�k����8�|ȥ���8���kq�#��cI�q���I��T��-����� TP��b��m��=V��1��1����2g�6t_������ڎs���E�~e��U8��ި�(�*� x�gR�����������`/�C�G�J����m�Ϳ��x�ƦQ��ӊ}�"Ui���� 7�n2�$U�G/��Z��w�x���������x��)�L`��9��TH�E� Jh,!�p?������x��ͰHe�mr��2*�&��E��q��M}��:l�ZW��U.?��������hY���m�9��ҁ z�f-�5�*���q#'�T �1s0��	��3�3�_�q�N�z�2��yQ��F���R;:j��n���m��~ <r�^�dX��.|�.D� ��uP���k:�-h���I<�&�XV�������Jd-���9H��I0�}Ad�	�ն�=�&e�:�g�J�oD�Z����sDMO��Z�Օ�_�2�,ӥ`F�:�����?��9�_�*��a�ڧK�a��%+9�!ݮ�x�$�d���)�*�aX���L���A���ݼ�l|O�� ��N���l�<e%`���v�9{���I�  ��f}G�hb��BY�4�W$�@	��t;J�c�vn��A)�b�P3�g,d5	�+h:TE`�%n��������'����Yw立��>�h9�ѭ����(5{�.�1Q���/��o�P�`]&�%�;�w3=�#��n+�r�n�E{�0�n�T�^|��V���jU= ˰�NC��ɥѮ<*GEO ڿu&1��� ���8�B��˞�����4_���!=Ui��հ=�z%e��FM�� ^y�����Fx�iR)�R�E���r�M8��Cǔ{g�rh�&90EM*�����ZEL����Jsz|�. WK���׍3����{�J�n���$�-��Qf8�� X�Y�_��^i�bQ�����d�"Vk�G�ɰ�-��h�������T(}(*�%u��/ _3{��D�?�ӫ=bo�0B�QZ��!+2D��@��9�LRA�S��M��I�H[��w��
j�SL�fx�Qo��SЈ��)+RQ���j��"(��7���W9�c �F�����\d"���6̧�J��^����E�3r���yh]G��6�Ejҟ�+	�p�迣�a�%����CQ��^�<��ϼ4����Zյ�	��ӣW���jd��)�ε�s��6鲲�a��杧ohO!��с�"7TM�7gB2�֝8��_�M��&	��D`I���Gyx���ٷN�H�ta.���,Gϱ\�ry�eᤷ��6	*���@R�q��pI��X�HQ$a}� As*q�<�1���麟�e(з��?u륡,{�lݖ�G&�_)`��'kH�+�Q�ӝj���k__@�#�J���='�X%X���~w���?{�/�k8��>�j)�%�y��1��q��Dk����x0�(�WI�<�Β��
}�q>oTM��)
���v�PEJ�U��EbZ:W�/ߊ�]-�$�J�@���8�P6�,�}���[j���Δ� �P2ًξ��?���p�[�3�5W˓���7x3%��aJ�����R�s�FHu?O垑,�T*�꾷��
�:�v�����g>��`'%�s"r�U֒`��c!u:#��!F$u/��j˛u��<1���I�-I��Ǆ�x!�+x*��/� zv��5�ʳǘ���;iE/p��x�f*3��__o�����a����y��p��?����	���"$x�2{$�O�	/؉ʒq� טm�����U��%�Zn=�Hv&��17r1�G��*��e���T6!�3�A�V���9�>���]Gu?��t���?`���t��X`���1Z@ܧ�8_"�hA< ����(��绿�Pv�>l����є��=R甚a?k��{!H[�a��Ψu:��DԂ�;�Z����gu�q{s�Kn.X�t8`�Bs�Ϭߜ����RA�q}�;c����#Lu�E[ro� 3���:	�@C�~��z��?���s�q�0�8�7v.���BZIL��Beĳ��K������r��KVY�<A�㊤�kW�Jxg8��ˉ�}�.9��f�}
Hlǃy���z�q�'oW��~/�I#�^+��J��D��^���N3.EM�[�G0�JΔ�[�%!���Wmbf��|6� �-7#��`�:����1j��`���>�}=�&v�r��q�F�4t�Z k'��'�u��[Q�����D���D���ܔ&�UdD���X5eF��sܿ'�)8��k�[5��s�D�w��W.�q@������5��Sk���R�"�sq֕��^\8>�����{N �Kv���?z�_3�l�Li0���	�j�ۈ%rzsY�C�֊Cm��y Vͪ�<a�t�\�ɇǵ!���� ��+9�*ʝ4v�{���k�մk�fH^���Tf,�>|̨oB�c%�#j�Yi���V@f[]��i�)K��/�v_gs^,��u�G.�b���߮ʤ��w��	{_�,hSG���Y3��^��qMQ�p���/.��L��/]W��I8�9z��޸�n����>(Ļ
.nw�7�(�B)�%ZE�8{&�ڮ �4f.�-��Q�v<0�kU9yn��>öܤC�3�s?���hE͕���i���x�����R^�Oi�YsM�̿� �Z ��9��d���П���x���̀.v�40kDb��/�q�k�tz���`��A%���Z�ğS�cE(BRpA<^�>h�Z=�&�*��($2y=��1�G�Uq��⺫���|�b���`�!�|s���H�GZ�M���rk�:�0h��W�&{�2C���/5V�1F�x�a{�v��rz·�z$,S�]�� �]t�!e����.i��Yx�<\aȲ�G�,������F	�|GlW ;�b����Ya&�2R�&-x)���������jL�ck+]hq��:vp���PSs�Ӟc���FM��m�C3�!����QҰ*Ur�����{�k�C�K�F�?%�����@��4We���ŖRS
1��ʆoS�����w�:�h���w�\v}{�7G~X�JA;�����FR잆�˗#��E��Ԅ�t�]I���G~�gz�W5W6vp�cL��8l���q�;GqkH��E�n���E�����j�r�v�ƄT0%��;����{!���+*m`��>�_d���(���B��z_Av�HiP�=cN��ZΈ���j�&jZ��~B�$&-C���|�l�3��� ��p l�fh�C��З6���\�����ؓkÿ<;Űj��x��0�P�)�GS���|�97��gz�����C!(,�ېt�q���SjR`�3�(����^1Q�����-	�]ϲ uו���g�@#ϣ�<�P�1@Q�;��4ʸ<(Yw^_�[y�)�e��*`��tɪ�'K>�W��Z夶gw�W�׸�"9���ǭKV�����I�NI�'c�/ʍH,��+��u/�_sQ��3�j]��u3�Y/]��ɓ��������ǒ`����T��:����ܹ :?�i�ό�YRu�>5�+���I��x���;l��u�"��ۂ0��&[�(��4}7�n�Š�7��=ø�+p��w�DH1N�,�ۨĦ٦x.h�a�.U���`�`�}�E*q%���ےN�Ls�y���H-8�_#�z�s��5��0���8cB���*�תN0s��g���0��:E����y�]�J�GW�I�1�#~�>C[�<�ş@q��ȅx>���3�`�@
j��|_Wy~Z�E9�UL��P:�PPEv�Q�~A�tN���03���I�X.(��`���{�!�&���2c �2��f�����O�����gв�̉�ɤL�ȕ�]�t#�Q�iP7!1�Z1x!����
GLc���I��l���xB��nv���	��eȊ?��L)�����Y�Fˠ^8��|���O�����ch�ʰ���?x�t���>����Fc��/��^�)�tpB;�>Ȑ���	cGD9��m���T=s9w�]�R�ԫ���]��X�J���ɒ�����Y���=<U[�|e��A2�)S�m��7��Cv𦾵?Zx=lj�T{y���\�~W�_k$aFgR�Uz��ͤ^�=������7�d|YB�P^9����b��F`igi��Ƥ!�P�����/Rv�v��_wض<�)��?�i_��L�r��3��Gm��Ѭ�th�5ll�E�wzApsKhw�hv0��5~+^VuN��-FY�)�#a&�ӈ����#sJ��[^�<d*�,�,+�Fd���A2t�,��t�T,uq��\���2猈���>�]XHOe�	Ζ
nS��DQ2����q�XJ�44�?�BK52E�hrO��k�c�N�%��6��ez�~f��/��n��� ���w���1M+D�6�Q씘1��k�i��d�����&�sl��e���K��H%,����Y�S�k�2/ȑZՓ�R���r�����8�Fp�~h�V������OMl���H��8�C\�:�9q�'���|b {������al�D��F�noprQE-O}~S� ���y��of��T�%���/�'���
}:=B^F/ �u�I��9���(�����t%�֝��0��Â�l���?�v���e2r�6���G�,ѐa�,���G�� 	1D�jXf;)?B0��	�&��,�ژ�p�r:A�̨�(����?}��g2;U��am���/}V>���a[qO�`�h}��V�`�L�Γ':P �EN�궷kG,��-8��<$H#���K�<x�uR(g#��v�����ɳ����j�/7D���		9�y�5_�%��C9\���������l%-��F>Zl�Xcm��s�.M~���٤NY�)�.`Pn�P%a�ڐ��]E�r�p8��$����kq׻z^���0��0ы�ZC��e��U��g���]fq�p�������!1
�v��@��@&M����tW�ߛ�S̫Ҿ����������Rc���Vx��Rଘ�0]%��w��f4񊱨"�[L��2v�0u���И�`=%S^�U��7"���6�9��`�ws��e��`х�"���j��x���v׹�}�4����ts�Y*��X��g��Ubц��t��1������W流����c�+z_C����N��g|�gF����� Nil������aT<��yx��06#�U�[��3�0�ߧ뻑�ͬ�L�`YTvS,*t���8��rZ��W��Ѝ����H�8{�[��h��������$�:���O�H�)�,�S��xI«s̘|�+ػ�ӏ�����\ь?�XW�o����نO�u%�$gFh���,�+S�@R�0R�Ѱ=��r_�U�'T�m)Ⱳ�d� shѫ�
Z������@�F�ě���E�>�����|��m�+$�_��>���Sj�}s/��М��^6��t�	�r�8���u[|&��2F�[�ሟƹ����B�H�I~�����+/Y�����>���R��4��b�4n��C��YC^�zS�T]�{0�(�'�!l߮��懲4���"r���Y}�m��[N��d��S눏:��xT�,,�
��+w�R�pdr�H��8V�0o�C�"hX�R���.g����ήה���^��8fv��cq�k�N��;c�B���q�v�Y|���������׿�5�y�-cyP�*�U�pb\�D*țr�������%D��d9$�6o�?��S0�Mg�	}UxV�'(N\�z���_���/)�_<Z��Xmi�t۳IG��Q��2�(v��۬jQlݼ����9�x�w	��Ь��m��	��������/I^&��d0���9v�E�4P�b��w�
��	�s�+��x�|�h���}2�18�d<�&�A#���������_BusJ��������yQ��_�Y1�,b-�RpaS��N���d&�z�@	gD�X	��t�N�+��J�*��1N	���{��Tfl�|�k�HLEoKahz�y�r��O��DcC��#�y�꽆@��e�W����$�^���/1H��:bݻb�"�w�F#7�LK ���6թY϶��oV0��;�����_`2�3w=��@��̴ �`V��ȣ��c��O#�
�{r��8G϶�FX�aes7N|�/&����P&�г�/F�Z�`鱽DM?�1���xF�j,��.`P�D��;@��X��A>4+���h�(�+�a<Hp7��seWi�i����kP�����ʒN�2�X;
�b,A
�+ĺ^��w�f
�	h���[u?"��_��|�`G2��������U�_9����`�GW���0ϤKBې�RX�n���x\Z�1z�_}w�t�B0��	��d��Qq2 d�����!��ф��{B�}=Sa��f\���nO�Y��D�NY�l���,�ݺ�U\d'mv�Jb��/�[��QGP�g�7�%�A�B_|�Dև]�s��B�fmtp��+�������Ϝ�\�MG�N�|��Y:`��c�Y9]�5��~&�U�?�������U���v�Q��
��>Zd�'�5��n�b\���F�~�r��*��-v��D�Ψ(�*��*�Y�Yu�����r�L>1����G�P���*��?m�r�\����qNNf�DY��cNPfy?�n<N)k8�m�C���v����Q�?��ǩ��Z��L�!���q�j�7��ї�{���		��}��gma��HDW�p��Ca7�*e��^�8�a�xB[x��J�"�e|{���4�G�������<(�{�e'���`��k�^d�и��w�A|�3�N�y����L��v���dk�\qko���r��� e�� 2�	:��iZ'��הּ?d_��}$*�9�-slc�D�JP�t2�f�_ܟ�0�5��@|]�[��黛�[�̢6��N"�NJ���Q�T���N� ��D� ��*��Ҟ�;��j��L'٘�x�E@ Зģ��˒�+.�U9�%JF$�U7'��g�5U���3��@w��_���W�,%�ݡ�
(0��uE9f�DJl�|J#�S�ד2��!�tB˞�l3���H��7^󩼍Y��kn��Zvi�AU�[�)c�{��i��uB2�|��.y��,6t��q�O�2�?:�~�Ab��`���V��o	?���˾CU��Ui=_ܪ.^(\��E�2X���ȃep �č\O�������˕хe�rM����o��ɏ�׌ߍ@2��ZAj���@�y���d<���Ϻ
��s=���̶�e?T)^E�8 ��=��Ub�j�B�L��]��x��9_Ԕ�n��*���7x9a�^���ࣨ�0�ݭ��8�m�)B�+�kQ�J;y�tC�%����I�����KAU���1��w�fe�N�<���+�cЙ�}k;0��^h���m��|����d�������h
��8�*az�*r�g/�o��H�`�?C΂�'ގ�^L�F���YX�4�
"�I��so����������ײ��xݼ�� �O���r�@Z}�X[X�A�?-��;�LM��4�)ϊ�˵c7R	Ń�Q"���+�J31�6/���m���.�F_���	�l�^��lF���ҹ_r�X�õ �D"OR��S��6rV<����#X��]퇑ԄI+a��hm�zf1��8Q�U��|���P	.lw&M����,u z5$9/b�k��&��u���z5VኯG^�Nƅ�zw#Q�3����ۏt��S �n/�ܻ���S,T�֣[�I�;�dŔC�*���xn���Ĥh��~l@X�t���\�p7��V�z�'!��p�!`�/�<�\pWM��+!����;�WP	�
L��b���-�/�EM�dٛi���a�8՟,�~���M�/����|�ӧ1J�TcuiD�f��ń*��ZKN�9Yc0�u&�׮�_�M�}�5��J1��B�"���o�d ����$�xE;eS� L,]��"G�'1-��O����xJ���P�Ԛ�k�>~�C��T11w�^ ��x�1���<A�>E2|{����Ş�/x�jf�
10��Z6�N9_�1c ���~fa����!5�rf��F:��AlȲH�h��6H}��u��keL� 6t�Ҍ��a/��A?	Z���#R��?�7|�q<0 {�)+�� y��i�S��u�.鞔tZ�~Q�v�7r������1ph���+� �
dr��Z���+9mL�ɿ{�'Nz������/`[��.ϲ:��P��V�b����f�*�4��Ŧd��Ʉ$�Aj�S�Ș��}��a��/أT��KP�P���@���x��p�Ѱ���@�S����|�On��[=�C�x�G�r��������2�ZUr�:b�T�j�ͯ�jgN� F-<R����3���ѩ2$�
�_^(�5pg`Ey�!����U��J�@���f���1.o�d�r�"��*q<c�%�F����2�pӸ7����|����|	X�b_s�����9� sv������jߕ2bj�"hSl}���Foߏ,d�/��h��r���[�i�_nԎ�ӝl�( ��\ג�DR�{8̓������s��x�[G�2B��9���Z	(�k"֍��	���:�Q3��J.}����t��55�f�5� DC�M��I�қ��g@Q�*ZI\v���Q:}�� �Z�8���I��D���)�p�~�(�X�����ַ�xb��P�����a�Ո}�;O\�1]g�{�ʨt�vq���+���j�8MI`�ۭ5���u@[�A��?��h�-ͨj�����s����}X.�&�d� c⮞5�����sZ�z����j'�8z���v|��*�'������ml�Ҽ�����e��R�$��O[�F2��<e�kEܠx:�w����D��k`p��k$|jZ�3p��ᝰ����Q��]�{I�
�T�0�qez����9UB��F�Z�����y�g�ۢ�V=GJ-f����~�;��S�+�{Iri!I_���x�)x����1�o����G����ѤS���6���
�;��`���}=���)���!�����-Ӂ�ĉ���}�%�ݶ��z���Ҿ���9�a_�T�J�F�����4����I=�"��c��2r����|��GS�O�w|���*��ZdM��yU����0WL��~D��J6���b�����J�VB�oS8^��ԑS���4�������I\n*ce��K6�I�FY*��d�v�#��ko�(:�Z��F�y7`�Y��T��!*��;w�1�i؛�US2�*L���E��C�*G�*���,�[��r0����84A��J�l���ڎZv���%�����kقY������M �2s/�Z���D;W����ϒ�v�Y����q����QL��{aR��i����v\y=���������+0�,�D�/�o�ٔ_�x�1Kp�S��ޢ�4^�����0�ɫ{p�L�Ȣ���@�@jWzҔOrf�PX'���>�j	F�$�^XUS��,J��g�ljd�5B;�!���(�m�<-d׸��H�0P͎vƶFI��ȵ^�a�AT��U:�D�7���aVS-�Bk����Qq�4��A$�d$����[DS���P�Zi��B���]�*�>^�����M�����D1�P�T��x4nx��SA&����K>�s�6�8Z(���9�����=X��T�y-�1���|M����vCg��*��Ь�A#j̸��Oo�Y+��E	v��}Ӏ��zyMS)�g0�u�>�UgUZ��0�=}�H��c�����3��h	{��c� *>��)��{�>ZMʗ������C�#� 5~�R���Hy��4�l�k�w��E��l�%_�	EP��?c��Y���=L���6Ӡ��&��Nۤ-��<�/a� rRG�Af��x��M�7/E_�g��P�0[��Cfy��1��ɝ���B��}�K<M��k&�������L&�Ld�����dG
@��/D�{͙i�M�����/ͷx�X������cѪ��<�,x	���FC��%������'ǋ��
p�M��=�J���לD9���϶�TV�cϑ/wYK�H�I˚�+�i_|N�v�	�����w����i�Y�:C�'���khJ�&�!L h�]<Nr��yn�y��7�@~�D�g���g�ssܖ������~�ߑ�ش���o�B�߄����-ݳШ��V������ޑ��h�d�� I���9�М�u.��
0%�e� �&a�f����#o��\Db��%��`�����2�O�!gV�QM����>��ͤK�ft���]S������X+���Я��U��9p���l��c]:���	�\���	iD}	�0BM?ug���� <�>Ø��<�K�����/���^{��K>����"�a�G�0���1�Flj��̎����^)2�1���=t�e���^.�՟Q�KiD�-�G��Z�L>N0����P��&P��?�~����F�ha7~vxOq�� �kj7�ĺ�Ә=�9�xº����%�h@T@�]v���=LH_Gۖ�+���K���C�Y[�$^ ��M��3�;��A��~��EF�XC/��D�C���.�y�f��Dh�QMI��l{�CZ>�v�5������=��@���to)^�3��c~[�x�ٯ���~ی<��槢�� d��/���T�n!}���k�4)Q���H\<GCZ��������m������]I�Cf��e�r�b�M�ԇ�~0��(���� HӵA�&iO���Ϝ2�����s�N��J+ ~���&��ڥS�}f7�\&wzF �t�mu7�����^��n��#�
�B�jra]�UFa��u��힑��|����(O����&u6bܶ���/(Z�¿]�J�P���I6��;$W�Lpp���'��O�q.P�?Ts�#O�v)��۲	������zg�u�� �lS$ ���bF�g�*�\پ��r˯�*F�9M��Ě�k�u:�S��o�R�@δ��W����6���`T�bn�G^��M =/�� �ś�tJ7��Q*������P��� �&�޴��_�����@���l	�N?�~>���<�9Mo��3����(�p0�J��N�N�B��. �M��tC�;Y��~Qc��H0H�OE�ucY���}�q��l��#��>���	�O�ECπ��7ein��u�Q�D�׻T�uwO[�Ż��7ku�q�K��6_�6�g�C��_�eGZƱ�׵2��G)�*X_�����\LW� ��	�8���F��^�+��Pɮ&`W�@摾�
!��ᣢ]�k��[Ƹ��ɾY�Qk�̑�h�M���=��o�?\��`�7)�����b�|��0��%�A���>���ngz�y	����R���W���}�s����,���}��!)�1F &�S���$�S˹�1eTe�5�(����i��`,U�9�L�N�
��
o�>ܵ^tm����j^R�n?�\�ݑu�{N��8�Y\�#��b��HT���p+V-����mLA�}a����A�`�^_H��B�u��f�_�#���ANm �u�~�I�_�a�.�U��� �O�:�vrB��v�ɧ���]�x����N�d6�,wc�_?�A��d����F����ju����2��T�ȭ ɪ��Nv++��p7}����.�%X����F�	�]����
��m����������^�����ڪ�[;���'�_�-�	@]�k错=5�y7�Ԃ�F��B{ڗ8�A�G�]t�cL�᜼Cj�H�V]�I�~(��@�#ךg�tx����h;��![R5��Q�4��H{��g	���xγO��]p5��i�rv�,����{B�OM����n�+LЁ���D�5�Da�[� O ��Ck���*4)$e�B�pdZW�Y���QB��3��V�-i&�ɽQ��@N0��JP�K�{> (�q����A����ܶ&���
*~0v-$�G�m�6?�aZ�� �~: a��˓�iL��LGP��T��\J�T�coTV��>�z��*�S�W��>��3�B=l��Ҡ���M�U��Ǐ�hRW�t�DA��_+Iڤ[��e�F�/E:E�+Vx=`��<n� z�ݭsC4)hQ �g���^Xw�w*�)M��)/��uLJ�\�-��U3#�Ԥ+T�?��ճ����[y�}jg'�|���g�_�h�������5~�R?�>�[��P��0��0zJ�2��sQ�F�$����@�BhL0J�`��(!� ����z��gt��"|��v?�>Idc��F��di�O��W�r7��2):ۘ��>����Ł�˃�|i<ɣՆX��x�F��7�*>B��IEj����bi��HO��y��1��~<	F��^����V�f����X��/5:�k�ʍ�!�r|N�<�'�$P�?`5-��mz(���ꦔ`y�B�B$�������yJo�e�8�p8z�j�{K��|?��S����	����;��vW�yuO�P��d��uA1<vn�i�>e�%��?���5��,܋��������/�S�Fͪ�_ �ʹ�Ѣ��p��,�P�?���������*��K�>|Dj������7�,Q��?"���˗4�`���[y��yP׌$���sy&�R��xx���Ah�E����њ2��?�:�W��Pv�L��Hh�- �Z�J6��Nl����:׼4��Cǿ�#�B�j�6sRG
�����1�L���$Jh	�ɤelS2�04 	�4�so0 �2�4TÉ�y�����p�?�<��Usᮨ1_!�%���R�KOw{� �A��Gs��n��4�:v��v��W�<�����@��������hq�fhZ ���]:�H�H릣���Uj,ɥ��'4��	w]t������>,U�3Ø�R�凈k��ؤq��莯�]��k}f�D��L� �u����CJ�_v���b��"�����r��$}t44})��P��b���g�4)�v�=|m*�܂׿���$l^|�d_"g�#���`b�2ةU�/�ezC��h~?%�C���#����ժ��3W�>=��@|i�~y� 8��qs�����K��W�K���g��>Q!������AZ�3��,��oiR4�Gg� ��Q
T�N��w�-S������pqkR ��@T��ηM9����Ŀ�e���2T@څ�
M��{X�v��Rq��0���Џ��$DQ�r 󰳹�Ix�0���#Brt��R� F�۠�z^����T|�yZ��_�/�+ �W�$���#���k7�DJ!=�{Y�Y
�e����{͇���2m�_OK<����U��*�2:��U{@p*�|�r�z���e=Ϝ�}\V�`��{Z�)����g�NV�|=���;���KM;�L�om�h�t%�0J䑝�f�nL�pU<s���I��:�F&(p,Ɨ�2Ȣ5�H��"��f���>�N��xn���ۍ@��+�	xc�0bt0~n��|h�K�n7��F c�g �̶�Y�Ҝ=~<m7�R�� ��ac�]�� $���d	͛A��<`e��h���t|��`�'|cZ���%^3H+�E�i�Čdx�a���������=����ZW�M|?��5&09��E�$s1����RXF�m�;�ޱ�5�R
��R�F�\;<k��F򁃤�\k��bU+�D+��38�޿ZƳ������z�m���" ��1�ذ&$�CgK��ub�����?2وWu��,��� Cr��V�*UJm�.7;��[�A�ڐ�\1�>'�q�GF�@˒�;Q����Hc�W�8v�^�RcsuzO/�@�R����zd�/�8�Mqz�����6��u�P��t\Z㭈�`&h%q/8��^I˩rr$�bE�/�a`���e@�n��P�C�x��!آ�Fec��8�LW�) L�	E*�_�Hl��z�S&��=�s�ĩX!���1�<�x�qt����{w}{�|3�j�E�[���vODy�a�s:�l��&��������^��;��$����~Z5>�����>i٫�]n��h�%�C��F�HG��Q�rki���L���rØ&&���k=�3R�,��SI���2�|!���֖��69H�YS�^�+�6Ά�[�� �j������z�m�C^8#����#�§�N����Q~<��I���6-pk �]Ԍ�R�\�w��#�9�S���M"���o��)ɹ���� ��b�o��F�_7�;Ucg���a	����5E�6_+D�M̂{e����g���J9�-���c�_�
u�g2^�?�~���Qʷ.6�__M.��>7Z�=MOG=dۗ�X:�;X�������5���`^�"������Aŧq�AJ��D^�)A����T�Z�9�5�]�y�U[��'6g�e�-�u�>**z"��୺�;��޴]�ݺ6�A}H�p�s]���>P$_�9�1�R���5t�̶��d%V��k#P�����q�hl90�6�{�2�$���1~�yZip�w�+�\�ܽ���)�2a�j�Јi�}rX���*Սr5����)D�q�8|?`�O�Z��q�%�:I���><���N����X��/�0��|�z�g�d��}��ha�뽲x?^jI$4�59�Ӣ�&�¦7�uU�X��L��)���b\�=��
�ʎ;�z0p5��9��jTt��J�46���\W�+Mq�5nː>u����>�(l����wED�Q3�bb���#��zIS�Iu��o� �N���=���\��:�$}#-b�*M/bop#T�>��{�á��ɟ����g&Y����DL������	z_�/wDO^{j����0�ڽ�hj�q���V���=��LlK�/�l"V�Ct*`�ۏn옰_��9��D8'?\��NwL�����4�T5������e�t���;׶i'��?"2Ck��H���@`9�ży�2ar��_p=��/Z���q��f�m`n��T�,�����hC��i�8?��ݲ�V�ϑ"��jZΒ3��ޢ2M�a{���B��V���^�v _J<Sϕ]1ɽ{ԝ+?*4��jP>=�d��mjYc��S���	�Uh��j,7��D�>��K�b�O��d)�cv��ߙ���u`uA�ӪB��&�?&�-��T�v�Y@�>-�#�4$~���"?�����K�1����n�
��9$�c_C)�e`$B1xKr^^-�P�$�����B�W�:�ı@����-y�� �s����|��9ֺ�t��ʰ��x�m�r��E��t���5�aAg���LKCpH3�X�J���=a"��3S����rg��Q��y��x�)ϹE跄���܎,H��w�i�Em��3��w�F"�*�V�X1�z�JE�X�7�D�EЗ>)��-H�;�e��+��>YvӴ�p?�G��\��8;��}�L�_�z��M-z�[z."{h�
<�����
�/j�9�E6m�\�g��'��K��d.���U���B�m���/�i�C?Ӳ^K��(<xM*|�G\�LxQ!QD�:kJ+���� n�7�<�'�]���?zգ�S�oGFӗ��0s�'�� f�g�ߴ�ᒼ$�Cm�&�V�i��7 "1v����aE�-��ƾQ"Lu�;S�
���IF����s��*��#I�*���+ӡQ@4��=�.X��+ch��\Uc`������:���������z*�&31��/�%�`�\NsXP^�
��$�b�Kh�\w��:���H�����0��`��BM|z�9�uo��g����(�����9�#5[��������x[���,����T��kf]w��^�Ӭ�rl
��#x����8��f�D�x��޸��7vy�Ŀ�y�J�TJ0ī����o�@J<������e�+yS|t�	�+��8�6��X;�xHl�[�d���9CTB�eA�A�~p2f���u]��>�%MVy'm���{aR��P�=8 )k*NV2�Թ��Vq�yV]�ܚ8������IuuQq�u��<(xz:�e������T2D$1@�#�!�ی���$^9ō�Dd��׌���'���R���U{;�+��� �H��eP4+7���grv�=K�AJCX��������̱� ��1���-�Y�B�6�8��L��Pأr�-���PpSݗ"��0�	TRh�m����]A�2�m���t��)�7m0%�����#~N`FO��]���Q=�M�S�N���q�+���]K}:�g���"���4ԃ P�%��c-�d������ޘ��eA����;���J�YoY����Q�(%�vsJ���WZ�K#8Ϝq�S�M)&��(ΐ���V�E������R7�ӂ���j�UX8����a���i�%�Iya�b��i���Ek6�<J΂����m.�-h7y�^m�h��N�ܤ����E��r�m>�&�1�Э�>^�+�x�o��C�Ժ���
?qi2�De|�������O��� �ߺq��hh/)���;n(��||�������T�L����psJ̡>�o�0N�� U���3Ȥиz�[���E=c���ǣ�Yr:��g�X��=e�I���{�h]�B=��5��Ͻ5�u�}�b���
�5*"��(e~��o=��o�2�Uѡ�ã��H���:C���/3��uB�9!�>���UXwo$:Ģ]3&Y�@ �=x��I��AV�y�i$A�X����*�7MYu�v1�M��;m���H������ڥ�![�B��nd#B�����s�N��)7�{�UX�H������Op����jR��
�	'�������a����3;?��%��^�Ĉt(Ί�s���]?!~��~����e��*�>�3?`W�D0��Z+�}{׹Bm.�6�*�����B6�I՟y1�
`p�OI7�
!/�=��h@"k18dn�ЍVxR	���G=�u
0�Y��D��w�f�����6�b\����N�H�K"����[
/��c�<q�_"�}8�X
�-?чױ��(/8�94f�ڟ�,I�M�eN���5@�2/N��$�����t}?Q덟FZ+O�@�&9F�
pqGYgٻS��3U�J@݊�(�Ѐn��'41�l�!�x<Z����]�+2�l�3�}&�Qժ�$ي��ǁ�&A8�[1�#�j���B�+�9�� N��Z�D/W�iy.��/c�K�}�_�~h ��KapCw����=�����aG���xI �T��>���_�Y����n��'���s��&?��ӽ�>���!��ZRr�Do�܀u��Qd�~���,���b�e�kh�iR�r���x�O}O����M�+��3�������d+K�:��B�˹ ��#���` 9����.аe�q[�n���r�ydޭ��Ԅ�$:3M��n48�|5h ��N͗���%.I�~?LA\��=!�x���qs`d����Sf���{^ܿ��_D�;x��w@@K���2|qrx�GB���>�9i�GM�����;%��B's�0�����7OZ�����3��}����+k����QN���U�Y8�0>wNɺt�,M�c��c��-|g���>VЀnz̼�y�^�}!4��w��y/���*j|��0qyr�<+��;<���9�P�u� 2,��|K�0;�'#t�%[ds{�A��-� ��<m�&�4aJ_$z/!�/��l�9℟�^����c��96�*��.��nD#�I�>�u���=����-{\�A��%l�z]׫9Z�����=�Y�rzM����*:U��q��N2J7�
j����֔c���x�[��ǻ����^o�^�7�.Ƌ�f(�O�9qo���:�D�딩P��SD��l�?�������i�n὾�
_�X-�cgg�hȒ�m�~���wߌ�Bx�Wo^�����j��S��,��{�̂g��i*Us�9�!�J)"�|Ş)F��_a!���c��t&/����S�$�&տo�����U�b�Zt�CcK��;��1~	�k��9���(��f����Z�A� Ľ��T��5���w����m�=�-E�x��KX����}2�j��L�2�Ձ-��Q��3Œ� SOy,N�y��:���Scu��6)���F1�rmA�`#��QZ�� �\W��]جw�)HI�I�?Ҝ�Q�(�N:I�B4���+9E�҂��3r�����H6�%�]:�{�-&A?�ȼ�&C�-]���ѿR(@�c0^$!HĲK�Yw�g38��X�]l�"wI1��~�	�Z>(s�Y�o�G��lZ&z��ҤXV��9�o�G&�t�;�K@U�2G��r�31q���
�,���a���WV{�(ɡs)��C��3�Yz�%��?�1��~�ł��n��`��H��V��J%ٯ��GqԔp�)�x�~��_�U��סb�[u�g�L9�gH'>��@%��.�:&�6�8w��\�S�7~�>���眽��d�R���;4 ��ѷ�.9O�Kvb�G�H��o�'Γ+�ɼ��X��CK�	�L��'�P'U/h��B�^�+�G�T"jƎ��6�i���+N�6Q�ܼX�&� ᇥ'!2w3����K��َ-�)��x���?>��N��j�3Y:�^;>VU�5�%�e��qȶ��ɭq1��0�������l-�h��f3�d���OS-�}���U��I.,[�wQ}8��>{�cqcї���8�qt���3ALPA�)).,����6W�|�"B�1��ıc0h�{�d�cēe�k��E7�]�*����jv�����fа �-�v���U��f��~�[79.ع��רa��X�
��W�|� ��U� .`��|�n$F�n�A��?�_(q�� g�0�+G!��CNG�rRQ;^�X �����p�'
�L��Т?FO�0��4�0�i8z�n.s&p�^̄7�8Y��`@e������ ��.�^���*q�h�����Xxm���N�e�����1���\�YF�����*�	f׆'FRw2�2D�ӕ��=H/@gN��{n�#�TEz^\`�{��ܝ����sl
^%eR���X�Jµ��{<��|;̊��7�sV2z�l�CW�-��j�=��8�4X" �v�߄ȅ����ߎڬ)(�?�y�h}n�X[����#6��|i[,	D�2~ǰ�ǚ�8p����0Ud:y�_ o�}���:A\·WA�Àj���y_�Z��������M��]e�Mٜ(�>-���X������u��������'#έ/��_Wb�Kو��E���+PlQ�d�Ͽ���c��V��㋍價��z����o������P#�g��ig����[x�v��$�x�17ߴ������L��S+�y�܂�e�_�nDk5X��`�����x�$�?��eTD�i�ڱ*Y��z��;�o��T��x�F"�v�Gن�i�����,�2џ2�{���̫Qr�Z��O�G�0�D�@�h���)#��\�H�2|�)M�E]
�R��pGF������4�ʙ����_ǋb�Dy�6Xz�3,&u&�EX�Y�*�Z�1���*PύL���i/fI'��FRc>�x�R�wsT��6�2����@v��*�$���������f��JPgK�t ���!0��[��f&�w��}=H$�l}c�d��!{c}�v��C^�	t4@��p5 /��E�We�@ 2�nj�Jˢ��-&������y�M.}GS��%k�J,y�-��&��o�S7�b	Wm����{�Y�lrFǷIxɦ�hC�؅@�LCD��}��O�U�2!��%�\N9�*�d���h��h�
b+�&���AʾՀ<�Z(;@wTmG�G�O>��A��fC��S��8F̙3$�{��U����>!�MLj=u��֋qNZMf��8�M#"
a���
�LP�R�Rp @S�T��K���D��\q��㓤	j�0�D!��l��@4���j����8Q$EzI���t���c�$Ã�?��z?���.���8b���p��#h�Kb��J {�*����_c��n�����{J���f�N�]	Qs�����Ȝ��M�^�5�nA����,�X[����U��H���� �
�w�����@7S���F��s���UUb#���M#����ɮ�C=�����*R�$��PS��x���<��{��<�#��"��B?WTO�|�ǥ�؎�9�A�l$���5 ��s��0���!m��Fa�mm`V�}ܹ�<O0���e4Kf�p���@���[���zN�K%����=��B���Dnq���f{�z���l��z����E_�l��=�^h�h�d�A5֓`�\V�V-�=P�%�O�m�k�̷�:~�,
�Jʁ	�ir���3��ս]�1�{���lG�mO�d��e��+ũ��g��Xf�c�p3�1?vk�.�0������n�}��E����.GI<! �|i�G�F�@1���DK�$�!'a*��h]���r�\�m�U�*��9���#qv�	��3�6b��{w��0������!�G��:t\���_�J)���V}t�\jm`�����U�Z ^���9��t��R6�k����[�"r�a"��U6�;MS��������)��g �<"����#q���j�$(@Q�#�aAܰ2�SE��h�y��ݾSNC�IT:�LS�����=��X�E`7��7u,�t~=������1���_�1�?/�N�&�����]�0�!22 ��� �ħ eIӫ�hև&4��N�:vb��T��!���Y�c�0�ǻ��A ��E��T��|��[��+�w��A�.1|��d��Z�:���1�H���#�u���� �V����)�E'���r���K�d%�;{B� �vCs̽����ޠx�M)`'(������tk�r)8=��v�����.�A�AN=�_�S�j���F���9U˷�a��-�S�_�Z �3&YX���!��6;亿zaa��t�ԩCE���c���+ �s+��Gz?MFj�O����O���C-�5ۃ�c�䠄�+�1'%zy�j�xז2���D�x�#CitE+�����T#`_N��Y��M����4�`E%�=IJV�۪���������2��tl���q����*%�_m1��.U$RP����0�_}����l[�V�$�{�/���0UŨź"�b��������ǬV��,¸7r{��~s�"�	)#�.�����
��<��o�{���Ř�D����Yj�eVL-���+�Y�YG@��C�.�(0u�Q��S��_�q@3�	t��b}��u�y ��]�;�.�:���5�7�F��$"Kl9���>�p/��a�A~gV�׋�sɭ,�4��`�A`�5>1%�VƺM�.a���7g`����#��bJi�|��3��L�2��7�yUk):n����@����X9���L�xd�(�h{�R�6R~@�[�ʭ1���� �?�",<��I*~l�0oȐ��@�-��Y����7 ��l�>����Ē�k�\/-|�L��&8�����;q��=��/�.nէRC��bBޅ�~�ؕ�c��|�; ^a[�hR���r?R��Q�Q��~��&X�Kt[�s���y������vd/�-��Y��5���kZuڕhsL�'�SŞ:��1�Z�s(����#i�A^g���N�w��̓��z�r�`�y�A��-X�!׾�Qt\�L�_���otid�%><��}*>#w�h�7���Aٞ�R�p���(o�C��?�АX|�n��>�V ěK<��ɛ������&s�+Y=��ⵋЯ��`�Xԡ'ٟ��#0z1�b���y0&��ԑaN�f�JB2��_�x�w����ԃ=����b�opKwdM:�g�{�㶤����25YA�
~7ſ�6�9��p/���~uO�vj�h%ӅL��دiM����Ȳ�9�'}eBK	�l#Ć�5/m�����������GI����O�`�}���^�jU��s$�ʀ�*z�;�����a��V�w5V^�1q��8�f��z9p�?q���p�Ξ�@��q�֡;�G��&5A�ߏ��n}v1f�%�C�I��S�[S�	�YW�| �ǺH[�3���N
�eT���:�D<�;�5�o��G��xK�;/2RJF���.gF������nȑ`.�G����9S �,��N. �K��!o���)8֢@�^Ҹ6�5����	,���!��^��H%_�m����1��<�?��������]���Nbr`��<�&Y�M�i�ˈ$�vhut�ׯ��=[��Uw���^N��a��k�}K�����hG?\���O4'�ɪ1^*�����&-����F�f���
�/�~�F�+��k;�I�鳝��d������kFP��+ϒ;���(�M���:���Z������l��ms΃f9��
�~v�"�����|A�9�K�_\��@�WZHa��W�3�fҘ���?��36���c�dC^ �%�K��UA�6�Tb�)[m�iר�l�\��_r�u6�n�sѣi�����(r�[�z���gxk�8D�����J�_��L�� ^Q��N8oR����BO��2z��	�1n!I�N�f�O(����d�vOM�)��ͭ��͟��-;�V;i��.`$J�<��}
��ـ�!m�16�K�W�0.�C��:ЇB?�.po$��/��0NBx�t�wSbnJh�:�|~Yc�ҒVAxl� ��\�&���pL�2�ހ��݀�E$�F/5�A����眆���Ä2�B$J������y�0�XzȺpZG�Q�?	�G���7��@է �m��nw�jm]T�f�|Hü*�'�9B��L����������< C��
��<�(�"C��̂߰>����R���K�[�,���H��`��&
�3	����+V�oy��(��ǹ)"F��Sg�ռ p��ݑ�s�E�JIq�of�㶕�$��o�J�-���ֹ�}����cNSPi��}���9Q��i���5�N{�����1�p�ٝR����uS�%�'sc�xn�hـ[h쨑D���N���2D��e�2�S�<ǡ��8x��<�2z�`s����@5��jZy�J�:7����/�LF�?ts�7����_�yU�P�x`B��p���m���j���k�?�r+��}Y��,��C�;W+dt{E��sͧL�3c��#p�:��%
�ĸ�[�h0�e��n�(էD
��؟��Y��eF� +�K��z�Oc�uƒ�J^s��jϗ��c�爁���[ �|W��j�4�gd@�azE�Žn�Y�!��O���2Ӆ����A��h����4�Iʛq�3��<�A,*�-zHa<�$/�%�:��z�bk���	s��(G�$5�!nc�?'�!����t�a>bR���nS�rv�R g�^�aP�d���_k�q��$�����j�@�`pa�D
m����X��ם�ϥ���^ۀ�L�b�^n�G�Jھ���y􀀣�hVF��������w9\Q:�#�m������A�?��=�BY��2�R�tQt!����|�"x�C��3B/uAy��(���EMb1ms�q����v�����/�T���D܀��n$)��y8Q��f�������ݼ���e(�{����;˃�d�y0c�5߹���]_��@�
׈��ԛ2��C��%����X�.�tyH�G�V���ltA�^/�2���=��? �)>��B7��0�f �<�8�봇����v�
q`��T����/��4��oB�f�A��,�Uӽ��A�p�k��\��Kxv�ave�77�L��fߛݨ��1�h�(�8Ƀ{�T"��M�/��b3Ӛ��[�֎�H'�1R�_�����g���ٟ��a��%K0��������rF7��n��]�jU�U����n����ܚ��XuK��$ZN�`D���bOd�N�k�[@���9~�	�ψ�[���`++_z��L��oþm3љ�S��))�_i��a�	���R�e�6��Wk�6V={FP>�)l
���8l5�G	�z����ב|V7]�m�5���놑qTY���>|:(�����dM���*���ƣ����Q�v �E�q:6X@� �y���9Ҷ��cd��%e24�����2g�V7�r�RFgSC�+n֩�X �4ɺ����h=��'�������qN݋����%Q���w��(6}6��Ao�iZ}NWMM��hחb�:�t0����]2��ϣOG@�e�5�緳 k(j����Zx����3g������a�k��F�\���U�7̗�w�u!>���lh��S��E"�BWL���[ڬ�ɠ������F�0��_� Ds�S%JRPp�n��lc��*|�v��L\�}�M{qe.}-� QL��Ϡ��"�G��f�.�����Q�����g"��V��E#I]ds��'��)A�@T�pr1�3x�F7�>��4{���_Z�Sqढ��i��S�����s���\��q��n�Q�爯�,�=�^�x�K�+	#dIs�ͬ�����Wr�q ��x4`T�b�O�_^mj�R.4�����
�w�8LT=Er�d(ʅ��f�����c�fW'y���G��)���~'3dq5g�H�Zj�T��WPU$ђ~.���q쮍67���A����xIUBi��uu`�:�j���d���q�X�l)T�`�b6��z׿T�VA4�R�w�hd��`1�}�ɖ!ED,�is�n��` �� \+L�>�7E\kv��!��Ã�ּ���N�D(G�)JD�+	�>{dm���O�Ms����o>�"��y��Ȫ��(�P��J�1qL:��5�s7��y�������9\����e�.�o��]��A��ҟ��tp�=����"��>EN{��<ɋk$ߎgP&�F���9��[Y}����`�������27\tTml+��s��� 4����c��>��0V�b�!Q�,�q�m�X���s��k�}�\2�J�}c7z�ô�o"vL ؆57��aԆ�x����w?�;�9�j�M	�.��ժ���/r��.��Z�Ԡ�&�6}�<��>Za�@!�`nFeE�?�!:��e��~��S����Eyd_R8�%5�y�E�fFF��RXV3����m7�.³1θ�%mXt�.r����8Y�q�)����/�6��5#�F_#�o�I�x ��@��s��W*�Vx�bC�ђÔH}��WU�����-��Έ��U�$ԙ	��r�w8(������ݤ�ߎ�n��
������E`N3P1�w�}�(�k��n�S���&��(�=�q~�k��c�4������AR���'&%>��o�DR���*�GH	uU\ܐ�c��,s�;�.d���E�#��((D��?5���/�d�z�c�����.����,���N.b�t��'��D���YRQd��W�*wbC��>�0¤�n��)�{]�Hp;y�e��'���
�H�cK��o"H��i�w:QX�_/y�oD��j�h���rZ�:�EOEX!�F�7+����G��qɉK�PO�t����p0�<�ޱv��(�Ù/��(�r��乑��fg��(�h^�B�~}'*L�v�F?=�����d�T�I ��}俚�_��)�^�d۵O��R���F�z�*���t���;��4	�yܿ���}��x��p�ؾ����qޖ��ʽ|撓> �aK�O�-�؂���4)o�c��!��Ѕ�����q,A?vN�/s����~���-"� U����\ԛ�g<8��|g[�ф�9V��49���T���̤������}���q{ҝ��o�^<rJ�-6@ܠ�8�P,��A�{���#&$��KH���m���"M?d�ۥ��BȋuU��m�'�&�/�J����c`'�����F/L�z~�ݹ���h�u��n[M�k{I'ݓ6�H�,T�U�%��Q����M	�%������:�)�Z���3��,�Ѳ�٢��Q���H�2ëI�d�+8����}A���-ܽ��rA5ס��;B=o��>'�?�y�'f�-ㆺ���\e��B(��"�>�J~���2-�.�B�[��pCs�oP�?��1W9$,}��Cd����y��Ad
��jPw�~���f�� ^�zj�;��#��a%>�Qs���_B^y�igي=��I���9k��m�ǈ�@��g�7�+�ȿ���-<��%�c���4T�&�$rAG��:�؀�vZ�r>�J)���y�� ��Jq���$����Dgꚝ�����|4&�B���0,� �>Q� �;!��n�cU�#�"یd!L�ɰ�'�5���� D@G������&?=�(Z�,r:_f'� V��kJ�r{�5�N�v,}0�����������hR�2�Hle�g�_4��L;�5S�P�w�x���Tb۟Mw uqf�� '�+�M��x���-^�Q�۱J�TEWVCJŶ��'�,J����P���M��Zor�zإ~�`�H�%gķf����㿸���P���i��\9	+��q�@�
�eI^��v �z��Xp�)��[xA����1�A����-�Άw듾kǞ�P�vq&
 LA5���~`8s��x�}#���y#�ʝ�)�i<D���9kG�&�����L��w�8�빷I����P�+����.ZH]3��3ŹG/Ϸ�_jL��E�U��M"T�X�,�:v��l�"u)	t�[R�y�	="�S�>� >!T�R������5y�a��W��h�$������j���9�#����B��f��<�u=�R
�Vŭ⬜H���}"���r�WU�]�`�����<w)ۧ�ueWd�j#�A�ڒue�@�*g��=ǰ��Z��R��±$9|kٗUyП�Ar��b�eAth�� �qg��`ĳ�V��d�l�u��,#Fs��&+-��M?{�:ɵP�FT��9#W�n;lx�˸����w)Ih���~	�P#����O�0)� �\R���aǛ}Ne��;�G����z�Z�W�2L&90�qW���w��	�G�k�?ע�n�Y���ۅ˳�C���p���P���ċ< ;���k�^5$�_�g�c��}G���%N��]��36U;�R�Bc���9_#��D�4�^iw�(y:3��5�Z���c��P�F�������A-���.�������ġQaR����֓G��#i �v]�C�d��P���E0ܔ�\�֗Z���U�����^;�Ή<p@�sd!�R �Ȅ��卋��H�J��9�'�tbye4�~�Kw^,S��M�?i���#�R�g�(uh�V��'uD�D�}֟��[*��j�,z���w]����*Lrk���#�Q����sX��4p=�D㋩tc��FH���?C������x�������W���T��z��O�����4�U��Z �w�A���=��ĉ�`.�ۓ?F�n]>�1�/�ޑ�c�)�e��b�fvĢN����#��_�Z=�;	�k����d○���m��&?X#�4B	N�L�F���b.@��lR)��0�
��[�ۅ�(�sXA�m"Sf��#3���Ԁ\�Z]����cO��
�D��w��{�m��/4Pj�����ۣ������Y���l �^N+]#!��i�uW��x��y�#�5�ކ��cԷ�.����l�em��K�����͔��| �ϓ-�#۸�Nąa]�E���&���Qd���o e�}�(�E>h	�[�"�>y�^��F��NL�(�*p�+����@�bJ�)�R���� G	5�޹d�-6g�n\w�sCM��o�Ľ�b.�>���C8w��n3�MU2�ʶ$.��c��;��۳U���T�t,U�Q)؃�h��������Ew{���4�nF	#%6��׊םs�O�����N�7kS⳥��h�w[�0��|�#s��.Ь�4(�`-�S���"Y���s��Z���"��?��{q���`�KM�����("m�V�\���Q��g��e��)�QoyMV��v#�W�a): �d&0�D�,�p���g�*�W��E�(�(T/��f��?��Z����L̊�tυn$$�m�x��(A��0���=;T%�2Bb���l�[��$��I^/�֮`c�՜>By�A9l����^�!A�vK��X������N���d�EK&�l9�}t���G���4��еO��1�'�w�`
:~�jp�x�"�����/��OG8�^,JF���`��A,�d�k���r����] $c_Y���ۏ��
����g'z��L꓎(����c��a��0v���Q�B\#d ՗3�:�e�>���$vV��H�c@k�bC�B����|�S��+Z1�c�xX�M��>���~��e��,2g-��2h^�I~�ϜS6��v���1\����E�&]��챌�����Q��6@��J��k�ȕ�DUc��7�OE�ח�,69G)���<=�.R�f�2�c�G��A�w��#��V�~���ŏR��ׁ������:������C���)�,
\^��i�Bl%�3� RRG�����:}[$w��΍?��������5JA��yǗ[#8��F}Q��,�i��y��-�7s �)^�{�n�M�:��s�Ga 2���/�"�8����ۇ�F��3({��
����Z�����KC�{���4����Y��ǣ��O��,9�m��G�97���HE���!�Hb�ޒ�����&}�LX��^U����-�>��+`k��������n_�����T|���U���5���VG:���m�~Iz��n����Y��aث����"�aU6|7h=ҹ�.�2����&[g,	��{W��w���AF�<B��8�9�(����R[M/��e��X�qg5����KU��TY9��������Fo���)�:�_���� �o�1���jBA���?����\�ޠ{Ǚ��A5F�J!ہXݨ ���f*Q���JW�~+�(���\(��d�`E���je��Ea*�L�O��|���3��ka@�a:s�0P߯Ө���Zl�hq�r��&-h|u����N)��f��1o�$
qm��
�]�����s���{�g�����o��g�}p���a�m;$��
1���P�	�o.NLgx�����Ar��'�9{k	m"X�P�z��qi�^�dBA_�|�Q��}��n\��$��F�������LC��.�v|��* �fȳ�'f�R�Dܥ
�(�4�m�-�8N�x���j �=m@�� *⠩�}x���%z���H�����RW��6��mrN�(k�D����m�W�BC�9�ٶAԽҜ���O_g������T��@^�,F־+\�W�yq�"���C��N43�߾��p4�&�L��XCw؁,�����ލ~�JQ]�#����s%ea�w����^DZ �f<�����U$nw�pɧ�|Pi�ʺ�kó<��o1��a���qS��b���F`,��=����3̷l#BwZ�+3h2H����:�Px��� }س�m5$�to��'!�d�R#��b9���af�?I|!����-yb�[%:\��W8��R�FK�����+��_�vƐ��`�I߭p�w3d�<s0��#����˱�9���۹\ʹZ�ٳ��s����$u=ղA�����*	`��i���Sϼ�]6��$��\Xq�e�6
-��$�z.��I�}��ºH����.F��a�Z̋�7i��U�ĠU}eEU��O�L�a������G��lb�AKt��Q	L�󩖐 �<vhif�ۻ�t�R��#�q�x�D��ca2#y5E���%�_���е3�<��n�Q�PZ�U���]�?7��ZL�,C8��1$��FA��oʖbN�oKѫ��� ���A+w��,	|�|	��z��5�Q�	ȿ�Sȱ!uX2���G�tkS��G����{ն��.�Ƭ�F�\���[�2�vz���c#vh���u�=�Ό�����-]��z�~�Sz��?����U<�n!G�'�T��������B�@��߄���`�Bh�{�Q8�'�2�#��s���������C��-7���!eN��w$��m�#��~��2�=���H0q��C�L��/�+��DfdLd�3���WR�	�gGL�>f�)���Q�q5�~r<b9�*pF3a՛��K:i�0��%��Ǒ{���
{TyYW�Ϩ���b�k\��8 ��O�(��[�}��
4����
��9�&��;⃶�m��cpJ�� k�'���B[��>5k;��/�R��7yP(	-��&�Ԛ:�<J�1�Y�}�1$1�W�f�U�(~C�j��_sz��	�����=G��E�؊���O/}���5(C��]����]kp6'���;� Q�	��5ޚ���U��	1���b���?��߬�d���B$z��w�6h8�����'lR��TP����ںи=�t-J�<�����w��xo�5 �m�����a�.�������h*`>�g����D�dp�@�>�x�c����QQ�<��k�ԙtR2���`_����+.pkh?�Ëm��)��֑����Aʯ��B����<����T0_<�d|����	��j�Q�n���	9��L9#�P�
�)s�����������=ylbdZ��Ol��:��`�b!� �r,�����0XPQ7G�5�k���\< 1���a�)���}Ē7���J>������s�-��G&�1�F�~B���QR����E�/��+�9�k���7��ny��/3Z�V�����D趋�q�<�YS��B���%�A]���;��3�@�[��M��y�_��v�8��E�_l2�)��,E&�=�B=]:�{��E�ɹ��0Wݴ�eoq@l��C_�;��tI�x.w�CkZ
uğg(�M�4��b�H�m���1񫀓�>���%�6%��*���fh"1 ����������a�Z�_��s�:�3���+��� �{�F� ��*���`�/EB]_�y;x��{���E��Ԋ�hG1�������.$�S�;�H�H"H��{��J$�o*%�>���I�e\�c��?�+�e��$�1a<ևpZGa�I��М�.��E�������l��l��݀�~����陚(Tn��Ƚ��Уۚ�a�w�C�L0����$� ����"nzo��~4�6tw/����a-��ӎ!���J�[&T�D4J����>�wa��6��,c�W�����Q%���[7���U�v���Է~ �\�k��t��V�n�t�Q�0�:<�w0[_ P. �����v˫D,O�Mێ��V��35�	�-�,\���:�q�c��*�##��/��mhI��7���{��߄�� 4g�9`5]��`���@�yl�.�C0[�>���礂�u�(MЭ,<�1�QfVj��j�E�����-��N�V�^��D���$$r�*|�\#�.8�iYr۱�)[�� "�a#�:^����&���}��`�M�m���t�҅�=�ֆ��#����(���%������V�i}�]{����:�?��p�r9��Bjw��'�*X:~�t���2���7�8�PP-dw�P����L��F'���I��?\������Z/����ѭ�m�ר�;��H���To��y �����N9�}C����R�� ��JM�y����~`�j�1K��S�\������l�WS��4��t�ֺ���I��*,f#��d����R����0=�zB�k����t|���9�G��@/-�*�&�Q�T�zV�w�V?��~䛥�$0�=A�*J�^8�.�0yzS���	�Ms��i����91+/��?��"�L7ciyH�b2�����BO4�Jm��ǧ���|\�m�S����뉑�-�fI�K��� ����o��<���D=vO��e��i��M�$"h�����9!0�����������<�W�)-	�5OAZ*�N�K��AZ2m�'{���Ŭ�� ���eo�ȵU���q�Aʥ���2��(�9k��!A>�;�-sn��<�z/��<�w��;k$uꚈ����I״���w6�x�@)g�a��h����~�v1{���X��Ks�X}�z�^����1�g������\x):ٟp��s�(�b \�Na=�JyϕS\l�4��/���zΟ��pĒ}d�j��u<��a�'�5e��in�9�
V�0�u����f��՝JfF�7�.):cԟ?�qyH�����YW�)�m����{ �1䞤ʂ� c���`j�\�����Rb]rt��Vȁ��F���K�IN�?���~�*���<�����M̍����s�hr�i�]�a��)�!?��[�Q&k�hp�]r��j�ɉ���揉�_UWJψi���w��5���c�'�oOp��>?�6�?ݺˬ�6~R�4χB��R9i�]D��l\Z)<��NQG���SZ�J���C���n�^XIx��`��;)sH�8|G�Y��/������!��m"����vy<sQ�-�^��U^_J�����z�$���Ќ���Z��:�Zi�s�$jP��D.'�`��*�Z`�¦�*t�[�lE��T�&���7��ScM�D�M�fI=�1�Ô�m!�8�4�I�[Ƭ�4@������N����`xqKoL�dAڱ�(�V|d��x�L��͟��������1���y6�������D�^aY��/�j����=\2G�g=(N���#
�����/+x���c6�')؟��_��r[J�N�."�Q�7�ն�jy������,�魍,nUô;���Xomf&����b5�K9����@��.�0�j����:����;��CE�A#~;����-���y`�А���Ewͺ란g�W7_W����pu�ʬ��59g�(c����OH0���A�D����S��B����dőK��!��?���y/���S_�
F���z�)�m@��ml÷ |�F�C�O�N�[.Ȧ��ȸiY��D�^�4 ;k:��ײ��NN��vH��p�/[G.q�,��b� ^M<&����+�
'y
�2��y��z�"�*<�f.G~Nf�����ޕ�5	Q!܈A�G�iul���T���)�v����E+>���24���v���=��mޯ���yշhQ<�+O%���0/dްFz�v�8�O*���G�Ng�.�=�D�t��`��R��䥦K0�tP���e@ε�.��~\���g����|	E&�eoi(��>VVm`g��W��o��jC�]}�Jc�ns��SF�������½D8�����IÝ�����nL-��bS�ړ��z>�dP��/���N��(�fE�s���xȤZ��1����r�?�I	��3��6$�Ovw}�gY &�����(�M���a�&{űa�hZ=V�'���J���?0��?�Q�lIds�T��lҘنI3,Q�<1�N�����C��I����nc�53] C�4�8��y��]���R� ��{V�\ DN����. �k�6n�f����@�A�7�S�k��yH��ce�98d��Za�G�Ӗj/<nO�4�Q��W�h�� �y��"�$�``�����.��Â��K���,�~Z`����k���OH� �ڸ!�8a�|
�}d����"���e4�e]n�$f8�
*h��܈!�q`b���4��I����ź�L�E%�A�Xi[����J�9&<�O��s
Ô}'�d1�3�X.�C5	���������Da*�-����c�Hw��C.��ӎ�s�ORu���[���Z���'�"�T@-ݔ�<��9vW��Ln�e�X�F{b�K
!d�W�ұ/���j'�݂?�*)S�"�����8@
{����734(�D/��j_X^��D���Y��	��_
��"�2�z���rq��xh��D��5`�CW쾖+H20O��$`��@9��,�8��\2�/ivU�
p�Ci�����"A�I��]��w��ɼ%v�N\����U*G�zo˵r3��&#�.���7���{d���,#W3Y�f���\?�I��M��U_��.�hTQ�'
&��f��+��^}�G}uA�tj�oW2�9�*�(pM�){��b\z���1�]��\��9"�����cW�~�)`�ⅥiD��4�I���q�U�2��s�WPiX}tEڿB�D��/4O��M��s�ytVmz��R	g�?��D��F��Mt�ꐆl#h6g��f 	�KTW���w��:�,�_o��Z��АF�9C�%	�̘	�/���'"9����+��*��J�@0l���7�Ⱏ֓�8��J��jYʛl҆��&&i��m�+�2�	�{�-����7Il����p�?*E)0�rXH�T�`��U�S��E#�(7���WгOe;�������-�PF&�����3�E�4gn
�"��@v���S��m!�'��:�-�z��W�;�:�P�3���N�Me��D=�(%��JXx7�Y�$�&��!��n�,�y��t��\����k�/���H��9P������t �¼)�o�>���9����2�Vb��e�Fr,o^"7\��A��7|����,����?����:���oc1�u��V�}�;T��܋U��sݖvψ�����9N�Fa���-i���
Yv�S�����wd���6���y�<d��r�O����٭�0,l��]uN���2���˾bcg��=8r_wF/�D�^Ev��L��t�d�S�bU���V
���5�&���e^Ϫ��6�b��<ҍ�<�5a>!��X���&u�$�]�-O��3
��ʣ��V��j��c��P.U�l���xk-�Ԣ��m���8�alټw��{�@�-b��u�ëc�?�3D-�{d�)��ȣ�I#i�ea��.L^�&˶����ˈ4[\���-5�#@���$δ���Z��+�T���w�Ң'"�{�̠�ҫMx�����6\����-��}Tkq�i�wW��� �!�i�p2�c{�~���l���s�vXS�=[�u��_h��G�~��-y��EC���"Ռ�鶗*����_�M;�1n�%͙�睌`�K�ն9;XC-�%J�tS�Z�2�Y���(A24�}��.愥��Q;=#��V*��a�-�e.e�n�8�o��kL�T�o�u�Ɯ���E�x,�
�� k���H*B&�#^ �ҏ����l�-�¤K�C?���_���a)���fX���v�6�@0t�S,����I��M9&v��������uo����X`�WH�oij�0F�k/+�S{`��
���7e(t7��,A_��?K�<��2�|�a�O�n�.�u�	hpU�_�쐴߈���]	� ��CoZ\��O����H�/�R%aQ'��ĩ5��	���Q�6~�B.U��Z3M0�O]�/I��6��(?���ޜ�1h73D9��@bZn�P�8bN1�
�}�DS�D�����z��J��px�w��^\l��fb�Iz2 �rW��#������ �(WןU|#�	hND�?�)�k9ʽi���c?��R맚e��Y=�.��^q�Ĝk���~�g#a13�����I�/�н�����3K��i�UnJr/�hl
��UΞ��d�g�TV��-�$S IV̯OB_���������W������(�Y�)N�߶d�����d�yT�9�4ţ���B{]o��_��ԣn+�8F8r2�,El+[u�@&aD���jo$o��%�/7۝Ԭ��j�0�$�/+I�Í�ɛ�M-�ǹ4�W:�����a�f`˅�w���=���k.K*M�X�=Xa]�����T�����3$X�vE�?���sX� �|#��rS�i�Y�ҙ�����d�� �Y ���#�E�d&�^'ą3�Ţ�+A-����,9���/&��]c���]P]�(���}�|�ׂ��x�k�AԻ�����|.&� zPx��
�m��Č��B�e���3�{X������]b
��#HQ8��I7U�H� ���l)���>�0��w���x��bW ��#��zQN�gr�;�m�gų�_\����LT�E��{��F(�I>�H\�6�b�3}��g��EJ7�K��84+
�_w�����\�8*��d.|ֲ���Zln~��fh�S���+�+�,{nyC�G�Z��Q���{���e�K\Pn;C+��w��	(���3���^V�aP�W�Fy����E�C�K|�GEɣ�3H�g��iq.���5�#|��eı�#�*������;z���������W�2��F�K��t�Ba�	���.Y��*��m/;0C���*�9�� �+�eB]&��٤-�������_�Sޝ�1�P��z��a�����W��qx'�a��p׈�Gk�Dq�BY�
.��L ��tVn�p��ܘc��2J ����J�7�#R�Pl�|��~��ps��t�5
4�T�b����Q�2�;�TmWs�jX�dj��:�@5�g�/*�4l1��RU�h���M����TR���Lz�!j^��(P�?�W�N+�$�c,$���!Hy	�x�A#�1�vC�x&"�������	Cc�Yǥ�$v��DJ�f����ཧ�Z���:�q$`�JـF��'���[�������E��5Qw�)�^/0�|�gq$��B?R��p���a�-�y랔�����8��@�ɝ��c�F���-���d��Uhi<�[0��2�u^Η�)wG��z��ڂ��pTl��$�tѻ�d%�p%9�,�,usPX ��vX~�{�f�?�p��t�����Av^nI���7`��R����	e3w�H���.�*���V��QD�Ὠ������C��bC��Fu�ndY�D���-��I�����+�5_p�d5��R2X?��g���N�t��h6w���4�J�x&_��Y0�,���HI����/Kv��q	E�efk�r��yZ��Mw��"��~0<��=z�Ytm�Eu�^vO6�wk*�rY5� ��o\���@�99we�)�9�bo�<�=3�D�y��;nj�6-`,%�w���,�+jA�wˌh����)up�
���!;�)��)
�˺s��s��nG�t�؆�A�.R�Sd$��Y{�yE$pJ�g҈4X�K�U��0u�薼>y�+7Y�P���3�xV$�3�}[�YE��@�
,]͔;c̹��.Lz�s1��0G�8Y���U(� S���5�u�`ĀЛ�d��)x?G�3�� e�D�r��KGv�Co@�N��x�jJ�U\���*�VV��.��h+ЄL�~n��B�^T���}��*Yd�7���w]}�/���z����M�)&!G�8=B���u��i-�\�()�=��)��en*War�{������$Q�x�/���dA�*b��h�?[�� Mހ�q�ݔt6�n�����nbX���7��|7bK5��t���I֊AŪ�`~��4�|���̀ �dBï�Q�#a��6��1�q�I|7.�%|�3_.�Ӹ�w�\%�p)\*��+Y���L8�g��](����g Xv���ȅ@8��E��r�^v0�@�l��,�uj'6�E�ثF�Qq~ޱ^�����y�M���s�0�1�B��E�,7���!e�X�bhڴ���o��g ��1�7�_L$޺�破'OB6T\�C��
��\_�����ۼ.�����a4��� 7R��E&#��DetlU���%��K]�����ߞ���As�'mW!Z���_��=���S`��f�� 8��B����yΔ�"��E�VeB��#��F;m�)Y��p��=�o�E��FS��c�A�����V�����@�Ӆ���8����Έ5�7��x���ڥ�T�x]���頫���9���aFÕORA��>1`c�ò��}�u�t5�"��J���mW��	�@�نH�'��1��|�p`�K�Q���CNn����;<���n��x��I�>���cP�p��t1�.�A� ��!$���\鿘�(�E���Px(�����Ǳ��������� ����MѩF���P7���H�ݝ���_�:�"z��涓����̟1�=����m}Qt�#T��:Hj%C�I}X����Gr�o�����(������::�E���0s�[ا.���i1קC��0��-m��>�{�Ȋ��.�9&Y�xkt�HZl���)K��wM��(B-�zډE�℥j���À��?d��Be
Y�W9��*�;�So�|0T�i#R�5gl���1���QT�}��}�d�dO�/-�X "�5nsoR����H!�Jk��%r.�n͵$�?Ds�F�����f@ ͮs��W(ႻlG'Gߡ�8���LvfR@��0�B�1>����r߷��t�e��y�<[�f�$��ّf5v\��N����;��"�|Jx��z���96��D��]$������VcՄ�9|��C��uz��ׁo��Ϥ!��|��G?��"��O�<br�@�C�[��.���N8G�i<�����.��(poUm�-b�V�����_�TD����	NĆnMۣ���/#��օ������mJu��]�u`��aa�5?�����$G�R��x�k3j���|�ٕÿPs^�>�փب=�RP��)��"�;E�&cH�.������E���1�Jg�}��/��8�����h��!}��Oy�w��	��*�V��燖b9"�.c-)_�v�Y�<'K�mD)'v�I�% �3^Z���ӛB���hM�"Hf��o�a=����	���"�lc]d"����{T�܇�J�l�l���ӪU>7O:��Q
�D�Yj��I)��#��x�*��uc�X�6� ��/t��Z�2%6Z�8�v� B�!|7!XT�<Xq�
���d�]_���m��rV�����:
�usG�s繌�,"���[Sv�6U�� h��<l�5��@��t��	
u)����n�2�+R��؀k�X��r�6�Q2'#����Gl3���wEcyd�T���bs�vRy6:�!���!�8�k7���>��6.7�\t3�A+���G@K(�Q
�� ���������ɕ�Z:WT�^��y�ů�9�V�h[��	%r��ac.Q�xm�x��KA$"�(O�:�1��&j�LP%��o�o�ewe�������8�TX��zhѳ�X�C3���=10HN�.G'R��/RLZx�3ɺ�)k�����{�%f�V���2�s�x�\�>�&�q3��Z��<�i� ��Y�z��Y�N�Y}W���h�G���𻢩T��*�
�΂��el+C���t4�"I6aE�G~��I-&��x���[[�����>��wd+������g�Y�!&��V��>�'��m�l}��������&����PR��,��VǕ��X%�,�����!�,�]��q���^����9��|¬Y�7ƭ�y�?]���+��ש�4e� ��	eZ�@�c�NZ �4������[�8D�@��В�6�\y�>�R��Y:���?*�W �	+�m\�T���+�u�B�T������7ܨ�!����B
�K��ʋ��+��F�9����g:����U9QҳV4+l@��+P��"x�>`t?��p���<�;s�6~��06���-������w����7�>��C��;[�BI	Q��_�Ч�(��S]ca��^��)����g�|�U���?�oE[m�0�rm(� ~y��\�����/4}�J���Yw��C`���ăȧ�"}�f��G�Q�ٳ��]ӭ�uդjq��B^ �\����pj�>�a�s��{�M�F�(I:Qj�m�5]<�0s�~&X�<sp��<K�_�"9tD�In������&-s��������n��{�K���E�@J���\%䲝@'@�Ky�y�J����e90�>�� |�b��p����h�o��0�@H���-.y]��
^��T]ݭ��1u�eM�Ԛ�I��u
Bo#8h�� S��[++\U�/�]`픅B��w��:o|k0?R�bd[�@��za|c�L6��86Vɓ����`}�&qD2������ώ����c6?��U�zD�]�	���$��=�U����h�m7qQ�m��;��?UX$�&��� 6��~�L���D�|�!���_��<R&�#�.r_� ,���p92;�e�KPj� 2��HCQ����0�FŘ�+2�FI�S�}�lLJ��&�>'!�Z"/���:�]�r�	z��(�W��.$"��)%��&3������j%ag��ڭP0�ԏ{�(��L򥘒m�6H��e�0��ܙ�U����Ÿ�?����ӊ����.��|U
��X<n�Nw�ޅ���=Ćd�^�-S:��T_�������-�a�x6`%"/��\�*�gQ�z�f�vT&��@�*7'HC�n���g��n0�e�n�`]V�����Bd&Wp������в�Ÿ�c�7�3gT�n��j�(ц
�����g����W�jG���e�o�o�)�F�>�9�-�bz!����
Z��f��۴����\E;�_���C�������B������Z�*z�ۈ��I&,�4���;��4���U�f��׵g�2��_�ל߿a��at}�2=� ��zs����������:������	bm�G|�Ѻ3mk8ࠦ��粈6��!�i��ڥ��?��A$��OW*�����duυ�\�N|�	��:%by�!)������"��x�\��� 0�{EV�類�:�-w�.�얲n!AZ>���#��#S9G� 6bP�\
K`m�b�S�m)hmy,����3՟wV�::�²��+�K>m�*͕/é�*��Lvńl��k���
�CR���Ƭ�R���F����H��V~��7m��6]�('��ڜ�� /�����}D�7.��H�I�P�F� ~g[��W'�H��Z�?a�
��-!|����2ZI�T�뵾���2��Oa<���E���ު���q�0G|�(�b1�?z�^��@�0 ���!I�Fm1����۷6�eX
�L�݄������t�V`��!D4ʚ��7���\�\n�Gm��}��:�9�������~��˷?]d)/�KB-�uﲯɮ9�^zw�6�UG)@5�?�Eb��~��3M��U^�K��]J�\+y\�N�_�e��Q���t���eF_[0n5i�D5����Bx9���:?�	z|�\͓!o�b��G^qhL��o�}iG*��^8���
��6m�8�qO�T{��$�t��D��,�ŷ�_�Y�����8q��K��JaZ�r�L�q�rY1�n�7��˨�p&�\�|(��Z��r��5�tޒ/Բ�Z��Ba�D���v!ho�Vum¡�J��U� �9�*����nFw�xb%��ܬe�Ϯ� y�YC��a*n���uV+�P���I��&����A���c>���˺�o�OBwL��v?|3��m�a�g��7��Q�Q�|�
�k�]X��^"~��2�e_ ��C��v|;�n��0TI4��s��4I_�����%5�*1L6��P��E���~�R��,��]3�58�{i��Zz��V���B�a]�����{ԀO܏r� ��-5�fG�\Y&����+0��b���Џ�����M��:������p�N1~=g��̮�s^Y����F�Z�"�@�}�L��ѹ�tFu_gҡ��L(k��Z���[����j�u�x�./���B缑�i* ;�:;��B)COT7�c�r.�h#1�W������x�O�r�?��"�*���fQ�ͳ:��*Ы����l�xu�;
/�a�e���/W���a�0$H�@��(�D^^WK�vA&�IA�tK�nt��P
h0g�ˈ������c��~�%���S�$�*�ź���N��i��Y2J0��?�x���}s)��M5s5R�$uEK��<gq���1&���]~��������m�g�DMG~�ņj��fK:��7�u�"���-T^����nE�C	� �|[�s^r��c��W��,����te��)I�A7�wl�ǔ2�3��̽N>��E8,�| ��$���	�;��2�Y��=T�{�����.ν�f\w
}�ƱJ'�:d~�����b�|Q�"�R^���"��.��.�hT���C�bo�����ӿ%{��>r�4#�e�S�j�O�4^2iP b�u�Q���H~h>�~�ז-�1��O��}�mV��^Km�@`�)t��� RvH*���B^�'�ڷ��z�� ���k���zqQ�X8�A!�I#���W0l?���G��/���zߗ��}FhD�7!Yc�c��o�c�:8�]ʄ1-i2c���>:iS���=��V�:�r��#Qx��w(��"D��L�zj���&����i��� ��a�f9�ƻ��f���o��:�㜓8�r:8�3�mbMbaUB![{`����1���?2����'߷ȻQ�/ˢ@�,�Љi �@@���A��tA,(S�	�D�����F+���6Ŷ���AT�������j
��5�ܡ�pkٹ�?q\�Q���z6���qtJ�s�\�qS�YS���u;��
��%Y��\Nv�D�W��������΂ش
�b�~i?�Rߕ��J�nU'�n[���XQ)G��e�w���ܤ��aoD�8K^*��D��Ȱ\Uq�g����:�:�.wH]��KM�}I0��mz^ǆ���J��%b�Uw����55���x)�s@Pխ���L>��`YN	����T`�Np��B�c�����pjeKzic��J�tMD�a	J5l�YdI�5����R����O�镇���:���&�R�I2:�e�+��/�e6��C	*7B=C�����kv5c�Ӷ�D��vL�J�Y�sn6�k�kW��@�-P]�f�}j6Z����1?G|��wA=�C�v���R�í�m 7Ch��-��J]�dQ�j���tJD׷�ѽ���fBj_�.J��}ؓYC8�W�?�H�s�����2@�L �Mj�\R� P[k%�����t�"Hh)����]��Y��\` YTY׉�7�Ck�8�m�g�����`ǜ�Es��Q*=�����./@���p+&ô
r�X�A��uB!�u��h�ΫB2U��"β������]��?V�)���t��va���*�)�V�|�t�lwy��.�`��jS�m$8���V��:�8ۈ-��2�{��.+a*>5�7R<I2���zPa�bںx�v��6oi�m�]
m�.�o]���0D?y6�'�!D3��-J#��%����y} 蘺z�!:�OՎ��+=D�ұs�������i
D�Ͳ=���|4�$z}�&���.����6.5z��ˠ��c��pL�I�5���S�.���x%�<����������w�d�N޸��R	D`^������%�AXa-�D1�>�ŚFv��6rsǾ��{ʏXbD\w|	�Ը��-77�eW,�+� ����.�tЌ�՞�����LK�i��1��4"9'��������|��� M%��)�NJQr>���Z�?X뮨T��.q<��
�Oȧ���]c{����¶��~3�C��	�.��F䀅a��p�G�j�"�����eM�^QV�tGQ�����v��n�ĉ1�F������j�����!\�b((
W3m�t�1�/k��@����/�/�� �5/�Q��$�ĭ�/v��XK��a����o�g����4:E9���DՕ�|+�Yv5'p@��f��pd�|�1���Y�:>'���}���Ag�~�x�gAiE�
;��}@��-I�x�Ht��B�/~+��p�V��J�K�{WVV?�$���{X3|�}�Dm��i1\d�Z�~���>���n+�"�t^��ؤe ����P=Al� ��O�%<�:6�0x�fi�Ar�Ee�V�����=Fz]��Ajf��Y.}j���`�	R�3$�����Pm�SC/���=�"��6B*��N��8��_�*�|�y^��M戋�]azj����eὌ��V'���C֟�dAލԣM��x��W��N� �P��èU�da��PNKv�Ι8�U:�P�;i�ő�)���{P�3�} X�9��Tֿ���z�e| ��� jN�^	���U�蘀���L���cb�Ưm!8�������J}y6��|�K@.�a��`��V������	�Oy◢S��>��?�N��������hpDk	�6�
t��������kK3��рxO9SBej4�M	���X5}&`���eZfx!?跃�vC���Ɯ�0r���[m���m �HY�S�Y
q�=%#At*�fMk~.��Z��c��p���0���L��m�D�x���Od��L4l�BA�g'���'t��r�+�t���#�d
�ߵ�&S�?W%�&�����%	1f����,�pIR%]�����9)f��}F���|�,�D�36�2Dj�B� 6p�>&�6A=� ����}��-ϑu?F�N�퉥_��������C��D�
���Z�T��ݘ�}x�6��'o!d��l[��]��\��q�E�)��eU@�a��fR-x�9�l+_��ş�YN��n���{��1�?��+&/"_،�����K:TMu��_u�,$(������AvsG���mEW�W���?��*".Ӷ.{��	�<6��{�B��@�[���]�G\粙��1z�1w�{�O��ǻ8��pV�^a����Ӽ\j��a�z,^�d��_�a��"M �\��䁉��xĘ�FGx^p�E�Z�:?2�q�u%�\N�6\��ȠE��������g����%Q����R��dx`���� ���4r7N�x=��c��ސ<4:>c��2�µ+��q^K��h�R��۷C��ٙ���Ŝ�&$dE�P�m>�ssV  ��b�x�wi�ZY'����Ld�ޣv귀z"P���P�G��=������@�L����@@��+pn<Ǌ�+ʌ]�����y��
>oV8?&����ćM�b$�R�<�(���/��zŅjs!�n�g��d�?��a�
��A�p�2V�&�x/`X��>)��hnY��w����g����wuD�D�{,|o>�i2L�j�Ύ�m��Tc��:�ӹ>�dF�-�g5�+M�rn�cM&�niXݷ��҆���Ꮆ� ?11�2<B�j�yv�hS�>��� ��J5����hr�T�sK�=���1�T���u�jj��Nz�d��hm��
s���%�M3��k	dk�g;;��,�	w3�*X����v���5�36ҹ���l��<pkᑘd�jA���q���*����%ȩ���-�&�wk�x��iԡͨ�N�c�}|q�9`�'�p*b�wxw�WRS�����R�;��1��d�WmlJ>�s�)�!���eз�N^�x��~��/�
�E���s�86)�X(�*�� 7�iz��7�VCO���et��3��q��{�NxwD�����AM��T�j��Swx&b����!K
���7�;�,Q���Ɖ��:�ͮ1EI�F�h��P�x����i�h�T4�D�^���5�A����
g!׭�7���Ά��w��k<���gը��!�!��|b��
��cM���LS���`�z�W86���Qt��&�]]IJ�G�P��H�eXr�xw�C��7i=MѬ�yC��אK��cvH�A��#�n���:BU,0�t������~U����#B�}��~�FJ���d��kL���׮Cg����J��Q�����P�=�!��X��'��D��i֪O��L8�e(�:5��4;���zN1R��T��>9�:���Uֽ���pwI�1�ҁ��=٢�+�
�jF���[�� ��n��ć(�ПTH}
�d&��"h�#�hav#ź9�M!%=�p=�AC�<��ܩ2'��50��5�2��>A�W;c�
�S���[k��1R��}�y�C�K�s��k�X#&G3����l]����!!� uV��O�G�0TG,]mw+.�8�E��t?�^�t�N�
8��eɹ����<.��u<`{�7�O��ݣne��Uâ�+^=�]�J�p�1t�V{�����i��*@"�8T`�
pI��H�d�(���z���V۩�dA��J\w�))�D�֯��s��0����ցm,�Ib}��A��ce�\���slpsptg�x���KȚB<�V����e��8A"B�G���H�-�H<=_V�6*@2��|�)S�R�kT=*�1_qkh;lx�{'���%��W�NOm�b�{ml�U ��oIp��C�q�wp���w�er2��v^��P��}gg�����x�٣!�ϸ�=���?��6D]N�"���}g��J͌׎K���U��LL�/S�O1e���q��L��� �/KE����.�9B��g�&Z�֪�d�^��bۦ����})����C���Uj^�Mym��=�Tx��B{�������K�	orSs��ڃX4!����f������WO�>�<$$S[�n0na�Y��2���Up-�}h"/Ձל���S�k�rn���+������Eovo-hra�!	���i+�T�2���f���	6⋀����=�X٢V���*9���9��Qpt�{5��=�̄�h%����BXJIh��������͋B���z\�l|sM�!�0,��9j��k���h�k>�x�?B���|�~H��ҝ8�G�N�A��1�r~�]ݏ�LNӶ�tI_� �ˇP�����m0N�'��.��oP�ldWUdRl��؏�� -�)��-���e�)Ϊv�wf�Gm���B�F�2)��m�(P|��]E���u�
�L��"��5E�Fp{�v�^�(��4�5_�w3�o�W��4QW��`ӻ3�%S����������>n�ߞA*'��$r�8z�F�+�S���S*
M���ꡖ��@PgT�n��H�5A��ϩ�s"�ԕ��/�Z϶���'b;��>9��n,
K\嘾�7���&&��{g� =����
t�<0%��/�?Kh�s(����ed#	��Mܖ.yS3��!sմ��(E���$W�|L^�߂@1s�<�?3��Z���ߓ�=)�3���YM@g�h�h޳��6����F�S�v��fR�����oی�/�@[�j"�w��E��z���xE�A���ʴ `F��3�Ki5�k�Y��<��3k�=b�ǁ�V ��W�5Oz�d�A��>T�� :uf��/�.�����[�v?�GC����VK'U�sڹQ��qK
��FlkV5d��3k4�1p�V5�yt
P�+=<({7c���^{�;=��/�0I���#i9@܈'�pݕ#R��v��=mN~��^�0E�/a��B+�t����~�5X��gFO�4?�Q��!�+�Yl90#�j��d���|{��T<��������U���F?ǵb(+H9�|\�$��Tg^5���sU�v�|���"�]���&�wQY6nHY�7^��H������~��3�5�z�<"���9<ڑ�C�� 9�^��˟=�Y �erUe�7x}c����R�r_L���ֿ���<R����RJ��s��u���s�W3�y�B�d�S��H z�J�lH���g�EO�@�B!t�L�	e�)8r��W�1T"��+!�YDTj$�w�Bǣ���M�٫6K=��JO����~�τ��՚ˮi$�$&�衬�Ӓ����Σ`��>9���Y]��.]�)�{�m*j�a
����[՘K��ף�����VppjP������DX|WC�i�hP�|T��FT��RL�3��4J[�k��6�	h�[�<Ȭj�g=z����]B	vD����fP���|I�G��,\���w~�&}��G���� ���.���`��{�g�]c2Lx��^�nD[R-�~U�jl�6�8:�$��XN��!���rE'ˀ>3Kr��*�r��=`���5+nX��2W%a!o��vr�=>0ES���B�&���葘Y��_u�bc{�.�Zjڣ](HMQf_V�NbMQ�VF�DZ�oaX�-�]d�\"����
�VÂ���sAp�
gṌo!��_,ZQ��{���m������QE�~1���N��.:�~.�0�-���v���[�6���kNLOC4�E���� ���t`�J�3�|�9�q�t��~g�Չ��c&d~uΖ��!�®�0�ܸ�1�C��:����_�={P�]�'O0���qQ��.�<�&'B�N��Q�v��3ӨÎ�ʹJ\��Y�{G�hI�_B�E����.�QZ�FմD�i?).�)��҄٥Y���jF�n?@>�q� ����2!$
K<Ǚ���Y���ب���}�7�3��Q}i�iz44�s+3O�F�8j��k��)�6��34�d|z`��N�.;Dz��č��{D�IDc�JM���9�Q������2�O�ޘ�h�p��R9~� ���1��/���(�#<��ݪ��A�7��5k([��$��2fK�6�ڊ�ۋw2G�p���>�kP�I� !����⤓G�� ��k�{ǉ���e���ޝ�S�
��⪸��.�w��|YK�Ry4��ܰ�jY��d'�b�6�H�"�83)�Ɔ��͸��oà{ _ȾD����כù�6�(R��S+�-������%nQZ1ͷ\�"OUI�����G��<���t��Bi`��8���t\�,y�Di!:~�qJ�@Bv[���b�b;\��6.
c��-}�ygw�!\��"�.3wkrzg�osw���'7�+��R]{�)��^z ˑ0��.�>,FA�`���,KN#��M,ߏr9g@thQ%�fسf!Uq��~8I��_j^[W�[(������WC��0w�H��R
d���T�
3����ٞ��,��	���T�]���䍢q����D���b��މ��3�A��D4~k}�o9=��F<�*2zY֛d�,-�!����^�����?��qM�Ց*��`���b�x��:��|kW����k��x�d�ȃcn{`����#�><�o���@4�pP�FId�Ca�7Ҽ,�k�v�!S��O*�Se
�o�c:��5oY.�7�c��3t�Y�|�DQw�'o,O���EY��,S��Y���\K�u���K1g�� pj�*���U�'%�3�	?�b·���5�3�/�L����Ѫ���L��me\�[�B�� ��ө�e�@�p%Ǔ�L��U�G[.1X����4��ةF6���{c��������Y��~\�NH��G�D0�7�e�
Q��-d��]g[ ��	�'?�e��;<Ki��~o�'(��UA�v������&" �HaQ�\z(�(�Dь��A����C6u?�uZ6��T3��yD��ǐ��eT{Ⰿ�غUa?��9Ċ?��]�t�&58����(���R|��-�+\�%����G�`h��|��^&��f�}��Y#���Mz�|ŋ{�(&��XUn0��Md����iK3�fP�A��g��8��r�,���g�_`r������I�ن��S���Uy(R���4��V#s�����'~ Z��A��|D�0F�t�����|91��I?T� k�vBX���C8�4	�}5��|�A��3&R���iDD�T8Ka21�!�BOg3^[�W�9*�C<��l��O'b�P.�L����w/��W�F��Y��J��S�~���\UQk|9*J�%�W�����h���z����Nܗ1a�3���1��*�|���g�i����`bU\������%FH~2�Z1>��8rƔZɊ�!/ݷkS�Ï/��<��YƔW�^h��q��|���攞�\�ڗY�xŅ ���t=F!��-a�a'$Ro�A0�<4�w]W��Q��M����G��O�I�Du��0���]�5�j��PU�$U�q>N2z^�N�)��g?�;��Jƨ\�����_Q�C�\#��U	ĭ	sq|�J��*Z ���ʠ�?��� �&�V���b&}���<gR�6X��D��7ݒ%��.�F�t>��!ǃ��HF���ǰI�� +��_�z�+_��d=a�w�2q���>{]@��h�=�����F�;`Vٜ-�HM��/����5_F�z*��+v��2�F������<�� _%��l��E�WA^�����=�oP�#�!����S�b����Ny��I+��P�(|���K�S.{(e^G)���:Pj6�By:ѓ�'�����8��(�rJ�qf��N7{��V%��|B%��e�X����l��J��s�����`�%��V�fS�)*HR�m^�d�"i���u̵ٟ
�E��qL�2�)���+�Fx��uΏ��6���
��V���w�K��bߩue�|�/�3�)��J�q�e�V��| :���	���V�&�� O�2+���W�����Y���+�Qd������|��4�+� S'���8r/��wu�a ǣƶhOG�� �|�T��"����1�Lj�/�5l<�m�J�Pf��@�h�nLu�<�2S/�=J�W��Sy�� %��i�8��Q'.�٭1Ʌ�����������]zy[Y/���`���L������-� ]����_W"?�h����X�9���r�W��`��N�j,��pw�P6�e��Z�@�0A]m�6���8S��ʘ>T���:	�deYrO�k=��#3x�OeT���a�ީV�wV�d��5�bJ�I�;�Ptx18V���v#��ºR�i����Ee��!M��Ms��`p���\%�!���`���.��~0�WqT���~�jC�g�]4B�KY_��^��mQ��C�\pX~3�ɘ
�/^2����@��ORؐH������I	F����T��%��}|K�vn#j�{#��U���:ꕴNA2eҶB���D!{@�B����SP�#�;�M�&ng�>:�X�]�g$k��Sf�&r�k�����Wv�C`ݘ�޴P��a�ٸ�O��!n��rӌ�焑���:B{u��2k��̡���W�׍�[�/�-�&�:�#gȬ%`lT��&��t�Tؕwtz+�IN��>��;�P�@v�>����N��}W@� k�
h���{�����BL�G	�P����݃6�ʟ���3��Qȯ%��m3�"�2u��v�4t*�ቼ����q;�D�evaN�:�����/��k��*���ĲśW��m��<�k��$!�W��!
��	r-I�L��~�T��t�����/����?��s46���7�g�z�����TN����!�_��iױ����㋠��b/��0w� ��Y>�w�As���MP�d��`)ɴ+S�f<O��_���gm���\'�EȧԴ�Ǯ����?�ݺF_�g���2�(p"o��U3��0Z���m	IةQrKx�ߒ6�Y�@�"|%���6���o��M#���7Yg�5`@pɻ�`�6��/�C����#R�����,�����a]��%W�Q;o��:@٣a������|76iF��w38�l���� VCr��ӳ �N�T@��4�dwA�	�<I�[%qx�$8Cf�������,kG�_%��g�|\$N� ��>j>t'B~'a�d��2{]i���z�C7L���?�JQ׊��u"d4%g=�a�ּՉ%�;������X�@q�L3�Š�4�'тhK��o�*?$�&���q�X��`�2ɯM���9H+��&]�O�r�ԭL�{�a��cS���ڱR[.��e��_E,���.�1�q�	2.����Ά��G�Ýh5������f��`����^UNrZ5��ї��ROG������К�4֎�ViS����	��f�zj�Af����`];��S{�u�N�����\ҡ��w���1�29�'Ȱ�FL<��/R}!�I@�.zy��� �.*��X�Ye=������@��T�x"*�7�U�5E��		,sdKߍ��1PvvjZ��mS���t^U��C�n)7+¾�U�ac�+���2Q�G����l3�:������a�uPoX��!�F�N�$ͱ��%��a�����[�Q�*rH;�NCHRk��M3����䏏��2:������w2~��5\·�����V�dV���C��� ���*���.T��u��Xe����d�(4�Z\_�-߭��un�S�Z�S�p��Yz�o r��ls6�~L���Gy���I���/���0��H���(Xw�b�o���i k��sސ��`���c<B���F5qwo&=n���`��P�j7��J�bIi������N�G�%DQ����	�.��� �*� ���s�8mRUUE���1,�Ž'���W/�{^;��e��D\/cQ�
i��d���+:��*S�2��b*�q��F
,�4r3M- ���Y**�p�����\G�%���VG��k��I�ġ�P��=V0H��5D�7w����m��"���5tZ��Cig�������	�NFAZq�ty���Xg«��X�'�k�{:I��1ʃ�ɓ�4�����t�B��m�y��%���/�4F�p
����C�mf�����j7�d]�C��f�k
�U��>�
O�b��i�����?;�$���`��Ƃ�Փy��85~�(���y|��e�DQA%i	۠�c2"����s�&�}������B�{�+�������{,A��\8i���J��X���7��lTP�M1��������?� 0��k���5����>��Kw��Q:O�dH�M�AB��*Z}l��=T�������_\�\��;.�!�V���������Q%AT'�/�S&o���7�]s�X�
ᓿ���?��ǹ8Կ<'��[�	��aK�?�a�iE��*3�΃"&���&����۸n��Cz���Cw�G�n��
����3`�U"�8�G'��ڔlN�����d?ko�"��sZ�ͻ���(ץ�i�fIV/"�@`�8�s�Y-pܩ0�⇐��N]�C���4�G?=Q\�B�6��_���@��-r�{f�m0Ӓ��9YmU�`e�Dw��'�b�ꄬ�f�<�WQP����1��5[�A���K�']��.��l��d�0Iu^q����Y��v�|��ҢV��h���ɦݳ.��Z�	��W]RX{��E� v�K&v��˯{��?j�?��=��&ZY%��Ϋ��2� � ��٪��3n�m%ܩ�w'�6�[v�"BLb����VNs�mDPq��p6����¶�)^�l�o�m�[��v��FG��+�'V_.�e R7j�Kb·R5J���楇T�{ǐ��b���"n������?��*�� 蔗�H�J��MZNh6�0'2mU�_��`���V�A�)j��Yݝ�&� �l��g�z�w�-������w�'���[�9�ט���+�k��W��W���Ĝ��ֵ���40!S��V�|�H{�Qr�R��c���gq������H�9=�2~���7}��Mm����j�:�_
$�XH.v7�A����r��eP�CV��t�/a�τ�2j_
�y��0��d�Z5i�}4��M����u����]��9k�z�����%+׶��C�<�J�,^@: �]�����2��Fn�ȫ@F�Gs�|�z�A+Y�B���E�ӵ#.�mP������xS�^�]|7ңA	��XX�=d2P�,�L8Ԏ���T���і+��E3���ϩ�,��c���k>4�\̎t�A���5/~���V�k�q�=d���k%�@�u�z�^UFѼO&�C	�~iS��ZV�?o�o��~�$-�%�[���J�n�!������0��%��⚅�ŀ����g��U����#ȸ�<4��?�vI��
4sW����)s|ʦ����#kgh��%�0;E��hV�#OBz��#�nZQ�r�k�k�d+�TRX֎�ښ�ŊEJ�H�g��Ϟ �9G��us2��/�%F���k�u�?�;��-te�_v����M3���n�N�d4�
�k���w���R���\�3.��Q��e�9
��)%앖!eēzڵ��ҹiMfh�vx@�/��!d ��m�7�����y�6��9�����*Fv��:?#o���Dx�����:�cדֿO��{��?ؔ�1�g����tV���z�,�\y�[�(�aD`7*Xϩ}�u��L���y��+��#��Q�-8��&�v����=d���H�3cM<!U�oR�C��*�.�(I�03�Ƥ�n�Ћ'�{�nU)�_�Ei�e�3�$�R+�듑��2�{!�%�������d�:4����U2L�SD��o��z�Bz�_��a���o%`�P�E��Zr��z�qpa�ol�����̡;������O���{kkޑI�w{�UZ����5al��yC����X�����c�+rp�Լ*�},&|�V��*�y�\��i�j���L�(����,�6� �<O�fRTT�-$������8Ш���su�Kfz��_���km	���WH�],Ң���R@�N�xl׆6J�7e��M���OV���*�I�S�0�)2�|�ܻ�bNV�J2�����7,�mB�I3��[g%[���Ѣ� E�:m/����e�V�dR��9W�U���(��m��qW�%u.R�/Pn����|��	sv���̚�d�y�'o>ԓv+,CI���DM�����m�Km�����;,f�^�}D{$.� ��ۊ\���*��1��;^FG�rA_* �&���G��+I*�~����؍<|���n~�k����o��+�H|}�n�2s�Par=E;��r)�C��<�_��L|)��MLg����^�a�6��(py��4�e��Sh��)�l䟰[�@-�/����eu�8o�������rTR�C��D'=���B��Sg��r�v��������Fkè!�8��y'��4�3�u���C�~�i@�1��~{�&?�~�	�lǃ1 9"Zʕc�>�(Q���f��ʻl�B杏��S����5��*�> /.��ȁ���V�u��]���X<��-Sa+M��(���l����Md^4�G��3x{�T;�K#"� �J	�}>m���h��9vPJ�b׸Zqn��
�7��\������po5y��z�8���Ll}S�F|����~{��Z�-v�T Q�ގ�RNAˊe�F�6��,t�p}6����i���)����X���p�n>Ũ��(��v �����y�c^�@Ω��',f�ʇ�4]Ŷ��T�-kK����[�o���	`<yw�V)��N��'- ��������BKX6�@k�&�C�2�eo)/_/U~Qq��õ�@<��ӓ�
��J�*>��<|~��H�t��ٜ�޵`�@�*�XPсS�'��QSG�n�ԧ����@P쨗��|`��mg% Ae;�܂Ӻ���G(��
�sK�_lΦpv"�����#۫n������ʯ�,��T���X�#!�$F����VE��GI����(�4Vԭc{F� �ޅ|@�5R���5�l���ه��{w�{�9rb�w?��9�/W���3�mZҏQ2C�9z*����9}�����v���+.��#s�3ޖ��4�`8t��#."����(��&>�d���(�6
��C�J��^��T ĉs@yp��w��w���߻�3a�Mmc	+r���#�~"	l�V�<�&.�k$��Q�9z>7PH�&�u0���خ	�\.د�P���,����v���
y$�꥘��/�/���9�o,90�����#�6%�$e�����Lή�3��t�Iez"����T��<\ b��D�@�:�
̀P���݁�w�O�5qU�}�4��%�$���{lRx0Y��UA���	��%$@z��N�{ͩk�P��F e���������N��$�6����?&�g���4���m����h��ؗ�=
:X>xk3�[�n���(;rp�[{5_�I����i877�e̥��2G=	����oQ��,�w	ю*��N8^��u�w�|ܼ�9��c(�}S&�C����f�T.��\��0
�����*�=����L���4�x	�:�Ȫ
�Z��%&���.��-�W�F�2��7\�ZW����U�ϖ�1ֽ(tv��|�+4t7iqG��L�Q-��������'a��� �Zp���S���V~$�\��ĈC�j'���<�E�_�¥� U�(Nq�0:HHt��5�x"�5.լ0�죾�=���]��Q�������q�+���A���bA޺�!7mmT����
�vp��C֌�i�m�Y�&�*I�����1Z�WGvWHӰK�_��l��cSN�g����F�p-�馚��%r���^���;��3[����HP���U��Zu<F/7;+S�H9�'�����Q>^:�L&~l��if����E�\\e��"�2���i^3+����v���� �ʀv����c������+B����ܻK� ��Z�k{F����i���}��g��y	\}	K�����@�������s�U����	v7��j�l�+���O��&D�����at�R�/��v�U$sMC�7��
`��� *��ç�F�����AE�r�52Y�`*�����m+�G�.�x�U��z�ă���d% ��T�y��d��F]�ox�2��C�XY�7��%�g�
��e�|��;��G����J��u��)6�M6W�A����_ىp�B��A�O����aw z*1�c~e<���Xß?V5ұ��B��Q	�E=��eCMr6�`o�$�w)+߬ J}ᥞ繀�'�s�paQP.���a+�����20�T4�Yӈ�����Rp�IY�n��w��l���.LIW#Twױ�H��R�|�lL�ڈ
!e�U�9���K��	w5�_�q��\jPd�a������2��F�Ţ������������I����OoT���DB)�=�{L�� i"눦
��٘�	z\V'�h�'�HP�c�u�����e�w��
�3*�6�+�H������?
&m;�(
�_�/a]I��[��8���>ѱWB�4�W�T&�Bf�$5/D�B���� <�Y�C�k^@�i2��Qs������8���1�<�R�96���En����u��%�p��6љ�G1v4�x�oWIl���}~e��{^(��!٠����ԛ�����Y}�m��f�x&$�����Z�-�����S��<�rN��8!|�,�o�#ƕ�Xv;B獍�#�-C���_�Z!��R�|��KP$_g���
--��*m�����0`�W?I�%	�H�����ѹ�,=�2������đ�U5��r>�m�D~Gy�n��FqΥP4Ȁ�u�g�ɽ�d?�����?����q����O��1Jw�� �րB��]�$�<NX��[���$�79�F�T��s_CTn@bU7�B�ʓ��`>�d�}lGg���r@��]��� ��*��v�vv���p�M; �#�[��l4^t�w���~jd4�'��#�o��E�� ��"+3�^�n6�z���}���|'�r���E)�)�������̈́S�'Ja���Lݥ��C�Rp�6;3v���+��4��Zjm#���k-��e-<"��=tK.FO:�A�ܣ�S3Y��bK)�u���m�A�� �[�:o����zo�%>���z`�8A*_f`����}^�3S]��h�^k�~�57F���7_bњ
��u��6�$�� ����_q)������خ �@��eO�}s�.EϦf��.M�tOE�[��U3�K�-���^x���i�!�z�&�wN�$l(R\t���6/
��;��훿�m�u��Qг)p�� �i%/� �H~�-�Rok(�׈-08K��#�!R�0�m�&+�C�<z Yi�IL�#_{cIx(�2�z �lj�[X�:��l3��W����u�����_{$���	w�X�G�?^i�_���3Qk͙~˒BSB��~�Z�de�̙�$�� P�E�Y��,�N��I^���q
^�"!�X�1d$~������M����,��~6�k^5f]4�堥w���*������.syT���eK�7ߔP�Ep�q8���#�Ք��S=�:/��e�M.�gɐ�?�ɲ�"&����*)X��C��6����z����K����o�V۱f�+��_��=Sʬk*�A�5��8N8���w+dO��� ��J���ma	�q"��`�C��A���fI��X㘋����Ⱥ߱�6���c�
�V>�4ɣ=��'s�˫fv=���0�/QC���)7��
1�d�~�	�iDw-���Ćg Ʒ/5�2{e���u�qS|G@ �1rA~jJ�+���U�����9�wC�w}��,�����)}���jE|{�Ͷ--�
?eUD���i�t��ײ*��.�i�'G~$ z�9�YP���Ei��t���V�|8d��ܻ��N^
�����~i��~�h>i��>G�S]�N�Z���`D?��:lኳ�pQ�g�Qy5����L��)�/����jxX*8eǁ�'����n���c��܃�xc�� b}���Z���_b���Z�����\d'�6F�h�aOt۵A�ZS���|' e���E��QU�3�E��/Q�������ŭM_˥�b"v���#cw
���f6����B���G_թE�ף&��q5JȜϤ�?KcjH(�JB��q��}na��1jN�y��4d���r��w�����v�W�eyW��b
��(u�[BZ���/�tݫ^���IL���'���1 d�y�������l+`�2�YMp��5?$L#0�m��d������l���w�0�v�D�R:�Z��R̭ՠ��W� o�J��	LO`�Vע�B��p5��P\�ѐQ�S>�v�%��P!�(�p�U3�R_����6}r::�>�+�'K��֜ '$���IWD,�Tɓ���>�	4�'PIcU�w�0�Mc�E����[���S+��;���jARW ݁ ����ˣ��΅+f�BD{������n4�ƹ�ݻc�����=�j���v0~�A�t�٬��/�iJ��9~�f�ˈ�h��0y0ZAHN�f�;#R��lo`A��Y�BV�f<j���T��]���Rߔ�B�����E�J����zW!��.��rD��ҵ׭m�e^�Vٜ�c//�G��%��+"�>���[qM6֟��hʋb��誾�)��bh�)0��i��ft�[���ͮ����
#ڪ��w�`�#���2��o�3�?���^;���h����4�axN�_�(*r�U�K������PǓ?�BS�.Y�өE��������$��iY�{ڼ�`uִ|���Ϧ��V
f//]F�]Ln;�Ղ<�6�J�Ԓ��I�N� ���4xb�dJ��FC(�AȲ@t��Q��'h��1Gv7�\�2���Ǭ29� r��w\JߵP�[�a�&��1^��-�ޏ�����}����>�;f������q7�J�<�kcإ�T����T���My�]T�``�z�n�QRߺ�/dZ��c�}F�(��r�7Lp��M;��Û��#����"ë��F��%�E��3;�q�-z�^���F*�����~�s��L;��8�<�~՚V�S��D$D�w�GPj�ɼ��Ds+]��mQ֓�0dw��As�hBjt��dt�g�[h�7l����؅�U�^�����
%��ަE�%ہn�-�"��,Hqo3��2��EX0�N�������s�ko��?�P)�L����G�Ȼ���0�+:��e|�x6������M{��nGv����F��7n��G���[9姺��C2��%�%nE���w�5$���BPv2r
b������V�&={�!��s�h��� 3I^O���R����b=��qfhި�3�%f1k�x�w�~g�a�z�E��֤e���4��w:g�v���Su7-�"E�W�~��0�\�|��\<�1��R��ry��^�z e���A����mb�s�j",_m%���"�h
�B':~T� ��EUґ֊M��C o2�v+�*஧w���{C�296 ��/�ӥb��^�"9�^�s?��r$��aE�b'�^�6/@�A�hx�%��\�M�_;�li2�g���n� ��愜����.R^������֬~��q��o���&��:a�e���	Ԩ���d�j\t�=���=�$���z.���N�Ϻ>�)n�Ǧ�lYޥn� <	��l�\�Qlز��T�F�+o�]�{�u2I=(=��ʙ;yD�r��AV��O�
�'g�u�ߚ��3��*eJ���|O��B�v��&bQ��ᅫ�����/��$'�������}V �.�Zcb@����jH���zs�ʣX������+�sa��Zg�;��b��l�^#M>�{�
fbd���b��_�K�`eXMr	�E�Ȁ��C�R��+��5w���ɉ��ؠ]�Զ��<�X�aIl���tx�a����r=?P�[=��R#��M\�;���tW9Q/�_w(,܈��AHSZ������V^½g�޶����M	�RٖkK�>�N�/Q]l$T�k4�Ǩˮ�i󫒷G.'FM��,�0�8�MT�b���F�r5ȡ�~?��u�w��K|\��ևc��4ѸN�F��v.+o���`��nsq����nb��� h�]�6D���6��洟=��a��)���5��"�U��|�R<!x��~����cw��z�%�f�U�"_K������t�$�۟ye�E�&C����MZ3���4J>�ʰ�zm��	Ekp�pe���;��h�i.4��x�Ϩ~����y�[���1���p�2j�k\�d<����T +U�=kGBFf�s���3�З(�ȋ�/�T�U�Q��=����N�Q)8r�@9���7)�T�3�mu�=Ϩ(�-�x�x�A�nJ�`S�d7����]�4 e�R>�\�{x_*m�D�������g����I0�d���S�t��$2��p�ٰ'�M�!����]H4��+�,�-<{��`�i�SQ�Gqγ� ����lB������Rm�p����f�+�A��������$�P�����G7�ͤ}O�r�	5+�_/�c�TD�:�SղL�Q��}�N��.��<cst��u(�����g`$6�k�]z�A�v��]\|1������3�GZ�= �Q �/l��A��D��"��e.�W�s�3��24���,I�C_��֭�f����B����:+Z�S`���OɅ�����0�}}���#��	��gwZ�J&G����I6
i��BN��O�I��S�Hf.���߃3ւ����
�N�c2"0�w�ܥ�Q���|2�vxn1�a�/�4�Y� M�e�@���CZV�U�� ���8V�JQ*�o���=�f��8C��-]�퇹[�%���S�VaqD�5�^��Gl�IP�� ��@�L����>{�jz��r~�T��
��!������ן�{\`��2�����mM8�d
b�X�2/�f�� ��6�����]3#��'/��BE/��nV`\'a�����҇��,L���)�y_�Qe_�v����+�M�T\m�okıt�
ةY�e<p:�;��z84tC$��25o@�O��Gޅ:�-:����i1%�0I/v��,ꑻɟa�T�rʖ������5)2**:�����+*9�d[oc���j�N-�7�3,Гr�uE�͞ي��O�ä�ԑ�I)ܢ��z�!�N��c�ѹ���{g�����$6ms����.��v�[�N��\��B-/�jPe��>&�xZ)�؋�H`�|.����*<痚�����r��^��'���&/栫����BH�A�"�_��_<}C���q˩}:ʆ+wڼ��+q�}>1��5Ȋ�,��$�̷cs��'ӳ�����cs�JE��h9$_�0��qk�@}�N�!	]���>���<c��Zk�oǍ1��U[DRt�����'�B��2��ĝ�bQc�y5̃�S�X8n���
f"wEZ�E!�C���s5�sɿ~3��%�(q*%���A@ U�y�W@������e��Ę�^�`}ͱboH�*��	�U�d�W�o �R�*��N|�G�nh���58��3g��Q�,T*���B3f�s:����:������w�7��tax8��F�V��nͤ�6F~�%s������{��>Tg��]_�4�V����_%����T�_#�������2m�wѵc~L��N*e�Ǩc~�S6�1ޭރt qK�&�� z �uugM�#K|Q��L}^�����Ac����#�i�s�������P�7��Ԓ�Xw�q��C�\6�El\���/l\p��{�,�2	���9yW��iS�F���J�C��2y�W�0�pp�z��99���Ȕ�T�[ȡ)�mݢ�{u�z����ߧD���|�c��Ubڧ��F�\�"�׆����(NS~?\ށ���M�:�٧�1E��x�^�S?�$�X�B�ߙ�3)_��GXB���jnV#G}y�{oQ���PI0O���"P�����Ԥ_R>���~f��c4~���[j������+x��j%�~[M���v=ދ�T�R�8|��e�T�ߜe���ip�Q:�3����$��Tls/��˧dK�X�T����>�O�!�;�q���wk�YC�П�<�*��HjGOZ+�� (�:H\�v��cpd�┺Z�/���<ɉ��"Ä�+Mw�Z!퐟x�Y�#g��p:+�2���<�,e����I�J*�ZgG���J�G�Wv��l��kD�[��3|��˾�*�!�/�G�9AMbjZeQ��y0O,�K����;!47�>~�Lf�:o����R�EN,ߢW���=/�!��gŌ)��m-n���Nf��(B0 n��p\͉k���*��O# F4d4��|yv������/#��(��;��kB�.�C�Z�('�6�`FL������ԛ�4�eS��Uz;!��f'�W�?p:���/���a��(�Y_y[��h��}H����V�,��^�Cѥ�T�[����7
�BmzȬ쁯[�1�V���;Bw��d2�����ݻT�M���^�ˢyo�]8��6��������~f٢���;�	A������!�G�L�.d���Z^qM��߅�-�e�·��Zk�ql����Κs�XJi�YX��jE��\!�j�S�^���E���������-� ���T�T����aB�.t3��ӓtg�*���g �zt'�wu,l���4`���(Kɯ@hfa��@a=�Md+���}�뀵c�����1���Pe�B}<Ҕ�rD;��U����̛�
��j��dr�:@�3�|AMc�əl�ypNni�TZ)ӱ�?�V�ir�i��vSU�����
���	7��8ȕ�Њ���EJ�G��@Y�@8����'��k�D8Vǔ�<$���l�={18�h��t����!�Ȋ��3�裏�X
S>6��Bq�PՋ�~G����r~	����o�wlKL�����:��� cb�s
�^�X��P�E�ǠO�Gߕ�)$a]h5�0� �~��Խ��(�u T�,�$^�D�V�����8�-�C��'`#���T���S��`2��7-e,�n�&�7����M�>�DTa:EUo
j�e��lZ���Vu����f���%�(-�������!=�����ks��Ҕ��x;���M�%���W��<�?_J���;A{����U��Xs�~�p�����(*[���E�Qo�'�ki.�R�%I�wr�Su{��/aS���i�@*���瑤 �ާ;�S9yq��$�1���
�TJ���!��RAjW}p�&p�K��H�S��=��-?���`?}�����\��|��ﻬ�v-�:@���޹U~�un�:���O�'�Us���S"���9�o�����2Hhg�*���a�]��|zhB� a55�.�N�Q�!�������R��������i��C&�h$�E�~���O�C]ui	}�9V�(�;:�
dR�tpc���g�"�y�]�]�_K��?hÄ���݆���"��&p�D
j6�p�"���W��)��W�"���#��R���y$DF�2��z���?�"b�4$Ji_4�N	�7���Є��Y�#r�=PW�ihQ*��7ͅCVU�dC�,)m=�/o����S�wBw���_�.R�\��~��^u��2m��U���\����!����rs9�*�Fp�u8\��G�G>�E�,����*VV
Yfz�vO�(���0B��W�鷒 \V�G"���=��×H1�1�h��|�p $���y�Y-�V�]����_M|
��e���H���u�Ca�Ꞹ=Ix9��\q���݂���Ng�sk4�ؔ� ��>}����w���J��-���$_���g�}b����Ȥ�k��ȕ����+B�XL�KU#������O��ו�G1·������7q����v).���5��0k�`��Ӧ������ϩ/01͓�# ��t�k�����NZ�w-��G��讱E8Q��z��m�~�e^�}u�Od@��+;��`���|G�y7�5�[^]��3{�s�����*�� g����1^�`&=�D��S�H�ϩTV2"�C������@�4^ie��7�_�R�s���Ob�w���ʂ��\>t��%���Ŧ��U�7��YJ�PcC?Ϙ�c�	�4 '�]5]B�`�6؇�o/l�D�9gN�?
� H���v,�嚫����#�y*·*����F�=l%�O� ��@���O�Z�^�w'�<�N%%�M�M�q�\�Q��7V�OX$������ ��cw�og
�d�H\��	��*�����T�C4eOܙ�*�^��Dޥ�X�Q��V�6G� T���)!�򼡱��W#b����Q��D���em���e{��x$�>y�B�}�c�Go�~�Q:%[�_�{��R�\�_�p�T<��'�����j����9�.��z�n�Z���i��R�z��N��_��mD:��m�v} "����&�O�R�w��CCX���:���]>�fW�h��P���z�.���uV��o	ѫ}�Ս�ݢQ�7mV���X��µ�Qt�y���g�k�dz?2ow���X��%[�bgT��Q�nT��6�/�T���,��д��<P�ٰK"�8��}��!!�O�Y�v��@ ��_��T����FB}���¦��P���m�"��@�Q2�]B��
�\�΃O9�՞���%�����$K�9J����>� �-����9j��U2�h�e�kn����Jt㔁�?�W"k���s�X��hw�p�o�u��l��?��OY|�~Kl�t��p�{\a�}@���G���S���S�����U!{�C7���2���r	Մ���� ���s��^���@��|B(�����|>�z�@��H� ��[,��7o	,[E�\��U7я���uB����b�y�#��+��]���UL�vE�'�Pj�v5/҇���x^�Ȟ �I�~U:�(���xϊ*�t�-ԭ6���:Ԥ:/+���$�5���T�C�`�4?m�}ڽ��_���|�1�˳Ok��+8q*{����;&��\�UZw0�k��;�N-�l���1��ۊ,Mm�tF�eԝ�qHw�ݍF�;� 7~w^ovʓΛu��Y������T�ɣ��P`� �q4�a����\�;��5��.���({����'��0�L`���һ����!�6K:�?��<g��5ve$ɸhN�t\Lm���^�>��7_x�������N���WDs�CuV����T�@����6 Jòz}ҴD���졳,�_+Jk�����>q�N��Gb��	W�pf4�Ag9�2Z�,z$��4�3���Ī,j��x�+aH��g�k-Wy�f쀸J�=��G���הt�͢S\��s٭�b�vt� s-_YE�f�����!�}��4�W�E8X�L�
��N@�˜[��N�_+��^�PDk�hR��_�S;�� ��O�J�^Y�%[���K?��o�kat���0���KK�j� ���R�^{�co��ErY��@�<�(�U� 9	�;�?0�
����F�}�V ��y�kB�C�ɋ�i�F�[�������B�B�C�|�b�;4���~w+�n�ܓ��%J&�.߂H����	�%s1N�I����e��%�'
g�N2u��m�֊[��`[�� eH'���w3h�*�dZ�:���P�W�
(���g����a�k�31��/�Lb�����!7jȌ7YM�Vq�PIl�k`��V�u�;�ms�%��<�o?��̉�=q�A��3�_�p)Ě�n��^r���^�v�[���2H(Υ����� �&���"4��v px�ko�i�ϸ}�����8�w��t�M���"DuDY�S7鋕��o��ICj�	w����Y�?��8�Ԣ�Ft�)�\M?͏i��
�̈́~0�Q�����G��aE_���oL&�A��\�����H�.���!x5�~H
@z�ѪO��9�\JTr��}�.J�/%�0���g�n_O\/ ����:܈�3gG�&Lw���t��C���܄�K������dw%�(���?��%(�I�9�ɏ2t�Z�g�v�C��#�P��{�`Ű.��u����I����)u���.b�k�]��pw/cj5�F�)�c릋�a�-��&)Q��Oێ��]���U��G)?"���˲�8cD*���|�J[�X/�K�	݀�oc�(�"fD�>d؋��Q�p��bȢ5��T��h�fHK�`\�4f�J
T�X�Eֿ�*����G|[�����<c:��ڻ4ڹ']^#wh� �%Ӿ]g��==���И�}�W�����$ɪ��Ft2溂�82��EyԌ��"B,���R�3D\Pl�����y�g�z&GzHI���.�ְ{�Mv��6�>V&�b��d=��V���u]��$��i2��P��e��9�~��@����q����Fuft��9����<�;�tXۭ1J�c�(��@�H�b(}�y<�68H�cp�O��h#�v!6���$G
���(˱�-W�^}�ǘ2��a����JhJ��#��I�^�lq���64���H���a+ ������ïo۲�p����&�Gvg�w3�VR�P �3�H�\ W�߁l����]�g���O<���7!�5��K�e�?N���+�l���辰gM�i���OÇ�:�������՟4��1�p��HWp� j1����pٜ��CI���h�;S'N�����N���kbs]�6�oE�_�?�S�g��&x�8�w|0$)C���|���,����wM^"UB
�@��;���Y�p-�$*�ȡ��Z����e<�=pwO���`_�������?Т��u����5[.����w�4�S�����x��,=r*X��[�{V7J�І鐬RyR���7U��^��^	I5y�;�2��L�����05R�x�^.��'F����W��k���/��#E�)H�6��s��q[�M<}3�(�
X4�� �!����Sf��8��d�6R���������5�ͻ���}���:��oB��v�l�ګlt$����� u�+*͟X�d�t��66���(�[JQTl��mn,����}&��e�ѻ.���`1t	DO��{.sr=�;�;�Kx��qt��7�9`^���% 7eR���I>gY��M-n���\ih��F�o�_Zc)Q
&��!�	
�_sf*�Z�f�GD-�uɁ��,QE��'�.�J|w�k=���,����J����Q8j���|�����ն,����h;�hݨoD|�>��ݐ��p����B=��#�9X���ǒ�
\y塪�pT�%?���#o��>�/n�����v00S�h�7
�T�ip��z�§�Mq���@�5h��s�b�|}r�,��hE�\�K�B��a�m7M�礬Q�g܋�A&���bQ�����}!'�A�N���-�~]����%�9�.	�uH����=�wZ6-�g8-��Bo2�h=}���Mx5��}I�΃XH__9��\p/�Tt���G�^��Vc"K��,
*1���4X��h����]�;81���H�Q��},��t��ڼ��HG��5��`�L�I�ҌO�����Za�)��'���^�V�!�*��+�N�F�E��0Z��G�O)H<,��SeK5
8S	ud:u�
[�i�{h�Z.d�wHo��u��!��|�gc3�IN�p�&�_°Z���9��A#T�):pi:��@J����������Hʘ�Y�	�q�P���a�UMR���d�v2��!x�*�q�9?d�
'N��V�� /�gҞ��D���8|-���Fg�h*��c�sp�N��q�aT��@Ѝ�����5���~��#ʷ��d��E@�-e��G�+��� �LP]ǰ<q�L��Y#N�/����5�@"�]Fkw=�X��qC��X0la�4|��Ĵ�O�	�2^����W���!i�����>�l�*�8 �]���so0c7xY#3�+e��YF���1�~�[S%�P���B�����}�_�?ʇ��~ֱ��!w`���`�j�S�!����@�ا8*�y�|[*���N�WsĔV�5�d`�$��|��Ϻ�yjd1���#*����O�����4�� ��x��2^2����fp�J�}~_đ\�%����_����<�i#ː�z���}1�`NM܇�t�>�X���̛���3��98Ŀռ�"��Tw�Y��S/��x}�`5���3<
��z�w��{����7��{,�Ϧ�u��2��TKC6��fs%���	�)�pN�$>C����Y��:Y+�<��������v���0���E��yD�4�b��������r���Ε�*�Ώ�`�}���Z�N9�b4|�{=�2�������.ȱ/:ܥ�`���M��I��c��}[I'~V��~bY�} r���W\*D7�����t�Bö���� �9��gh���;���?�7�6&� Z�8�/�>����9��i8727'v4���Oh�O�����g�x���=�X���$s��:���q=�u}�5}��N��k��Q�T�1��$rp���*x����
P=0C�a8�i�	l?��og���)ʲ���MbTc��x�ȶ�����>��֮׿-+,!�*��IݵCxo?;��6y�u����1O�+�3O�
���C2�We�m$����a	���-$�������g���KӐ&4��.�iD�����0'@��P�:��1ȑK+���td|��� ~��՞^	���	j�w�M�vx
����F�R��>�w�Y�,NVG�8H��^��s`�Ý�%`M��*����+����c��V`쌄jb�gZR�_��+���a=��\��] ��c��^)UE	~Pu�v�D�g���A>����b�G�B��3sӶ�2�(�n�
�ݾψ�~��B�p�id%�ު
����	��+�|���9�F�5Q�����=+>�/{�i�������a��,g�IZ��B�P��Rm⩃�&���ӔD`�cO�>M��S���_��C"�����C�I��FN�UŌp¡rxR�L�m�6J'�t�P@��L�Ɥ*���w�Mo�^��xl��| �XSPj=2�׉V�`�R)��D�8�b�<P�|��'z������{]/������\����`h4,r�eo���r2����*��A��V>�<N$�O�H�[����c;}}�� ��/�j���"�B��I���������Z��F.��fCa���Om�*N/j�\��@�1���fP�#�j��� �#?�ݦ�v���c�U��Iy=жB�	�U}�Q�-�t��ޔ3���6u��74�4��o!:���1��,�ԙT�9��HN.N2K`R��H�3'��|}��8=�\f0��0R�=!Z�c��KL6xݍZ�k��I��6J.n-���=]��>�,����9u�ŐPy��[�ʀZ��ɅO -��Ҏjw�<5�{��Yp"�f�,v7q���9:ԁ16�<OUI�}lɸO�j���*ZB�gÊ��GuC'U��M�h��9l����PR��Z�P��k�J���4U��f�Ա2܍ﬤ�%][�Q�Q\��а�N�q/mj��x�Ӆ1��EfZ��A��!�}��U'��?wԭ�2�W��4�Uyݯ�{�ٗ/w6���*Flw���{�M�Ͻu��y���`�|A7�c�rW0M�Lі�f�|<-1�)(v��ݚ���Dr��W3�!�������v�il):V=�����C��Ψ�A�1�����8K��,w^�j\�9���)�Q�����%��ǖ(�`�R߰��݀ՌO5a�Ǡ~��������=�e.l��Y�ڸ�#�yM���I��V�ǂ�.J�v������޻��Hw%y��3L$�:k�%./:[���!�ir�9O�d+	�۸L���ExN������m(��C���?��j4�Y9~�(5������cC��|s�����Ê	x�66<�O��hZ����U	z�Cl�Ր� �1�G��/%�Z�a5M�u�Z��)�ߢ�����V0���t������c��;����-a�쾞0L�HVPZ��l��[@��t~�QF%�A�	z;N�� �LL���v�}\�D8��@  5����@MHh`�.�Yn8tM�#X.�OW}�ɲ�8�IYKNԣg��!$��K�h�(��+> @�b�l���ن#�0�+��>H�&N�(�8,�t���K@���6e��D�7��#Z,�$��M;Kv��و��EHY��*��(!�� X�.��qءG8�;�^���)!��&�����,j�[��񂗽߳�D�D�M�JU�������w-l����`df_�O���C����Qq��&b?�|}^�}��]D�<s�6�'ˊ%��@[^pͼ���r�~x�H���pRp��������|�%�B�3U�J�z� ���/$��Z�=���D�IIz��)r%F[g6wYl�i�%l�\T�i��s�L�ҧ�$���J�~�ì��JjS*����0õ�4�D$PxT���D#i�e���װ}��ڜW��ˢ��!cbF`��67'[��D��ؗv�ǟ��c�A��s�G�Hw���2��[������ύ.��M5�/|�i�8��cU��bzlu&��.f+�Q�ڽUz���c��c�YS�f�3�G�'�$�v��vs��M�����;<F��WP�Qnݍ���A"t�C��;��[���b��b:�5�.T�`&#�'4B�ש�\i9��+w� �L�����=�TXX��*�gF���	�a��]���~������ͦ�i�r4�ÿγ�ȇ_���H~������՜b�S��f�j�`.��j���O��,Y=a��~b薩eї	�}�A�C���?������n7�yzI����C^�r�H��0�V0��S9�� &)M�!�<.�Cr?/�b(���'���V'X��Qb�������]�c�U	�/���7~���)�&ԞO-Y��"~��z�Y�R�W��n٨��_Y��s�m��dW�^���,Pjo_���@�љ��^w7�!����. �����Iy� ��C9��/��r,7}��i쟪�
�oy���O�����D�$��\"o���b!�T�׈��wG^Ƿ3?|c�5��C�|O]�?���ԗWA'�{d�Y�[�ִ�`D�ړ�����	�D�ak�_��׍�}!?��N�!<��������z<CL�<Sy�/���H\ ����%� ;Jaa�=6�m������[#o�_~̢%X�1t�dY^�Ũ�!�9.����O�R|#����hG��cN��pe쐎���ݝ����z1�8Z�Bh@�<��ɿ֑E>��Q6��й	6C��>/~�F%�	��
PD6=8�Sy�PPQq���	6`��x�UMfr�/�,�w09I�� ����Έ~3p�\���m&���G`>��>E"���f
;�'��.���O++�%Z��(�:��3Oz����v��r��ٌ���G _J����Q��:�|�*({xz@ǘJ.�"h
��)��F�1=����P���T	�D����Z��^H)# }��xވ5��!6���x����Q9���B֡g�4�F΄;	xM��e��&&��t1!���B�W˾n����p]f��a�qU/�����	�cT~
jW�EU`��'j 	օp�oOu������������p����1H�_�[a߿��M�U�|J%Q�����~d��o����i�l�ۆ:�0��%cV1d�`k>K����-�I� R�s���VQ���m7�d����;=�^�	� %�����|Ƈ�,�LO��f�ћ�D/�R���������2�`]X

wsV���ʚ�����} [�Sצ���~��1R���Aa��@g�]��R���!�+�-<��͌�d����r5��M�k��]�IB�2�w�����1RԝLT4����'P��m��K�1N����M쥺�2$^ޛezO�|�H�3�[[u K=��9��1���	�xgB��z�5�f��	�2ߵ�0B�U����HhJ�@q���
�OW]�}Vx~+��\���ED��r	8� � 0�Fs� �o�u�ۉ�l? G�;�Xː]C�N�K���kʼ�K�U6��ř���jP�ųQ;l$9�h��O��1-�����{%���	��Då"�-h�d�u��U��Q|�Z7:<y����yN�@�g}�/X��3}�6�b���Q߱���Bz��t�0��C��#p��:7��.��g�{-�i���/O�R�]X�N�2�:^$��~"3rpк;�!����Qy���c��g� '�^���a!,aga�;�MQ�^�Y,<��-ࢪW�+-U�+7��aJ"��MƢDyDz��O;�A��L�w�Ѻ����_��5b�K��mA�*�F��J�,iZ���n��!
�[<K��t��	V`I�A���*1�+|up����l�$���p����nI�;�V���|!�-�z��D�Ps0�OO��^�!��9�gQ�B�V5�
��=~���8AбBQ�LF�V?��Ɠf0m$��B�����b���;m��Ο+êK��,v�ؽ
*���>؊P�%�f)?I�0�- ��!哤AX�@B��$ޟ~-�>o0�[�)���;�bܥ0?i��4�v|��y'{G�FqK8Gʍ>� ��n/B�8���H]G�g�֏�~�B�Q�G�K�S�bB>%t[�EE��ʙ����\D�-�bHKs����.���Φ�����%f��y;�#�3+��0�h	�iN���C��X�P����<k�8`Wy�3\�j8,�h��� @|,�ٮ�d��Ch�ʀB���;�AQI�g�l9�u�-k�_t�|��Lb�``+Q��Dϙ<Ux�{�S�a��{"���RF1��Q�;A˦_�\h7:�[[jMo�Ärִ���~{���1�P��h�i(������gX���#@�"���:��o��\$����i�>l.&mX]a��7EeT���6������B���h�	�6ZU[�5J���L�$��-fe��9�6Z��"�|9����$R��ΐ
�u�X��ŌV[�i>0O(��c�e2�7O�q��^Ǘ�l������Z�ߴ]y��"�v	�:�ܗH^�Ay�K����d�6�w�K"�B�2��U�&�8����C�]B�r���^,�B!�3�L�]��&�������uʃ"3,�`u��w��M�.m>^�?b�ڈ�ҫ��ziw�9�Sy?	�??(3�Z�h^%�^��C^�d��A^y##i�C��E��m����g�УzՁ��B���{M>�Y���=jG�cgYsI�P�SA<v3��� ������YI��>l���sbϰ�L��̯C���6��\M�⥧�u}�w>M]t4o���]7�!�A���r�K�e̙	��o��	�TS�A �^"�2N@y�#�Si��L�����	���VZeʣ�����C!�����҆��zWF"�WJ�?��#ԯ	�v1O�k�C|RF���6���U�C����7����� �9�3$���f�+z�Y�����'�V��փ��̊pMC]�BJ&����t��d�K���3��Z`�<��� \艝���T��"�={�\
� ��5|�a6Ū���ϞOS�D�����3��8�;=�u�,�=��ՑT�����8cUO��j)A�:&�r 7������	���WL�Nו�Ž<}B��j�����[p�1gs�W�����+Fm��/����g�K�	N��� :œ�/�|�[�)��d�}�3O�j��ȯ�1�k=;|�Ɯ�����wu��JK��Qp�P�mqG	|D�>���R7�NT0:~c��yI-��ƴ9�\��򄠽�OmR���k��2 ���>�YCy��A�{���*`PY���t��YY�yo��F����C�̥��v�\���	
R����m��-3)^/>�\��قg�1ɜ����*lBq�iY$^�:���:�(��1o^7�8��S���O�9`ݹlxY�(נ;�̇=Q�ܒ�P?���7���%s��R��s`j]�d�h��l̓61�s\.�>2�d׭d�#�Hy���K�l�� �I^c�R�K��:%:��Pa	�����sh� I��X>liT�x��9Y��K!j����t��$a"K�Z�N��D3c��xw���b/Cv�����M��Iv��n�.�R�-5���¬H�����U�0N�'�S�G~�?���P�ȸ��h���AP��v$��?��	�<�o?���F��J��r��N�'q�-$z����[T��/����Tч8��0�K^�|ǂK#{`���t�K5p'y�p%�����&���&��U[�/�t��#�?e�w:�1�ˌ	�������נm���x+����ޔ16�-O�t�A8��/؁(�8����kh�N}�v?9����� ">�*ץ��pOh��fj�jL�F�~��c�� =��Zd-ԃ�������y�f-���Z[p�n�:&��+�!��������.#���z� 3�����5׹0
ai���HZ-\.r�U��$�S���}���sS�$���%���T`AXp����C�+1#]�+y�Z���<�&TU�9�������3g�1�6j��<ݴ�,���k3Dޖ�uQ��ݡHHNt�(�a�[����hd�E��Ma�N�\����b��-�v�i�C��=i��Jo\�@��)h���g%2TE�T��"=����X�S,�jE]�Q��&�Ⱦ��3ޅ#a��(��|��3��S�yd_.�RtPE\�Z���No�l`ٍ���k��e?#�� j�V��$�NM<S�&n��2���Xd�1���&{x��)p�?�QĦ�z�+��X��q�rF���v�MB�d��"\G���>
�� ���6*��Z�:г��ߞ�Q�����r&z����pp?q���p�ӑ[lr������q�M9���D�,�Bo�m�%L�;�Q�n^�fI>_����K��;X4��ԚG���ZV�w��#p�I4<�YnYi���tƺݿ3�e�b���~]��Y`��Vd[��Of!�w�����+\+�z�}�݄��o���$:c}�g���9��N X�1M%y<���(I��gO�.:��/��#>��RJ�8�˘��!�ǂ/�M2���=�q8�4oٶ^��Z�����^.�`�J�S|l0|i��N��A�Ǣ�������ϊ*�~�9�f����;�ɾp��,l�P��g�t�5N(t^���i���6����}�U��]ID��Z����=D�c��z���wO[��w}�	Yx�;6�ݱ���˲�և��(�]�X�X����ia�.��j~���rMX�&� �8�!׉���,k�ǯ�ǌ����xLKُV!0xջ���{$,|u��o�/)ؑS(k�ؑ�F��]Rt��e�&?l����l���P���K��ϵ�Fӊ��0m�h����p��׹ķ5�^��y��S`[bOv�)�� ���߼�i������Һ��/� �Ol���h�Ȗ��ӌǫov�����@��`)����>3,�Z��Ԅi�s� ?�_�eq��=#�)��*�ԩe���2+C׵�/`?RW�l�����߃�����s��s�^���>�5��h�<M����0^Jg!���2�Uq��2#��ԥ�1�����Y�<��Z����#ˬ�d'ٸ�$��4x�|��[�gLY�㰝�or���z����]��X�� ǡ9��W �bx`b����%�����$�sK���{�d�"��V��E����~L�4� l�	��GhF�c[w�Uc�4����ŋ�kv���7L��,��O�NL��#�ggSa����\�u��x	 ��^kY1/��-!2�kT!�u����IY�(?b�9��}�)C��� ��2�. 3�5�t~�=�ZJ��.(��%@C��i�� �Y��q�<~����� �1������.��e���|֘!���6M�գ��I�ik�݇CF5�6���2�8���0X�C�t-x�sd�6?w@�P�8Æ��̮��d-�%�e��S#.�d����i���d�B$ț7�t��k��n��N��@��-�r�S��Q�����9�cǷN�����,Ŏ���x���:	Mm��^�E!s�<ʔ`7�?�ͻ���I	�6e��G��p��X򾠮��Ŵ��B�37VC��j�#��g4N�0��`h���jN>��<|�W1�֞^����t]2-��+e�iR>J*
 �u���P'���gu���vO����Ȝ��N�R�g��o��.�u~�a %�hc`:Ve4��$`�O�lಁ"�Ȳ��F�N(��$�g�t��־�
g̑8�é��:�'�L4+G���������If�����GA3�/J�q�g�w+�Y2.����K)z�X�qG��&n��(1�5�	�2{�m�L�U� ����19�I�;�d��u2In��������h�ҳ�Q� p(��(��!8�$1lt��g��ܔw:�$�ȷ��z�ԭ�9��q�zd?2d����|��XkE��u�#�=��K#�5s�ʸ�z�j�҂	jf���#�뼍�;Ux���u����_ߝ�����艦�֪"Bl
,�L���X�
b��	zS��&oAj�'�����Q(�?1��Y���7���3���L�ƶ�L�M�]�uI�,~��YsS���k�*y1j��O�Ъ;z��K@�a��m��i���*9X|*(�����W�������Y�d���oQsEL��Z��uO�����N��(���k����e�d`U��J��H�x�sU1�X*4��h��ڪz[e(JdQqvֹ$�ש�r��������:c��(ԇ���R�A�+B��:�Isx�mp��67�߆��V�/P�%/ڽ4��D��YG���VU$jP�m�r$����egQy��+)�d��u��7��[,�;�S6��,9��΀�G��c�pjK�x�j�`�	�����FV�H��z��N��ER���!�@�@�[��x%��8�K������|�:�X[������e��k8�~���
$�p���N�ʴM�d�f�P� I�5�77��C_�׾(�pϪu�Ɓ���h��=�����b�s��x��.�i�)�2��g��&�x%=(��P�q��Œ(,����7�����A���g�p�d^���7�e\#�A,�N�Lt�+7�-��)ՑJ{��A>�0�A~�c*��DAN`����O�*hS�6��/�z\�^d9xI�������Њh���u@��	K;ĂN/�٭aXQ1�~�U��N����ǕM3x��r�%ʯ�5���f�+����>�u����M7��c�m��Bo���N+�%���j$�y�[�R����T�.������8�h]�;��:�y�y)�7��=F�p1�H�S�z�3�:�a��@�nd`B�N�Ϋ|;��|�?�V�5�'�8?Ǫ%	_M�!CZ�ԀL�V7��s/��P����%[Oȭ�OI�z��jaGU��&?�|Ɇ[��cuj���-Z*��+݂�� ���ܾ炽!�2v�!���b����@��p�Ε>�ԯ4����}���.��'�5e]�y��N�\���)�loV(^+9!�a_A����Ҽ0��`���6x*`��{���Ki����^(��«$A{��*J��Z���Hm"����/�'`.�+���>(%X��4�Wٔ��V������B�ȇ��fs�8 1]��^��q�ě��2��~��Ԇ�Z�4�s����i��`��ݯ7��H+��rF��A����ᕁ�M�ߘ��ʨ��BǤ��Gr���K�q����6�3�rnAb���鯨�y��a6�4;u��(=��:1ˎ�~̱�j_�8��#+;������]�n�����s'&�A@J�	���	����:b�.CrU����t�y|FG'��>�0\-lV{�t�)}��`��su�l�4����Ƴ�T�ߦ3^�׸%�=S8��@� �>�yE��1-��YE��"��Au�g���7l�#�{�d+�u"A�D������A���XPN�V��O��#0�3���Ҿt���W����nL�'[t�{JN8U2N����:+��{������.�d#�ڋd%U�8YVsO�� e4 I��RK�3�Io[�҅��~�p�#���'�K� �Z�@�×M��ëJܼ"B� ~�h��z��tj�QV��� [K���M�Y>.�
�	����m��lyS53 ���'��o��ſUr++��	����+�٥��Lx96d�ؠ�c��^��yi��rޮ��i��/�b�����E�DTc���o���� ��j$��F��7Hl�a� H��A�-�&[�d)V���Ҥ;�]r�4�:Ɯ5��jr˪�\ݹs�kP�0�����������U�H�Q�.���*g���W�Y��Wر�x=���z(�[�����!�FZ{�*M���BNu�� �H�C�M9�2
�f�w`U��]˻�,1m���	<��,�\DBA�|��U����΀�o��]͹wlZ�\�Q$}�#�#v���foq�#&S\VJef�^�d�
QN���S]ġ����dwBu\�:�s��$�A\��t�4yD(n33�F��]5L�҂�źq*�	?��I"�$�@��aF�����%󿳴NP�H�Z��^9_��� ���m]�`�e���!7,��6�rN�q5�r*�6�ȌN�J��=�d�:B�h��a\�/\`c�$:a��Zj�1�� <Ժ���!,2'+��KT��f����o��S��7Ը+��\�ѭ�gf����l�vj�(	���Pԣ�3D��1��9R��5=��i���1�	�%"��Y:��?���!��w;+�/�������ԛΞ�m��$�W|0w��������xA��J�
��c��DP�꠨�3����a�f�]HMKx���V����K��CcS��ln��	QV1)�d�ZcT ���\���a$.��:��k�EA��~���x,�Γ~b�n��1������"��2���#O����.�P����Ϥ��p��5�";��x+���1��3*b��ߐKK��h(�!��8tv���EF�=3v ��.�M�J�.��2�ݔ+�D(��_��
%�~�Q�E4B%17[c���QM��Ļ~��X�[.�Q�"ó��s�Z���NR��w��0�-�B��F��k
����L��,R�H(�Ȑ�ݯ�t����1:��v�;l,d��a~��D�\�'��t�����2,��ېh���D��}�7�Y�?��<�7��T��m��3{Cv��dc��3�:��߻�:��|�Ts�H�h�(焌�Di�T��;��4��8�чF��}�l�-�
bXb&m#D��IO�:ӜJ������m��:0�����&����l��#+<	�eq��֠�c�;H��p���?�V��b�uK�_e��v�T1��?p�*���Tow�'9��׎��W��~؛ �wX�vO�)G��""�+�8�/}g*V�/:�߮u4K!R6�K�J������/�h��	݄V�N���f_� D��̘�{�r�g����S)9���[�PH�ꪊ=��l���;yk�d���Ì����d�����W
��H��CC���r�C��� ��MW�iL�}Ұ�:���k�`m�>�<�l���k�̬�=��f��t��̉.խ�E�+OzH��>�Qޘ�
c�"Ƒbk7�M; V�]�㹍���_��V�����p��LS@�h?������7w���Iu�i���o���,�ס�(��c#�Q'�E�9!��F�^��X���q�0�رwE� N�
��@�`���;�/<ÿ���C�J��M�k�|�qUQ����s?��n;��Y��Vg���\��\'C��������f�Q!�mT���ٿwh�v��:'i�_�T��A�l3��/�a��03\�S��:�l,��-a�1�W�IB���M���'\
�9��]�cU�Rl�*Ksķyq�I&pUqא}�r5l�z��"��8/o�֞��dx���8�����,�|���XI�"��B6eA���1�qzג%_Gc����m�x"��t��U�e�fh�b�d�33�� �ѓ�؍�\Y��P����u��-���Y;ÖH1Qb��o�75���)���X�h��
����y��=�A�a �:|
��W��{����0����Z��Q$Bq���� ��Bo,p]9I Ģ=��E�*��[$ⶪJ� 7jo8��L^'Ej�i�3�z'�2�+��!����D�ǁ$�a�q�i������#O�DU�x?��ӰR�)wz���`��U���\Wم���u�9�:��h%�ׁ/(�N���bYK��nui��ʴ�D��Eʰ1��O��=����.]N��Ĝj�u��*88U����~��Qz��()�����R�ux�-�+PFS�Q]�3�� ��	����:�n�AC(q��\����X%�(A9- L&׷�|U����V?�lX#A��	;(�i�j���������C�E��:2�����a��S�|y�;9��d��{��'��m�@��b�^��c�H�&���`�B	�v���i����Z�ߠ-��y��o�����>%�e~>��@���8��j������&�UO�fAV+��S�{��5������/2��i��d8��[��&�� �D	[���0��Eh��#�`��7k�q�V�zRE.�TJPNq����_k�� *��%���`����'8�#y�/B�w+0�C��m�}L�a�JY<Y ���
��&Bq\D��#S�wX*u�J��G�����:���P4lVܲZ�:��rΜ$�x�B������&��I_n��.G��/���Aoį `�17E��R�۹�r�6Rb�c�y�E>/��H�(w��4Y,�X�7>x���O�Jm��16���4�ʤ��r���a�"d[��^R
�g.d9��^��%[q.X@ �	n����/F�1yU�@dle͔i�����?p���S���;�q+m�_~3�&�1#�	��"���w���׮ #��#E.@F����hl�x���'_��f��ex���:Hf��L�[ht�9�wU,���_�N���W-j����g8]��C5:������Z?{+�Q���	y&��Fm�l%P��Ge�Z��	���v�?�KA%$�~Yp�^�w�'�n���tA;nA8G�!�eL�Z9kq{@֭2�0k�fh[�r����"y�Zl
Vġ-<��pP~I�>��aWO����dݢ�Y]H�X���=��ʎ�`�:�������W�Nt՝D���D�X鵨:C����W���B}tO���{]��j���9�Ǻ�aߖu,�*�-��$��C�D�3ƣ _�m���(�^,?��঎�S�i�Y�XLt� �k�a�FaZG�MU#2����Gd^E�|2Q���/<?;�i��D�Cy���F"�/�-����������-T��Y郏"����8&	�}�,�SO��jO��C���Z@��3$��'����/�7���F,������W%��9�ȍ|I�z�̗��|���b|a�Wp�J�,K�X������Ff�8��]�g���?���" ��Y����'���`��d"��$���vq��0W�%�@���4B�)�93�c������~;���*�\'�}G�w�y�����s"~�����ެP��.����{�"�;~#�̳Dx���m]Ee����P��J�7�n�)��C�)����7��K�:��x�*#�2�ꊖ�m cϡT^��u�l���޳���E,��	je�5�ێ�JC��&�@�C�hllq�`����X���+ �[~Fhx�Zl{
�cs�@�J:8����20����#`�祏�o�ڇ.��p{�B�'���[d@��7�-�i*�YI���K3���r���;?��6�vP�Ķh��$H$��VBqԜ�#{O�4W{�Hȳ8����i����3�@�b-����:�� �����wZ���77�_��|DQP�Q�=m۰��9�j�_�=�yϓ\:3��!�6�%E��=�6^�r��{910e{�5=rH%�g����k*���cYy� ���G�Be'��t��)�������/��kC��H�#	�G��d�R�L�����"�{�o;~��?�'�ӓ��뜊�_�'M��A������ۗZذQR�^[�`�=�c����Bƙ����u�]�nDv	m���#~�i�D�My�$w5����H��/on����E�O��\�n��E�uW���O� 9+L��1�#���8��t�bս�:W��(��g
���e�b����O��_'���p٢���O�&2��b<�p2����a"I����3G���,j���N�z�}��%�	 �%9Ө1�Ңf�nJ x��I=B�V_�K�@������2	�0 �61�F��0X�iz��������V���4c�C���QzPn���F�_��juS�3H�Ĕ"�C~�[~ �Sʜv�k�!��e�G,�����7�e������P9��^��3�ɺ�/vd(~�DJg1\��2�q������ꔿAl��Y�2����n�o�{C�4w�&eш1���D��3��b�Z�p���4��}|������ea<�����u����X�A�k鞜��L��Z%�T���t4�E�'�J��'"���F?�<�v�n�a6%����}��'Y�@�35��]U�����J"M�e�k�e�ͻWs	������cqR:��zn��e�9���������1���ͬ�D�=���\��krՠ��
���"�g���.~䎐������Q��Ȧ/��<hn��ʟ���6���b��a��2�0_�G�h��$&�x��o� L�Cֈ�#��H��3ƇX^b�B��qp�." p�z|��`2����rʕ�Ũ(��C"�s�+��2C���1J��2��#��W�@������s�[�1c��a��,�#?&Z�3��/T��/[(�Tǩ![���ҭM�����o_|���֞�-P�M�����F�A����Uu���tM���ޣRU�̺�2�<j&�)L��������F�}nᮡ�̢PnV����������^D�(bdq�jp�ؽ�8��.f�A�딴C�lC���*��N�.`�Q]+�ŭ��I��4�2�~�����e�q��k�����/>��x�t�j'6���ov ,�{��T�#�	��~0�#(- �klɗW���X�K������U�h��e�ĝ^�4�ҿf��]\�Q~(-�� ˽�d��"�_�T�#�@��f���{�L1�xuFcQ%*�l}�z9�;QM����� �v��q�^����ˠj�����+�5�������ٻ��$��9�F�!+�Փ��h���&b/�Z��tž���߶Y�as��c;�Uw�C�*j��Ó;�#�����5���_8`�,?�G��Q3y�r@Zw�epo�8e���"+�� $�9Z�:\K�(y��$�i �k��.�H�h�X}!��((��R�p��ҵ�j($nq�v��x�˭��/Z�=�K�
��=Go�. N'�~<6�y?���>'9&�w�B�|�aI\��+w�~j���>����>3Ѣ` \��Ԟ�cH*r�Y�[$�Q��;��^�֦�H�����f0��a���DD͉�1��η#���N���߰uR�����$qJ��4��o�� �xٜ����nǋ�W>+�z��&��e>�.[sB�>"9��?EU?>�ЦEAc|��7|9O�H]-ҩ���qk^�O����a��R��%�Cl�j����[�U]vF��ՀT������t4�h˟*8�|�xφN���yъ̽��{)���`%�c�2����߻Puk15O���4��cww/����t>j�@�A�+ե"S���^dx��"o6�w e;��/�q�g)����>&���T:>Z����r\�%�Wx:�?�\�٤*�%󐳋��!,m�j%�>9������Zs��c��-P�����^u�WB��vlA��0<�ʾ� m[�����̴�n`����e$�����P/r�����Е���'+oƊ)�Z�ֱ�	X
��7A9{\���2t���]G��b���Lw���=	���]:�3��aT��t�Ɠ�;hxJ2�%a����{�D:���K6�iɂ/�F_/a�A�"+�����`4��g��I���׏_���nW�$C��:2#MqC{�����P;Gy��Q�!���oy4e����4b�2m���РE8�!����mi�r�2�pٮ�e�:�Me
p�2u"uڇ�ۄ���A(u�p%"�D:g�q&���S�J5�+i��(����m�����;���ʅ��dG�,�.���G"�6���/��e/{~��.�Xk:S���H]�x�kӨ��>+=�>�f
��-���T�~��&��a�N<a� k�b�.C-�1��A�3�m�0x2��8v=�Ͱ�3���VI}�)�]I���%�����t_U�Z{�=o蒂Fq���ui-V6�M��"�"y	�C4oika���~*��]�ĂO��Z�5��E+�L4m5qc�e�"6�m8�>�80������&}���<��`-�[���D?�N1S�bm�\-����s_�#a�U�%R�˦d�$��5�g��k�F�E�T%�9r�zx(O5���>��,���#Ր���C��VT��t���Ȕ��76_�ߞ f+���8�ց~擥�l��n��=�����bٴ��x��@��)S��A�F�H,}6��/�c,>����]�^�Ղ�tJ;*�Aܣ�cXIQ�A�z۽�ݥ�6Fr&#�����;��-��:X�ѳ�?�/��o�ûw���/��nw�gPqr}�G%� $�#����2A=�5	U�֣r_�z��OGx	 �n t��>y����j�H��t��j@������o�,:����3�����2d~��Mk�!��g�҇i�(9��4�;%���~o������ů�_-���G�0y횀8�T��
6��R��}X�>�R�;���t�%��1��ƚ�܀�Y	p��ujw.��QTdբ�Ќ�Ӈ����*fH�������}����<cݛ_p���aS<]���)���մڹ�RF!ty�ϵ�Yu$�>��q\��:9
w�ۨ��?�ʾ��C��B��d��f������#~S�t��X�`p��ڭ^�����߅6Ů��O��@����כp:���q�(�����O�b�u��1�P��yuEu�xU�7A��B�e�¿�sD��5��7��3#��-��5n����B���b��殺�N�t�,,��5�� Tz��["����@�.��͵�aHŕ��֧54�F1 &�y,{E�u4B�ܭ��X��v�AHLM�"+S���;<��Y�J]@�8���ʰB�	Zw���w��ye/:U�~���@�z�s0��ƚ�YFR�5�%�у�THձ��"|�[����M[ɐ�)��ף$.��~�k[H�&�\}t��o��=�=1D�t��u�fSV*κ��<~�n�Q���:����
F��\��l��ĥŉѥw���}�mSV᪘�p=��'��>�
#�������j��J�c�ʹ�Mk���P��an���$��O��LV��>���7Y��n�c�P�@ɹ�&I�;~���)$��ʁ�ikB"�j�P||�{H ��,n.NX�ӭ�eL�Ҭ�KqE�s{�m��W�e^	�!<y!�/�z�$�[�.��oT��ь&������j.�=�_>�I�r@�ɩ�r�乔��uTm���X+^k�f[W)��QAKF6�"(ܑ��{j���+&�S��_��E�6;�����Qh�tp%�S�ڲw��W�c��M!�q4AK}���ۂw�݊A%�b�`q�NK/��嶴[<Ї�JG�������%����K3M�D/���wÒ��ֆl�|��9i�.2�պw�� .ö�!%�-�k�Y��:�avn���O2�/���K{ @8�wAn�Z�}`�So�q���d�}qӕM���XP�Kq��N��Y�9p4O�f�y[z��yB�@�G�Ӹr����	Ĳ~��Z�>I����e'������͊��G�ܠ-�J1`P@ ��Kyh�#����?R7�<�@�f������=����'^Z%=Y͵�5�����֖ai�DPr��%1���i7�2�2Jɶ�>�35U�sW�������Kl�Zo7�(��T��}'| ��Va���@|d�t���������i"A���dm��(M^-�MU��Hc����@� �(���P��e&�I��Z�]iJ�2&T��ܼ�̼�H��h!9�<�o�ڍhN	(9�Yװ./��=LΓg����zӨ?ؗ��e��9<.��ۼ ��+>��o`�σ���-/��Ù)NiL��$��+�c74����+�"��!���9`Ob*���$x��H��Ok{ic,�/!��g����o5[��}V�'0��#�{�_-K�`�p`�R [�B�^��k]����io�INx��IX /���v��%������}������6�� 1�Z+��y��mЦ+ߚ*<�}�����0���:�K�Խ��9>��Nn?a�s�Ћۢ�xߡ�>�qک@�/M8hY����$�~�3o��e�h�>,܋Ր��j�a�]��t��#ᛯR��h��"����-R2T���[��E	��\֠�;0gqf���,*�宁�/=G>�y�g��:ФR�lYb�o�DH�񘾐`j��F�ha�F,���ٯ��mX����qPúGw��`!�X	B����}F�b҇��g�[�û9�k>���b�v�Wڳ0�h�lACZ\�3���k�<�Z�K���5j������˹%(�7]s��o��8�'����l.��e���18�rxT`��l�m��rr��$9���B��e�  mK2JI��.t
���b�$�ѷ�/
���,{��ՠ�M��gS��i�4�_�[C�#)0JG�_��w
0Ic+ x���`�B�����G�R"z�ev��!�
����#������7:���~Q�Ў��%�𗊒{���=�
�x|9s�]p�X��S� ��x�)���j�	���do�E�EĬu�\-�*����I�Gb�d�'�k�ڍ�T�R�FY�3��.�|�������O�]7��K����1�%����[W��Z��C|V6v���4C�Ȭ$R�sV�;��LՂ')�9h���GǶKnx͢r�Ā�ψ��z��i2��o)p���|.���Аc��vޫ�ک.;Ɲ��6��&I� `3�ʀI �D�$�����V��\�9j�	��@|:�,�J�`�U �!细�'C��#��U��IĻ{4���',�L��@*��R��=T�\�����k����xl`aB�H#6Q�)��Z	\���"R�w��'Q��&Gܣ�X���}-*���WH� ���8�P�5�܈Pk	 c��-��X�_�~�k��r]���p�4��kE�m��G�ƿ�_� dR��\�"�(�
 sS\P��g
b�?�_��~`=�{N��ލt~&k)�dC�G�Ҡ�+��HOz852����<����=D�%(Km�+��/�B�4����!�7���#�r)�W��R}�63�a{�|�� U�	�]	6�(��)��qV��`Σ�/�+Ms:%��F�LnH�Ό�qI��T�9BRz�F��f���ņ�IӊU�bp>V�j?�o-(Ķ�>he	��`�2�#Sȝo<g5W�n��E�4C�,�F��)nU6zU�	>j
��䶑,=`,�@r<
���o��&͜��̧Je��F�A��5���6Z�ˣF�,�X�'uy�[����`��=}�\�J�c+eЦ(���쥢�����'�*���E��b.��ƿ��^�=)� ��k��	؎�yk��d�;�q�t͛��l�ٞ�!�L�׭[� t� )ȁc6s�z�^�I�`|�x�t�2>�� `�$��5+�V�C��!����������8Y���ӧ���V�V��%�=<'�@�WkWk�%�)dZ��/�]��~�,�;�v�{�'�w���^� `+�Gp|h��kĪ�W�2�O�W�Q� [^X�4�V��H�}vzЙX��Z(�h`� �� "��������l�l �@�9�����t��w�1�#�1��V6�&����v-e�'�c����� ��L��2M��RX��ޜj�-���a�pݷZ{����ǉ��h5�:O�G=������E�Θʽ�=}������*���Ɣ|���j�����7'U��ߓWI���<�tg
3�A�/5����J'�J5ܙpR�Rթ ���9&iS6�ź�.ä�߮B' �U�M�+x� X_��Nu�)��`��` <� �j�S�P����Zp��"+A���sMae4#U�t�q�M`NȰ�a[_��2��^�kxx:�䨛c�lޙֱ�3��/��@�����~w���������xz��Zl�,PAv6�	gW���;ܦ�Gxmq�G�!�b�L�&���%TY�P�up��4O	��`A�߲���x�H��}W����Ŝ��D�FQ���8k�d��mW��xg�W�lԸ�Tac��3v%b8����%�Asf���w�[���zXE��(˔Z&\�����^����t�Q˳!r��y/h^ 
%8�4Cg��;[��+W�W���U��-��F^ŭc���"�)�b1�Rej-N�����p��e�U�-������Q�v0��-��r���^�	���b��ϝ��I�u��)�cm�I�x�y�5J���~�����UԪ�4���Ң��h*�]W�5f����J���s�dX��o-�J}ϵ�ݿ����Z��l|
�N�"l��t?�D	͑%�!��T�{}���͉����T^ƫ�E���O�_d.�}a���:a��۠�04��}n�n�y�B��b����u�d�����1��%h��a�?�������-p�+�q� ��+��0of�8Q�?�W�DT�vU����6��'����١d�?�%�������_�Py7�D�U����{��C�xDKyK������D�`��	�0�7�N9�P�p�����?N�vr/D:�K��{����?�kb*��I�em'�J�>���ؘw־B���Tm������{s��0�suUדW�a�M�F��N�&(aZOCBƾ�.Bg�1GW.'2R70�=�~Nޫ3�1W	��(t��w?�p�e�͖L���4	����>�G���[s[I�?
�(ݔ�)+��$V�F��!�SFۑ�Au�m��H٨>ͽ�8"�?��S�TVÉ��)*!�Y��o���÷��/��0;|0g���NH����} rU�{��
�Y���+(#ꢺ
ac��b�5Qʶ�y�\��n�L�� @��S)�Y>|�l%�(v 4��It��E�̉����sQV�C��62I�lL�FJ���,�^ڪ�M �h��߳�`cV�ߓD�r;sWr���0	%�Q^�Ϛ-P�V�ȉL}W�\��=3d�6�|��<�_T-�B�}~x�ϔE6%�h�LЫ��rg�oR�&�^�=~XZ���l\uɍ��k�3�L�?��-S����ņ"A�
k�D��Fe�עGC��j�$ �~)��6/V�F�G��fG���ޅ�!�P������Wm̲u�H����k����A}���U� z�(�}����0I��m{4����p�C�_��K�ӍOp�DZ"��4 -�8��ppkΈ�/�5��a�4a|4+n��g|�v�Kr��T~��6	��7�����d��=��@#�9F�*J}oP1X�F-�6���hV���O����Y7	O��L�������c������B�
b�̈5��˚'b$m�|5ЋGs
f	�u�I9���/����`㽝׸��n ��a�3\��xV���2>�z���\�(أn3���JՠAk��"�VbC{v?�S�1�?ח;��i��r��-�	z��r���U�u���/��a���B/�йa���n%�L�g�K��y銷�X�P�ځ�Ɔ~�mbL=x���{:�ze̷�I$�d5��+��e:G���?��=́�]�_m�<�~+Y�pp�c�l�զ��.��q6ė/q�N ��x�Se�h��.�]��.%�V<��A�!gl���M@��\6v0Q�tY���4���"��$)A;�ǮK��t����)����nt��Mz�טc�t�P�!��vD�nX�iήC����Lh��ە�H��ghgj�V����*o5�z�7^���[�����pb�f���J�|<i%xQ� IA�?��^���������W�$�hS�
�ݚ�.xO2�73�D�;���~�YwGB��+���{��C��� $満��S{2I�f�{ӵr�B�)x�B[���m<C�3`�5�\��,-�/���D[��\�d�O�V�i�s������~���#��Ǹ�?<m�<@5�-��&C���Gb>�>����W���`��� ��)����\T�C�[�n�?��_� �t�+p
�i(���sz��[x���8/Q
�E/Z�2�\���EJ���%�0Qb#1��5⳦���{mV���w.�f��a�O�L��Ю�L�����sQT�n~	��m���5�����=�%���Ѷ��=��m�s�Vw��y�;{�:JZ�&�%������������p��뙇AF]ϣ� ��f�u��y�2�S�b֠�_zm��/*�<�g��̼�-���Af���ɭɅa��$��!��O嶂v����(~<�}��х�����c���W��4BrV���� ��}�h(K��Vc#<!��C�� ygF�=H����=n̂�Mw��#5Tt�c�m�76�u|g��=� M����ݰ��)��v]�&������Ey=ꏭ��#9�Z8)��*�p`|$�䛾�J��!���з�ˀ`�>�7+��o�Y2"�17��D�y��^��)����i����F���3��'���Ey��
������N���_���B��4]4��2����C�����M��	��Kh��7���[	��2��xB�\~�&Xx�����&3�D�x����&�4P�G�k���j?�n��QTCTme@��HLf��1;���9�"Y�H�N'=��m�&��N����(�JO�v�����I[I�)�(�
'Hz��<=>q�2���n=�m�����N |�T����O�-ik)}@��.��n��pi�,�@�	��tbmoۚ>����ʕ�2�jM4�|�9K
_��Bc��?+�x���u����C���5P(�Nt�V�C�G�k/��]���@E���)X6���D�6�����Zq�p:H�*'DK:�i�"K�pc@�J;8X%N���*8��(�;I�!Q��'�r=l��sj$Zj�/�[4���ŏ����X���q,!�A�f &3����S�S}~��ǱGXY|�D>����f|s˟#Mw��s�y��7Q��WZ���.������\��=�ԚB6�L�Hq��7p�KX��l�O~R4j�V� #�mUL 2��K$'*r��bG:������j_��̭�Po��{��F�rv,7�L3����b��0$�o�1�@�H{���H.9�p���+M�v	��"Fk�Y���w�P?��F�Oa�C�^T���u�ş�*���6҆YJV���:�l��=wٌwͬ�;>��ˮ�
_�>�2^���w�n���G�˝t�d8�F�����~��=^�bN@+�&�K���
�`֠&4�0"�����ɏ��xl#ާ3p̂�$U2Oٷ�^���v�3���XL���?~�����|�*H���o��-Cp�<��@[J���q�7��؜~m;�1����@��^4��]K���R�эF�N��z��C\R����g����u���6����"��/+��e\��%��D_�x�3�v�,ϝ̪A9�/��1��=�៪��Q08���ȾG$_-��@�l\����`����ܛ�Y�(}��څ��(?[\4!���msZ]5X��������4�Z�R�W?A�~<0��@(H��9���0Q�l~r��JР�RE�� ��7W;e�
&>N� �|]h����Z����%�ͬ�jk����.�-�?+5Nr��� 䗍�5�G��C�����9wq�S���j�)�������������d��:w�=ql�iM��+4�����R��CP�,owi�K��ËE���}����'��H
��gO���7�� /;�͢z~�ހv@cg�X��:S�V��<�(��5��~�2^��&4pD ��B\�%r�?._o"�Mwty�B�c{D��ejJu��9r<��ݼ�[&�e��(ݢy��O�
��&�	?��[��R��k��ɔ� r7�i�Y�CveM@��e~������&�Kg��!�қ��oθ��=L�>B�Wn[� �V�����]��F��kz�Ů�����?�L�7"�Jt��d���J|�i��.HLñ^*��>�7G5���&厐.^�%����ȥ��ק����ܗ>�N�!7((�*Ŷ��O�U.=�s<2��A^��$�oM�����d�=����~��+�A_��+}�?�r~�q�� �x�P�Xf���M8�{0��A[r�4�}I�i��A�Ƚ=��8��g���5�i��u����V'�,L0�R�>��<�%�wd�2�/P�����<Ŷ��X
I�]p#@�s�ɇ-Tmʃ03�N5!;��}٘`�U���n\�;0�VW�jc���O�p�MG*�����G�����4c�-jZ���#�M�C�6������.qs3Ėz�ҋ�J���ǔ,r+㏰���������˖9Ϗ�^�^�ޕg��g��^	���I��M7�~�1wZ�3�ܱ����r��T6�CI�M5����s����6����V�Yǎ����#b6ո-�̒��;ׁz]�d�T0؂ϸ�W0��\�����@��M��<��K���0�����]4�@������~	��0��9�ꋻ!,���Y@7k��#P.�����+E2f�/wy_�O��Mx�˨C�k���Q1���\8�jy$��en���}Pbծ���Fj���4���ˉO={Л�[�� ?Q�+14��!|�V�G��}��B�'[�Usd����m~iW}�����%��Ga�Lx����]�"ʫ�N��BۜS��X�`�笩Vq�����| ��7c𕊲@�T�	�f��&
�|�A��0��5��9���+=�5�e��D9�t<�������1�[=�gs�u~�:���L���b`	_�T��3u�'""��z�O��U0OK2����M"��J�#_�=d�JvC���YK�.�lQkD�Mp_m���ܐg�V�}wzI����-_�V��n�ִޝ��Ã1t�p���`�
������	B-�$R�'�<�g 2�}���L�hp#: ��(�%����rϛ^#�&^���\��t��HlB�TQ�O��������"��zu�-��;����E��37���b�b�Mn�8k~r��Kw.Q_�c�a&�ߦi	�b¬�(���B��&8��ߧ-�+�u\%?�\2f��4�1�8[�����]�K�^��0���Yxn��N1P�)E�'�S�8�=f6�2�`l\���yY��N87�r֐^9�$L"Pf��w�"/����2�
�c�9�ʇ��q;ɾ�T91���C�^���?��v�������FU�� �3#_�FS_���y�^Ck����a�����?�v{��sV��wao�8E�x�jge+Z�N��ܵ�����I?�J��o��!�IĬ!�N�
f�8bJ�\��	�}#4W(�g�� �:�#����Xj���D��mas�l�`9c!��l�E��n��)�t>�L;������vM�3���;T©��)i��N����H/˥!�����i q/�->� ӎ,O�W��T�+��Ϡ{F�Ι�äm+5�QBF:��ȃ5QH��P-c'H�q6OF#�(�W�:�k�2�d"�%U�_�Z�Wd�vQU��,(���ׂP5�OD�u��ۼ �N���o����
օ�$����dԔA�˦%�cziO�)��/>|e���������<P�8���NT!�F"�>M��"h���H �ӍSw�_�&	E��<�5�H��-j#�j�q&�4m��	�;���a�'l��'$��}q�y�ew����o5�[,����1�2҇'�s!���!��|-6q�YkH��y��������-Z]&Qx������� ���_3�g_G�Y��҅����Je"}G�KC�FO`t,U=ң�E�M�WS���������<�O2��	��:#��._��[>�'	�9��������\��"��Z����P�)�c<�E�4������0������z��Y�5�5lD�l[ڦTc��	�*2�;\�c�R^��.ݭ�.�����!U�H@I��[�f�]�J��o((����vr��-���'�An��J��)�"4����!"\s.~j����=gl9�V���̐=�=`�:��J�2΁���rcc�L�@��f�K��l��*����S��a�������>g�s�w�,�6e�)�� �U���Y�g�������I81����r������03�~�%���C�T�HbB!���PȖu��f��I&�ٽ��*�{�w�(�X�h��kH��a�#�bm�eS�!y㽦�L��C?K: ��U=����}����Y���I��oޖy$�X{}r��{��/c���Q�Gݹ*�E��[�G:�nD�߉���r���̣m ;������M�\_OSHRl���J�`r��
�7n�*9��id�Tt��B���<�z�y�*�^3���双�r�����\Knr����Ӛ�0� ��}�o�"3���f��_���=���,�zO���}s��؁6��H`�l��m���t���e���P�jt�s��ө��!͐(��&�����r��r3'$��k�{I)*
>�i�'�.fһ��58r\����'�D����
��ZE�_�/���AH,PE_�{[�\��<��о������f��K�׵���f��Bک�Ҍ�^�lz��h�*E���s����e��O�_���d0P��It�,q��0�%B����A;�zʃ�ڰu��*�P��l�<�=�������YF�򾩝G��j����È&�x�;�������g���=A�~HTG�����J����ę�r�^˖��H~҅Z�c>k7|�o��{����+�A�^|�OC�_��%t�1�~%���T���Eɟx����ɵ���Ո�:7�É��u�j�z�0uo�,vC����4�./R 'z�<Ǎ�� ��o-]=��DNěHR�o��V�`,��+ve�bHx�e�x.d�!q(c�	[ƶ��>d��3#��-SF��m7��Z��F����^�ю�lz�`6X�%��0��H˂� +��[�g�V_lzNY��~�kT�^p���>�m�����N�C�;K(#u}/�����T����ݑ����
��*�%S,�ubC��T����e~��$u�B�خ�>�PߏKW�P���",�Xxf�8p+n#�%��b�zې	W@P5�^�d~R��uk�C(��#��z�_H� �Hy`7W����oO��4�!�}��s�G�q�U���,�_���~�U�G�o�V7]8�ś���M��]ш��#��p�,�2��W��e�;�:��2�G�*�
<&*Q�Ldlg��J,Hh��I����b�ݫ5�cb�ڥ,��}�O��cࠪk;q��#H\����S�Uv�U9]����������]-�,�A9hU��\F��J�٥?X�8��X����������%�G�*�6�����Ӹ/p.@�`1t9�V����37�c?������5�4J�H+�5`4^@ڻ�\V�}Y��^�d�\���=����b�O�O�wP�Y}��A�xf��P�t�^rc����;|=K�bˠ�$�>kE� �g�/�'�l`��ڦ�F��Fr"̚{��{7�O��DGM�6�Q�~�-7a�ۮ,i0�ۗ��1ȹ�7Q�d./ؤӹz�Dd�2�y쉛�T����d���Zΰ���{H��ѤM�5g1]��0s��~.�tDo��_�y��UNE=���!�%N��_�LӶ��>�9C����wB�x�e䎻��w�2_<�b�I�i�I�ny�)�M�>
<�C@*�z�d���4w'��o��վ[|�M ���>3�ی!�x���ܛ6 sj�[�뎱dŐok(���i��+l�m���eH-�5t{'4�\�[��p�-_d�d�Z�wk��~�5{|IU;|�h�	��R�}l,��Ŗ�C��7�S��(KF����m��_�s%����BۜQy�����^0���!}�@��#c��=4>���x\�2Dx]��߆�|0N��t�5JG#����ӆ�&¯�^V2���R��6Ba�w��riE�E�N:�̌����W�2E�+���{��C�������4��q٭<�h��l�q�n�E&]�(@^�YoS�N	��&:(zV�h�|,���n?�ǔ�e�pij�*�63#���hn;�^9�5-qN��Qt>��gd0��b��M<��P�ԣW~);�Ԫ���o�ai���N7��g9�ץ�W��,q�X��7�4�1(Ijr��О��i��R{�vODg��!�Po/�\�t"9�$�T�9��؊��D��X��Y��%:��2��h�FV�y�˭�áj`c�p�WV��hG��a~�$?�o�˄"]4�Ҹ�B�ZG ���x95S��~�;Vaj�a$D�,A�%dg;����(�$ڪm�e�c�}�ޑ��ަ��^�It����Ў>;�?u�D�Iq�b?ȑ���>���{IS����5r�I#�����	�H�±��F�=dd���b��DV+_��*35�"T'!�N��B "���ڋX�3���g<��Z{x=6����EX��k:��J�&���Z+	�q�q�þ��%M�Q�������Y,�w���:���jeWw|Q�c�C%�M �l@�u����^U��J� ��g��I�����D<='�gWf�Z�哼u�����E����S(&k-��J��N0ih%ͮ���V����2���!żAn#�v�}���{��~��%���H3v����oVy�w��>A�O���z��ޛ.������3zj3㵑��Bp��6�\H�E�c�.��Kr�b��4�D`�"� en�d3t�Mp�&ޖ�2R�2U�K����H]�pg E�c�)7q�4^�
WG�aw�m��R�<���#7J_s@��A����0s�*��.� �Z���fRk�O�ԘV�)F��Xן���X��蠳7j�"f��D�u��In=Ԏ�1��^��	x�1&H��f����e˴�|�1/t�#2��f/
��,MW�ϋ��]Д�_'=�3Llu7:�_;������k.�{bאIL�kL�����rhD�]�mg:WV���إ�xƱ�+��r~\�H2B^�!� 8+.r)��D���.*bRu�CC�S�Ha���j��[P�2��z��"���8��M�-}�J-��>"I�_���6���[ˊ������#��C�9a�[Hp����A�Ӧ��+���(ã�����%�J���+�0�Ņ[�x~A��-�և��t���5�����zŰK�~0m�R>'�G~Y6e�Ge L;(,��@�P�E�݃������#�L����}(��/S��ty�p�7�����@��v �$vˍ��I��)�i��T@���B�@x1�ρ�m�ƨ� {<?�*��^D#��0��V�l5��O������2.'\}�q���H˄CL� n 
7�ݳ����2��yT���x�>���܅qud�<ô� �Wnz���q��C6�|�65�[�ciS���i���1�ս�����rs
��h�QU��f�I�O��Wy�����~D<�š��+\�Z�I1>�cxv�$����w�Xi�� s�(G��W�G� m�1B<�M���[J���L��~(����%�̰��cH����S}��.Y��<9 @���i J7�<Jb�7��9���y��St��X�և J�=BSv�:��g�)�5^<a���{}���EX#�5C��̼�W�cǜ�MM��Q�6��Ȯs��Y�����5��}_']��.�v}xpܟƋH�ؿU*w���y�i��7b�.�3����A�lp{I@�RQ�!��У�ßE���6E9�[E1�y�C��U�P�T� d�^.(����Rj��5���A�֟֓-F�ǵ�`��ګ8�nN��#yoL�zw�����S�a}�^rU]'ő�ޯ�2O�n�gM�)Os���B�ڔ�=����Qx���bJ"I!�^?����(�Q�;�&G*�@�sѵ��i{X��W�����Ǌ�+���
*�O�=�DePK`�H�S�����V4��_��
u�X��$���"�1S�|���a��:g��t�N>bM�s!W�#?�T%[��ڙ�Λ_��K]����.D���~�W�yKԇ��4����i�A/�Y�"��'rR�9�2�d_�6���N�NݯH�����?!C�`]���(�\�Ԭl���L���d��&��sY�]�{�{:��_��;��仓h�xu����d=���N9��4X�r�S엏"��&]]Ȍ�A�Uw�;pe��o{��~v ��rx%r\zLB��6�R��S�NK��)�*���5~���)W��`�J8TCY��K��+�s{y���͇z���<Z�r�.�~�p��Th/G-Re�H�;u�4�����*��{Tw��W[�\�Y�`����R.��|��1g��J��Jh�����z�## d8��ˑ=�L�F�(����[��@��4y9�wv����$Z�-��l e�.2�'��	W{�s�˖\�\�2A�@7ru8DN�6���'�;��kב�GK硾)���c_I�&`�K��kԒ���������5Y�c��߈^ъGH�\.՟�S9q.DNЭ��0UK{�G��q�����Y°��1t�ӥ���"<*z�!2��@ƭ�;�s*F��]���ш��{�Ш�bځn��p�Y�-��o�Q�����}>>G"Si�UV�@���B1JB�;ìq_�T�8�� ���'{��k�iۘN�O�^��dlψOc�gږ2E����G$ ��}!�o�
��8�b�GI�A��n��85�'��e�`�͡� &��0� [���F�%ޞPW���EW�p4�6��v�@0���qo_h}rnTD�����l�:�ş�|�$��;�^P��
�RIm�ܼ$�b'���-��,8g�럒�߆lwذ�˭u�)� �ʡ 3����D�oR����"���hi+� ��֖�o{��� %ێ��wў�q=�>W�9\�q��Ucj%���Wh�2���'�\�%4�Z�6��J�N�
{w'H�DR�}S���$H���sF�B{�4��y�������HBun�C�]�V��7���ӡ�&܍�����$p�4�3-�O�j��*��d�3���J 81������V�&���g�gE���)zTt��o����5T�D�]f�V�BV�-`V��H��P���9��q,]p��>�\9So�ŧ@we(�1@H��+���3�X:v��V�x�;T�t��Ou� /��|��� 2H�7�B�����ңo�4yT&oF�B���f|�oNIm�����/��&�.Y3IcO���JF��`��~}_*�"[Y�~�3�,�G�!]{P��3�yz����ec�Z8��)�sƧ�v>�����=�Xc&�B�jo�3O��!�H�F;?[� ������!���ǋ��Q�\�}��(���tT:�42`�gG�\W�U��0ؙ���cr�?zrM���7HD�߯��N��;�>�^�n�������������=��at�'�A@l�6:�J�GSxg�vp�g�����8$�:B:���"?c�^�c�mf����/�0��H2 )��tR�EW��(f�j!c�.1��������,]̡�ӝ��)שH��=�}����s*�����L_2u���e7~��#Ѻ� M��}C̦�/ysڒ�ܤ�%�-�S����RwxC��В��
��B��>�-��ؗ��k7{o ��5�"L���VR��ɲ����+�\8b��e/D��r{h�ۍ�BU��H$+*�h|���L����n��%v3���,6q��s���Z�#�7t־�8?V{�����A?�ȳ�Q��̎��q�m�����0���p���A���zw�qvⳝ2`8"W�\�Nӄ�m�>�o����=]w��b�{�K�;R�e��245� +,�ra�*Q�7o�]Ph����V�,�05�n�,��J�uG�M�$������9�������K�v���w��7�P������I�jLD{*� ֞��3kʄU߽i�Дս�G�_�F����!ɹ���ُD/	i�]�J\�a�Z�l2xF$���"��`!)��p^���
<'L���*�83
Yӝ|E/t��u�hV�լ�r܃�2�}��ʑk=8�&����O�2L�Ł�-V<E
��=/�L?�K�3Fe��[V�=�߯-��u�_>�'2%"�bM�r�_�n�QJIf5�¢�;��[�;�� �*VC6����*�T�w芻z;Q���6_	y��5�Obl��j�!N�T�Rf{��"ذ-PzM��W�-𛪘'��v��/��u��B������K�Ή��ظd���+��uD�F�)�$2�������l
��rR��=)as�f	�I�u�m0���� |�F�� IVwf���{�7TΆ�+6��2���9x� �o�� �[�L�v<c;L�2��E)I���[M�2X���\�0s�kZ̏A;�{���xn��èc��@��8�6�Qf,	��|~�h�ܦ��Þ�+j��Nua҈4�3w�nC�l�J�.~ɾ���!'���������w��ۉ�r���L2L�P�(4��9E}V*�c��3������$���-0�=�p���]�Σ��8ƓI�|�z��J�?�Ծ��C�=���CR�=p�����J���IL��d���dg�}ɱ;��a �/Q�=��Ҳ;��S�e =%9��(Ub� ����f�H������o�����P�>g,�G-��;H��d����O�����s�������c_��������d�b�M�����GI���Ro��6z�Ӷ��qT!�)~�a)\zåOs#��������oL����
/γ|0����
Fo��>����;W�4Z���I��s�(?��]�j�r]�������E5� q ����-7ɋ6�[���惚LϑsgF ZŐ#�5#Cx��rHS��7JO�ܙ�:�cǊG��RG&z��|Z�����XmL�v�AV����B*�(ܲ�1�{O�0�u�ت���*������]�mK^��W�r1S~��"��cA�g���g����Q�|�������cW��ϸ�@���t�!�Y��e�G�C�U�{wA��Bz6u_b�Ή��"�0�,�aE�Я�w�ٻF�^4O���U�^�AQ�{hc�v�D�������|igb�e�a��k����t
�f� �f���7=z��N��ɸ��E��F���:<ʰ��i>�\1j�ޡ��U��x��&���8�1�hm���3�+���d:t�rU�,���-���t�;�v2��?�a'h?%�&�N�����8��d�X��h�e�Z�d:V����K�=�[����N�	@�4��J�-߇j��E� ����L�� g�Rb!a�X� t��<f�-�� ��j�iK������ސC���r=�o���t�:�ME1�#D�,
�n?�����$)�|��L���j�2�����	NI��	�cW�P���%��uܟ�*���{��૔N���`m�V�\'R�m5��RI��a���p/��%�i^�0z�I8
���#��5�V. ����"���KZa�%R��R�e7'j�,�E����6U�X���G	�3�{����
-d7ʃPg8U$�6�BZYy�b��!����;U��AJ�k.G8O������Lθs)�x��z���1uG4�oɔ�w����e�p lf�k{�THk�
L5�$:��lv=���HR�N�v3Ps�S���&R�D�aB��x��1Ip���v�P?����1*4�X��S^����עCu�NI��X���K^H}����tӧ:f>xn²��\�X��K��2�څ��H �RA��3��r<���*Da�x�[B����������Ԣ����$ɳ�Og�K�������l��8/�`�0�c[�Z?`'�l���Q/���¯�C
�ۧD.����u;��&�+=cݚ4�Vvdp����>�8����@�U,�w�>L䫮R��ٳ�c��M =ޏ0�Ͼ�+'�xt���4��je��M�Æ���t���W��G1;m��Sk�u��zw�8���N�W��9�A>غ��=�ǯ泔��<�U�#��\8�S2�rO�l�@�%�P��%�&p��Oq'rP��c�5��f��Q[�D~t�7�-7׬���d3Ğ(wn&ސ7�3��U����Z��,9�AY�9]S�M�`YJ����럟��P��w>;Gf	"�8<)?�"8��rŢ�zijwbg��1N�o��3uN|Aɢ��ˣ��B��g�c��rS���Q�3�*�A�;�3f���k�$��G4��5����MS�%��l�^C��Y��h�NǙzI�K��̱Hc��K���	�~��w�B��d�b�w�l�^���l)d#
�`��a2�����=ɷDtj�=lun���Qm ��i@Q2�l $�S�\ޑ�2N�뿡�� C��D�x���}>3r�=_���'{���0D�<�^@���u���D�_��h9���@g~�2><[yߵ�p	>~��f����?��G�A�=��g�r�)�w�V����4(�%,<�8ϔ
F�T6>�+�楠�e����V"�M+���q���᷻� i�[\�3��FM:��H(������n��)j
G;_d�YAA<���N3B3{����|i��h�=2�8S��\R2�љ|�%>MA�Rm��� �=���;��W��'2]p����F�[XK�-S���$��؅���!�	S�Խ˧x(�+�D��,| W��Y)Y�A���H@ƶ/I�a02"�;~->X���˖0?�z*Ҝ����NJ(�w�Ԗ��E�(�l�~�sğ�O2�XY�h�4�#E��ĵ9#�>bM�>'{�F�&��߬h1<|�:ϛ���W��S/'��BǱ��1n���$C\й�x��y�	 ��m�]�!��1H�$,z3򼦬M��3?�1.ap^��T@!��rb�C����K����9�J5+:��rU&Igb���>��W �@�"���!�W<	�[OzO�9�`q'+�l ��܆�TXmݽ�5}*��KZNg?Q� c5���<�1��n���o����V)U�rz�E�$C�R*��$�&��L��VF�1�;��e����vW�I>L�|P��D�s�r�����6(��Վ�o�^/��a�>La��:�ZM�7�@śQ��1BܕS9^�� �.MQ���i�v�)�J�[�&�;�@�]0��`ԟD �Z�������VA���d0�wL�2cN^O�r9��*�:�|th�t��c~�z��F%���bŒ`$��c�o�p�"@d�n���$�Ϝўem~��C��jK��0����
���:�}G;@��:�y��١���ݹv�ɒ�xS��x8&VՊ2o�¼j��y�^�I׻�w8`{zUOo�b�s|ج��O�KkG�}�a�Z��i�� a�e�Y��NS��S�Ogo��p������1̋��+V�kX�
�4΁��hq��}_t�)����"��;��҆�}Jc�O���4�7G6����S>�Aq{D�А�ž�NUݬ��ҕ��U��Yr<����T�4u�8��e��/�7Ox�{ J��{��̞�f�P��q����]�m��Yi�m_�R�g�F~�} w��!������6x��ٖ!��/ ܪ6�셔못b��B�_l� ���<F:��҈��E×�A�8!5�������jH��v�:ͫax�ĂBӂ��E��N[͌�P�1��ep�p�N�s���^�Ͻs����c3�:�9�M�Hlي�S��H~2���a��7�}��am&�x�G��L�Y��e�=�M���gg��uԏԇ�]�u���EWǳQ�Ӛ�A�{���F�8Z�9��
eNQ���
��I�����r~j�*�S��?6��R�P�Ұ6�����3��-{9&�߻a��M� ӽ�~�źm]׺�XPN�s����ջǥ$�`�� �>n
M�����C�5	'���ց&
#������9�7!����{"���M{���5BL�*ޔ�o`��FkQ�y{G�Z
��2�Z�NB�]�0F�n�*��	���|���<7�F�����=������  =���ſ�8oX4�H@��1k��ML���#8�Q���>�{����l�j��n�r|'_	Wo�yã�1M�K_������3˯iu���XA�G�5 vwF/Z��iq9b�p�n�'S�1Å,�,�%��?��2kN�q0"���'o�vImX��o9�	sg�	r�Q=w�3�����- I�V~�v�K_t�Չ 0HjEf�91�E]��K�.d,@¸�hvsQ�*d��~1�w����+����P��;���
HeP��g7I�)�ӹˎ.<��B�z+2��N����������kQ���40���'Ҁ�qX�+���Y�Cgr8�.Am�z��¸�_��T�R���3�*�o�c�Ô��H*�v�������p\�\=��9� E�d�u�X�g OlU⹦��/��������g(5d�d9}��}�4'��TS�sBY�Y<VXg��!�#�#y)��1o�r�y���k�:7�YG��!P�K��c��/��1
K�
	��/�T)����}ˇp8��K�Ǚ7_]��E�J����)f���>�G��$;,�����ypJ� �	U,w����d�V�9)�������EL˟��#��{ܤ3�Bf���FX��s�VN�b,ߣ8�Q��%�	�s�dT]7�<�F���'P[��b�5�d<3L�|3b���/�2m-�/ܶ5Cf`��AWphϟ�G0"W��X͑␑��,��j�F�I���~.�7����M���ۣ�S�&)D�r�G<�����x80:	<���[FIF����>�HAkJh7ص���K6�JAexYȜK�����k�@ѳ���5�`]�Z����o�?�B�v������K\��Ңl�Q<\����PwD��A����!��P�0��4$�uϿ�J}D��	��%`���/ʄJ�8B���:�9����5j؈�cG��׬AM;U��f���#��������ƽSoa��s��B��Ƥ�0��|	t0*���S�3��!�3KVx����D����0����q�� a!k6�����s>��8���i"u�YȵYZ}^;�Z�`?k��a�"������5ى�I����-n�S����gT ��� .��v�~Zc�v;s�lif�:���VF������:�#��TP����w�-*4���$����Ij�IS�*O�N�c�w2Wy/W69O��2�@ÌQ�=�s,�2$0��M[$�.��)��ф+���n/�?A[���<���<r�I��M��Ǫ*b����Q��ѭ#�fY���X�ʿ��U�6��`�@bɲ�=
;�">99�-@�P�ǵ/�3�=e�6bRs��8��B��������N�u�����t�^�������,І�5�1���^����\+�Z��b�9�����0l���Ua<��A	���N��ȝsfxE��_����i�K�v��b��^*5�T7�ax�J��nL�M����ABov���Ha�Ǳ���B�����=ϴ���B�qxP��:�;C����h�?����N|��e-]bM�8��v	Ԅ}e"̨M����T�ͷI���V�])������h���&���P~5:5�D!��%����_8��お;X($���b�����H���<���uٹ�h��@V�T�_T�o�{վ�yK��ӄ`*z��j�V� �8�Y��	�{jv�«َ�Fz06�]�i��\Y�	l�`0�L�J�h]+D���3��݁Ln����:�n������޺΍c<��v�(��c�!��/���L?�rLj�mn���GM ә�on}�x%�L۲Ϭ*dƔf4��}e���rV�����P�56]� G�E�~���P��f����1��|����F��#F͍��s�g�����~�j�	P�{�!Ks�f?p�A���M��?�#�u�q������1���r����=�df�ti�ީO�����/:�Ud���CK�>�������(�حco���9x-��u��7ᔒm�-^�<^�����ZgxS6���c6�c��J�^*�]4��9i��N`p�P��J�%m,J���o �T�"�@B��8BO�ɔPY��A6V�=wh��լ2V�7n�y`8:���T���M���������xݥ�Pr�ʾ�LP��X�K���d�TK��8`TT4�[(�iz�.&���0��ioc��u3�_|Y����7�Sd��#�M�����ʈm����i���1?�M��@���_8�ܭCCU�}�sO�Ni�<�"ym�a{Xm0�f�x�C9�.{e�H����`�Y��$P^^\��p�J5y{�KE�k�i.K����:C��ˍ.��f�ADg��q�B�z<NK�������(�l��um.����¶L��a�DOt�.;v:'�gH���J��{�L��) �k�`�����9�����95R?�~��z��8�G9XI���мG,8�E-g�B���F	ė	�������DN^Xb���j��m��p����%�U�nw�=� I(=�މ�e~�2� ���Ѧ<:�x�r��r��Ǟ>��l�G��P��'o�TIp�*Jd򲨉�M�4�_(���L=!�����e �Al��[t��ҟ3.��@��q��YG��%b��[�պr�wz���<.��t�4YID�,k*�����t_%sy��Zǎt����PupV<Ҫ_�þ0��a��Yg�����}B�Q�2�}���wg���������g0��b�Gڇ?S�a����[��n�C�cl����h3<}�E��ta��Du�����_i�g�-ӬN �l�hԪ>�\�/C�O��Q9+/3��^v�w�rD����%=��q��?�Xg�<W~Z���i/�����S���`��M58�O��3�զ�?+�D�<Z���*C�w?d'Z���+��vYvnm��y��$�����r�b��fܠ���%�
?ֹ ��N��(�<�Y�z�"ƥ���JS��R� �����?b>Ą�M $�H��A�i"
��W$�9�)������i%�����;sz�U��ÍA�J�J4J0�1�	�[���N��ق���R�N����$�l�`�8���L�4�@1����hm�O3��(�|Ӏ\�l����%z5F��^@�A8o2-E��P�㯹g�]8l�����?P�9��Ǽ��K���HBk~$�[=��&�_�
5�o��xxLK{+�F��n��D
CEHb�V�3~�bЖ�D/֍2.���!��n�Ns��^�&mY��eV@!DN(���.j��6�q���(�v����ߐ?v$/���L)2��SS;uz��ڊ�3n9Z���i�/xu�3�v։������Ǉ��h�z�����؛����I�eS�ܭÞ�:��\���Ĉ�Pr�Hf�%�%l�q�&^ ��S@yG�*м�0�Z]{��/��f:P��*B�j+��/*�,Ry8�LbUr����,��x !�D�?92���P�Y�U�֦.�o�\�2k��3�BR7�kͱf{1��Rs�>?�J�w�/]�zg�z����c%I�>A(@���}*>�*��R�䖾h:�s�я1qaQ���є�I,��l�6�sno������f�,�$�,бM�!���w㱿R9hnkf��j���6w�g��$2hD����PF��΅%=�g7 (^$�c@����ٖl��jp��||k3��:ͨ�YI?��$�+��_3ޖfm��!R>�b�*g��0��+̗N"��K��v]U��X'��� �7BX���5����{Oca����O��)j�2nz��(�����fڷ7q����b.�Č�\�L��Z$����]�e,9��T, (hY�
 *���F�F�q��V�,�� v�:��벫[��0=+��0��iFH֘:t�@��<��wΔ�֒.ߺ=!��|2-5�Q\>���5 [��ր� &�+���\�y�5�
㙇���W1:0q��)D��h�Y!o�k�5*:�ʻ@v�s�G%���"���{}�j,���>Њ`�1����ЮO�>BaA=�86�b��
��=��Eh0H����>|.^�>�$���0{�[5aY#!_�*�N�kEB���Tf�N��o'��r[���;2��������w1��~�rw��-�X��]!�}�T]e�!N��[�)��Q؍P�|�dA�dM/������A�Ζ��5�4Y1,�k�v�F�ju#`��QȽ�F:�a�q��͈w�^�{���r�L��� ��a���҆!�äO�u˾���K	�ZA�*��e�1�.!��X|�1C��,D�U�1�w��*����������ߤ�&Sᨃ�w9}�<�.{e����$�q���EX���^M�l2��s2k���(�8�����ښfn�ߧg��~�U3��*,������B��(e�����^@+�
��f��ڊ�elBX:���$��d�JCx��ci�q���S��-�{�S��r��m���T}2q�fLH���J���70fB��^4E��vlV߶4'�4o�@�a�(�va�g`v�sA����:B���H�¼�/�c+�H��y�^F)�ZJ?����mEG!��gV�3%b(2������?�~��W�5�}���mǍL��/����&�͖e� �h޵��{��O%����L�~o2�LPݢ&���j�3}�c����/�R-a���.��d���u�$��������n=G���E5`6��$�>�5O`�A,�o�Df'����G�!�i�c(X	R�3�"Ut˓_a�u��k���n�?����Ī[���6�
���4��YP���1o/�
�0}�(@l߰�y
T��Ŝ��N���
�I}�cx�x<"�o:p�r*�J�D���?KG$��1�����J~������i%[����+X\j8E�$�Y빘
)�S�5�nӈ��4yq�ѹy�̝��Q�~O����E(��N�gKDeq&.F֍9��~�
�v��M���9�j���zd|~��2 �X��jo�`�nD�y��Gk���/I�1V�N��n��v��FV�ل���g��¹�t�|^�օ��QJ�+DP� {ןQz����ɽ<C��Wj�I5��&t�`B,s���T�:49�F/�˘�#.�-/j���� ���afp�aC�pa�K�aR�J�n;4A���6����D���o;�l����X��� ��u_�Ch��$#��42�)Trf�����	�&�?{̓=V��p����>g�L�`L}��O�(Z��>5aJ���j��UJ���g���:o��=dT^�T�euIt�OB5R��7���(�ʘ?jb(�^r��DђM���k�~-R���H�I��T�xt0�kI��d
S�MF��17�+��ln~/c��~!D�w����!F����2uY�9���U�.�7�~~���^'@ܱ �J�ںd��S�C�y��k���L:%m0 t�D_w;8�0��Ր�I�+#�z����`5��R궗r�T�Q�$#֫���uF>k��PQ/}��Mt���φ=\v�s��.rw��p>蓢�����bQ5��g��r�hr�-!�18`�⠏"���ر@/��{�i �Ì�A�a��H�<?���<�	�Q�qv�$�RE~s�J����ABob ;��oN�vK�ݢe��ѽ]6l��|F��OMN�XQ��Sv&�$'���<t����\5%y�%ޫ��C� ����49�����Eȱ�.%uNS�z>��s ?��/�M����D��c�dD�lZ�Yza2.� ��}�8q�5�#���ݘ��e�4��CwrU�:�}4���\Tڢ±�]�{;! �Y��zY��%��k_��l �>4��n�5�Eß�{���3L��|b⑎��2��b���g�i�wp�MF&�BY�,�f�9׎d��R�x�>6\�peQT 2�y����i��,Lh�i�)!Ԏ3�s�T��k�t���x���jZr(}$�BbȦ�= Dcs48�BH$����_�2�"��c���0j�!9J&b ^�kT	F�*��G*����t������ǍhD�0�77,���a~�Nǔ���)E+��q��ƈ�Q%E�����s��u<�����#|��}\�xneG�IK�|��ضR��ͦ�TNx�&�<X���~1��ځw}�i�n�fQ��;��eH�l��W7���ㆃ!�`DK���A���q�8�tj���~�w��f�E~쐾|����_t�	)6����r;������T,��ʀ�%���ll	e�O�hU(������.����cI�����@�U1���A!�uMH<7��o5�瑩�~����'Q�*S��
r���aa��dꄑ���M�3}u���uL��(Jj$-\�6���A�t{�5����@Y?�|:���j�n