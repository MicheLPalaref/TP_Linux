��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�x}��j��S�b_�)F�1�(d'Â,L.��ꙺ��e�˭'�{���)�Ilf\�@,�y��Z�n�X�D�P��c�����=���]Od�w��yD.΃��o�gc�5HFJU��d�܉<41�]�j�Y����SǷ�~U&�=�h3?3-y(���Dç���a�h��Zq@B?8��dM�u��<�4ҁK橢ŬV��\C��X�����i�+5����r����(��<�3�@1>��
���$-�}r*�\���	�DR�����&*��	]��E���Z �j���A��^�vz��@W�܊��B�f��7$u�A}��Y~|�ѝۊ����DH���i��hx���RJ>g��|�&�`��X�蹕b�vDB��@K�7���ܪ�B��ܼ�K� ���������ˁ߱�>�Ҟ+�莪��;�	�H�*��<�!��ML���� d�rY���=I�?��wX.$̀�o�HoS���:�κ0'j��b]�B�M�%!��x�yE	>V�������%�z��g�D>t]��U��_�U�)s�t���}���&�����r�Jz��J1���y��%�P#/����%��2o�)lr�����Ƅx�Ĩ	M���Ч8��Z�+(�����!I�*�<���!���|���jtSo���B�9_+n�f������҂R�Y�#2��V���Z��
٣/ ~bD(}��	Z�e������s1 ���$��+��p;ތ�L��ؐH-���$�4
�{N��h��(��7Z <��.�7�q���>��w%$���(u�J)Wm���`��{�{$|{c���#؟U���ҳ�� R���c�h�8#/��HA��A�/����t3ա���.g�;5A��j�p����l���no-�JP��A�R���V��{��o��:S
y�#XJ�m}0J��$�~��`��ƞC�ʆ�zp�?�����)���v�c�	�_�ٳO�z�Lfy��Q~���	>Ց�s��3A�̬�t�f1L�~Mӿ�	�����Pm�{�;�������@�å�����k�2���]�/��4/����ׇp�"$8�^�w��Mj�~�`�j�	B�����"{�x��k��S~$�w�G	g�I\��/���&."�<���9�?>|���s5��- <IH�.�>��߇��uo���9�]��+��w�z�W_���׾��_Շ�lW^he�9�j/`�ch�M,q|ݶ��ce &���`��IԵu"�CN'z�ܵ�>I��9� �W�����6��^��m+y�VWAr��Ϛ��U�]��$��A����%�
�HϸϠ�g�cS.���q����ek���E��l1�����.w'=�,Zf=�#��i����9�]��2;���U#Ѕ5�����YӁ�O���ujc3�1�,3�$-2��UZ̲��)R��C��O����Q$�?k%�4�Yl���au�xsC1!� �l	m��HӇ$^�\?b9e\q�ϵ
SY�~M����J23��yOZ�q��)/ɑce���I��e�%48z��ki��伆�;��k"�p��H䁾.#�X��6��SW�r��C�<Cߑ唔h�g�<)B�e?�d_5��E�*�P�ߴY�z	�]0N��'e����@-�pLRəʏ�e�Ζܠ�b.0B�������#9<4҅��\4t�7-��p�BD[�D{�S.C�t>�I�`R$XNx���zݦo�[R�6��w(�\|9�h���\ǯL+8��O���*�� *R�<(�R|#'�ړŠj�-���Y�6�lz�HZ���N�R���Vw��.�L�(;��hD	G���if�·����7�(7t�a��1\���/��M�����ga�/N"2S�ώ�Q��y�}H�A�W��+HVte[��c����)�K����~�0t���O�\$h�����>���Tnp9$� �م��	Ph�ߤ^�<�Qx9�Ѭ�4��=��yC#r�rv��צ���$��p~ِ��� O��>��9�Ǔ�$mЃFW���A�k�:�J��ߘ�է\���ڙw^�iζ�o7D�ku6S��D�)���p�|��L��:�0��Y��2��|pC�Ջ�R����CK�-Q��Ò�>e����m)�D�KP;���FRQ8����3W(��-:\��
���6�����(�M��ZJ �z��]
,���A0����������`�����f]�]A���P����F��2��Gg���4��:|���	"P|qsd"�����j��p��X'o�z�Q"0�Z�զ����ʛ�Uذ�?��7���X���lڬ��ރJj�!4���sa�6Vs�U\P��W�c�	pQdR+� ��m��ܭ��q�
#��s��F�9E�9�9���B�����55�G�*�������=g�����G����j��'�����2)EZ���¬'�<	̃�&��w�e|�Ns�	#��  i��)y^�.C�(��e���2�<��CYaX#M�� �Z`%�z
��P��eAJ�F܉�e!pb�)�B,�k\Тx����ͽ�a��3{&�)���~s�T�Z�OMm�����ù�Z����M�Adj���'�7�C��kBh�9�p��{3��8o��z�W}N	6���s]\!�l�L�o�AA�%	��f��� �t��970Y����̆@߷ [&P 
���@	|�-_NL�r�D�-�P�E4���]��y���h<?S�����Bզ�e!��c�n�͓:��p&d�Q���R؉�C��ۈ��I)�j�\R�Th���5�>m4������F�Y�|KK���f+�V��~|\�#��~$�6�%)���!rl-%�t�q7�G@_*Ţ�����d�HǬjϵ��ԁ#��?��z"�hw$�=��6@�{݌�������Ra'����y�G�u��ٞ��Cr�LX�&�9�mY�Q�s,�X�`��VSm���Gf��d�(��Z  �.�?� 5����g
�TvC��V�)y'��R�@�,$/���x���*A����PB-THc��d3���hʸ �S��н"�vե�X���~��ks`
�b�>���ќ����\<��%���'+�0ڷ5��{��_mS\b�����v_YK-������O�ÕY�G�I5r¿QH��}>N�!���Z�s�9�km��a����`r=���/q�7�?O�5iU�A�<<���)�QWxګ\ 6���=j��w�_r.ȞR{�˵��Y��gpԞ-S��:�'������H�t�+��M�!�G�\eVKS�U%$�V��t�Ϣ��ǲ�(y|�ZƳ����:��`-���4�~��穮)Q�⑮�N�v���D��xG���t�R3�#O8Z�ܢ�t�΃q�/V�9����` ���~�>�h��G"�s�
4�&e/�a�	�z����������K�bE�a&���5_���`w�7e/�y�����=�#���b�
�`�2�?�&*M)��qI���)�fbNǽo�I�y�l����(�v�I��%������U�|���t4@���G3N���(�{���ڢ�뙺0��v��9O��[�NN,�dT�|�QgZV�A���p�}����5��6����C���[p�e[VAvb�Po���G �Gy��ey��B���+�Q%�ͫ����ij:�FA��d��-��_���n����o���I��ץoDB��V�H��B�'�w"�FܨR�I[�&1����Í���ްtP�{َr��Pz<�	��"<C����t� �1M�z�K��Q
�c�g*�h�1����O8z1�D�.�s�b�,.�c��ȴ��--#A~w�l��eZ?g�iQ$��[ ����5d(�dZ��m�k�K5���o!ȵs7� �u�u!榇l�����s"�"nVr��+]�E�#N�)�j�4]I�(_��W�DaI]l��]�%E�w^�xa/p��{9�B@��`���ΠPT�u�Ck��'��i ��xo{nʶ�$����sT��>\�i�Y,@�@	ӈM�v*���n��LA7�QdnNg�Uş���j���T�3G�G
@'9y���h𤟒�N���Dݗ$Z|k�y��!�q�ksd�@	��L��HL_�����9�axK�K�/��s��U��V3'4";���(�QZ���*c�(����ye��c�t ���5j��*2h|�}� ��n�z<Ti�Q�7�:'Eq7|�[�j�L;0�}~��u}�N��w��k���S�Dq�u���졜I����������MF3$��Z��El�b��x�����|�����A��0&e��ƙgi���NB�fJ\AQ��xL9,�q���lA~�D��lY�^��R�{��� ���F8�d��gf�S�#����0ب��5X��5� [�zk%��7*��-؟�#)@�u�^�|����7z�����XU��g/l{����c��om��~�p�*QlB��6�n։[i8"���e��D�ݒJ��ww7�Fe~ǝ&:J�dR��E?T�H~�d�!�a�E��2��D6�?�sXFqv��>�On�&�q?��q���4zt,�s�k�g���}s%u�-#zҪ�$m	��*�&�l�؟�
|�B��km��|1�/;��E1�j�n]������x5��X�<�q���7�,'�l�c�e�e��徬-/:3�C(	�5� t�� Ӛ��1�%�����p��z��zb�&��jLfP֮G�<�0'Z#�����W�U�$]A�vDQ���Q������d��1Y�> cL~G�-��3�51W�n���,�w��M�X�85a�����I��:XjI�a(�����"����$aMϷ5���a���&��J ��S+g>3بDU� �nnE�vie��$�(o- CVo�$\�;[�͘虽���G����D�j~"ܲ�n�lU-��ߔ>�J-�w�o�8��Ԙ�=��L��+��QHO~�E�o�1�����9[���M`5\E'i�"��K?�B�����v���`ӆ^Cv�-�?��e���/�8�_�[��D�@��a!�9��V&'�{c�+�KZ��ݦ���}}��a���H�N�&�O^82�,Oq#rb\�_,�:mc�Sg\���S*+��~]�3���)XKi*��Z��r�m��+��0-+�����Z�1�����uc]>�����;moQ���}���h�L�rLkjQ�Nl3,,b�کy��m���/����ɶhh�/ȳ��" ��K�@ҕ=�����myԅ��&\Y{xaL���T�]�J���Ox�)�h�$��e����F:��l�c���f���1�M����(
�h��c� 1猷\��H3� Fc�m�K����N	K�;1��¬c�?�~w�07(���LPR�-W�C�^8�F�͟PU�Ϲ��������yDo���(�D-.�T�t)--D��Լ��V��B�t��RC��łi� ��I�SQ�G Zw��( ���K�w�����_'�}	s<jJ9ޒo��r_�+�����d8�]�n�_c8M��"������mO�Y1�O�Ut�5�2�Ӻ>:�����`��>HJ���^yG��ƀG/y�>���P�a֎Tw�?y�ʚa��-Lp�&�|G�q��?,�r��w�eW������r�@��� H(hM��b�H枣ajwc��j����\�S�N��T�;�$9�Z?�?+��+�6�Q���tp��u�-i�L(��!FQw*�~,�wEBњ�l����ɢ��H��!�V�h�3��銊X����J�O��\5��_���j��-T6�-l|�]32u��� P�^��7�v/<{=��W�é��l��=q�Px��?�؜$����׷���Ѿ;GO����x c��*�۸J\Q�_��+�T�Ƃ�I�*�:V��:e�|TA>*JQ/�L
|Ɇ�;F>"��k3A���J�*Ԍg�����H��M�c�������i����ClEm��O��&M/#�O-''`q��1�۾�=��\]�tߥeڮs)�G�@h1�������E�?���G�fO��6�� ��O6k���	��;.��m�S��J��<���
��|9������+�U:�[�?����գS�v'~��Ǐ���+��+���S��^F�{�u��V��2w�QQj�!]���U�!�y �I~$��#_�>����cY���b�H��ņg�B��o(�ɫD�"�}���cHp�	��_dx���&��H��Oū<�VL�9�� K���@�P��uۮo�+= (b!�\Fx1ג��>�a�%)��ǔ�Zo�N��X�NƟ�rb����F�\j��?���h�*�[�U�7I*]�R �;����_3b3c���8A3�V��wԵ�t����t�ae��\>3~�s:�A�c@�B����X���O.�$9KV���	ҏ�:�e&���?�J����᳆'�P��uL�}MiMj@6J�*�R�`R����c�:Yʧld�[�5��ۗ((!��9ݹ���Ύ�C��V^�JjO|K8��+3�?��g�P�|��ƀ���v�'��(U�����M�=���$�|��q!/��Ⲝ�~��pF�>��*٠��N}ca	�Kg@%E+>�!��
V�8��15	'�1C�3���&��ÿqi��S�z�Q��	��ۋ�^��G��x4b7�5(R��4��ݯ�y˱�>�F����N�{M�C�\���wmű�����n,��Ks�?�A�Pj�Z��)mO���;xU�T����v�q��"*am������zIČSf~N�B�[�2ٴ�p��CO����+Z�4-�"����Rs�~)o���J�$�
�[�&}�{}�X�����!��/� ���tW@qm(4\~�֜����.X��d�;��������kf���N��&�܃>i�����Ε��e8�����z�Y8'����h���S����4�X�������	��p��N�����]#mV���[ʢ�� ���k�}<pKe��H9Z"��)�֥qkk�a������C�bP,�m���:B�$���<(4*��ĉ�\�_�r�I'z�i�"�׎� {��]m��e�4��կ�d�qͳ+��~�ldWag�	:��L56cv�
��`�/���o"'�$.TX�����96���ɣ#��
���M<)�Ih�	'J �&[�z�Y��E�ʫy�;���������Դ��@�tv�v�&0&������A����ӏ+��G�)^M����Ȣ9+����F�;9�+i)���8B� ��\�m����J
�(�qx�B���lAdϓ���F��%���ǌ*P�8GUi��5;Y)��h��w�.��N�Ζ��� ͎��Dt�X���[5!O��L#���<'���d���O��f�|љ���1�h�k#r�y>ai�UMn$�v���ZD��6e;|M[*,ɵ��<�E�F�&��e8��!jW�7]��^��k��P�)�Om=�~l�i ���i�]Q]� �Qs6���r�vu�_P�#$y��G�N�Ŋp��w�w��58���;�y�Fr��ċr;���ǻ�;�U�:�].�&I97�:A���n5Û���H�}�Lג�_�;�����m�߹�9�Q�7鰃ߞ�^����������gi�3���&f�-��/W
Kh����Y��+e+`4���8�`D�����U��ʑ )'��<V���|]7kj�\uh��8~g�o:���B�K�s#i��>��4�n�H�)�X����,����zC�u]M��\�K����b��t	�1]�W,ffi��mWN.̔���˱���<TQ�K����0Thg7fWtDHYn�ȍ`�i����W��h��m�|�#ww�v���rp��u�̨� ����k���gx��'�r57��:��*��BF.=�YA*h	��!ȥ��y@PZ@�[����[͇E2�yt���cvoπB��@�T���7�_�ӜL��.�`*��߬����6�
���D�0�^�����bՍR���u��;�����V_:u$��^
�jS�K�`�Jvbp�[�8�};T��/��g���T�KӭK�협~ z%�o���3Y` �@s�4�澭���N�zl��������o�)L��UD:PU6�m�P��!X����'Ƒq<8�1y	�q�F�j��k��PO4�O�ڐ�3�Y&��c�VV����)X�ޑ*6�C.s��%��'�☟b>�3��ˇ�n��:��:�sb<˟�UG�� ��HbSk�of��G����A�߉��"���������IL--B� ��;��h֓)�@��K������M������ӃV��Dk��t�0Iȧu8�}�!!?]G�H�G
YN�[�^��@)2�6I,�y�e��@�<�0�O��+�\Z�������LT��0��/�������*r>��z��-�sRQLE� D��hWD�p��Q<�����Sb�v�[b4��B��Z4-�(&��[�>�},;I��'<�j�q�.�p���tO8���E7(�pq{/��QNE���.�bͣc�19��y_4��~��U�4���㉠Ki�gb�<n.�Ч]�����kt����L��zLV<�7�4��e�9�@Р�u"t^�L�д
��%hOF�h?7��.>.D�D�y��ܘ�7��s���"2�ˎ����P�hx��p@�bF�=v+9�E)�t4�9Yxs>�͕l�@�t)\r�rWU��.���.���kB9q�s��3���9L!.[խ��W�Ln�릁�O��N�U�}���UT��|�7�i�\I�A�-l|���.��87�?]Ӿ��b��he?�%�2�_{x��J�t�|���Pl���%�ɽ*�� ��Z�����u/߉���/��<�`��S�r�l���:�L��)���܎�΁��#y^� ^��ݠn�6LY9ԷưD��%�����a�X�Y�uH
f�Ӎ����&��>�H	���`d8>xT[��\����4��k�q�L���ˆ�jL�K��{E�aRh,Qk+Ŀ��f���ώ�VE�*A��n�5� <Ȕ��&�QЊ)��r�&��O��'K�q��:��i���y���0j�ܑ�!�f��q���8�Uq"¤�fP�%��q�wͼ` ��8@X�T0�)·{�M~��OG��F��M��J�+S+=S��(�U��[>��-= 31F�or�`
i��WOf3��t��=AP$��h��q���e�ι��tn]�����k����a��})/n9q�.���A@cѬ�|�ւio�"hQ8\�F��#w������<����w����ї�݈����x=2�["��>s��,Ӵh�n�S~�a��s}��lO��?�J����mP@�óGg�RG)=����B/s~b*����Qݺ�������! ��v�?eH�� 	ܘ����4���"��P�݈�(O���(毝tn�cW�i���` �����)#O��$��)SfL��RRV��Z�O�3���u����~����6\�%��Ҟ��@����5��4V�O7�hB��{���@���Ѝ����XV�=w���gT���%�G_*��#p���'}��$��"=-q���mL��Nmnj�WH���S���=1�#��Wo}�:-�pg��_��s�h r����-!�|���4$sRô#9K�	N/�&�`����|mt�>Lp���+ȁ��h1���,�7ʑ#����.%-�� ���;3>�����e�Ny��Q�|�6!��#��<�Ʊ�v�L
�H?I��A��B$��_X��hM��w��+�T�(�Yv�ܙ����J��٫@�I�^�#MB��٭p��"��!�~��o�ٸ�Y�Ҽ箮݈���wWA�>��y��¹���q5V1�E�L�2�F���K6 Jo���������`�Zϖ��e�'�Z,'� � C*�3z����A����� :�/��Ik�Kh���t�vl���Ā߿����]�.�h/��d\�`.����5��s�dg�r�2G25T}�|G�:y/UW�l(vv�9Pe���u��W߅UVW\eDF���T	��R:�6z��?ZJF�;��u}	���פ�*ܧY�B�f�R�ͅg:�<8l��Q4�l�,9�(��"����_>�p��8}2)�?�e���	���е�H����"�eT������K�O-O���B���''�3�a�Yx�r��ya:�.A�Q�v��OUz���ފx.�/����/��]��R��8��������oe�""S��#�<x�j�T .����Ϟ����� !_�wt�� 1 WH��A���F��ߔ�=/�'gx�	^����d&�T	E��v�yg����Cc���no�L�Bf�m�'}�heb�!NX���$�(\�����c���W�Nį�Rә	%�?�UR�&h�Fӣ�+C��5���:f}�$���&�}d%��� o%�ԇ{�K�?~��m��.��|���(�͜�a��~��"y/�nq���Evka!H �9�w�\><�b�j��t������ֽ��0�xq�g�.��"��5�a��иp�Nh���L݁�t�ݎ�2�<�բ�̛�Z<��]7v�J�]�S4Mf-�a�vo��B�S�:�M�5���8I��G�!�{���$Z�5 ίIn��e<���K�
z+�/����ɀ$�/*�����K�r̯ə����v�O�rSE�BL-i*� �����*������$î$)i@Vs۴�.L��<���3l��(��i �~�=>~�_��M(�X�迚�ak��0�?Q�*�