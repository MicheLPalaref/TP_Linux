��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW��3��+�M|�Qb"+��#�g?	t<�	��M/<��eg;���B�`}Mh�0^F
1��<%��a6�t?�n�+�hX�o>�AJkG�iQI���*@)������f��%�~D�����ӘFy��P�1�ɂa���*4ŭ�7��(j��B�v�>?��^.Y$�G��C�t�?��Vć:�`���UC\~>��������&��_�}�S�ˆ���9}��c�9��-'��:|F>|A�\
;_9�/������3=K=�
�1����ʎ[���ʂ��4�گ�I����P�t�{�
#Pr�Sm�Q(ۣ�IOKD�#	{Mc�ԏ�N{���)�Sߠ){���W�	#{�!��]Y� Ɇ�3(���:��A�	�r��ޯ/�J.�n�O �1ޔx��4!����BL�[�-&���0�p�����a2T�)��9h�Ew%1l����������sq����Y��GR��������x�W{�J�g��;��V�dX�WY�DZ$~�M��y�Fm�Ln�x3c�:�D�Sn6�рy8�s�nA�y~�
û�+هcC����2�;�N�
X��#䁙����b�pa�$p��"��͊	>6�V3�E�LC{����UH��XR���t�H��g/�Q�+C����k�J:y
0V�%b�7˪�f@��m��Ǘ�ˁW1/Z��<ʁE������_��d��R�v#��.)�Oi�8ʚ�H#TǟOFj��ĥɽ���Z4P���/_��5���h��8ig?Xf-H�xJ\�=����H�@��%������-F�+��b�Ϳ/�.l���I$pN' �'��+����<]�Tȸ�$�Tϓ�Yd�g��;3�MP5���Pt(|H���ߖ>�W�j[��6��_�9L/`�* EA_�+�yN��qB^ �A�|[^|"H'��Y��+�8h���lN�r�[�$d��h~����7��p�Rە��`�/e�#QwE���o�JQa����ƀ��E"�4�8�D]�,�y�v!��9Ƈ|j��B�o:G/�Ta��ھ��Qtc׻0J�I�J�n��ߍr�_�L-���gqg^@N��k�iնM���$Ӷק|��#�����S��R���{U8�i�;�hVͺ��n��x�h���̷��5�6�kj�{�'M$$��-i�Q��=�*_3�A�p�9�~��h;!�4�niT�XTz�=��(����i�ܽ�b�,���KN�1s�O�|9����� �4r����Yѐ���B�E?k)ʡ"���Q�8]遼��	��WSJ$�=<G��;��c�fV�M(��ܡ}B/n8���J�_gi�KW�#� )�	���͑"��	 ���@_0'��\�`i�"$�Z7-����d'%�曯p�#y�H���$Ey� o]:���`]-�G#���N���8�W�}�R=��J��=��:����׷W�����W��e"�R\��?�M����X�IQO��b�>��5�J����{1�8h�ߏn���3�|II���ք:Y�X|�ߎOK�R��n�������]rlM�%��<��lp!!{m{�'���hj�0Lr���[f|b����P�:|��!���K�Z¥.o�:h�I��o��ڲ)}�ރ��:�b�NRT3�x'EhR��u�'�V�꺆ZϲS_�O^zQv�a5+kV�^w 5<g�-i�r�]eNg�t0�V�	���U�F�9	zU��`G�N!�ej��g4�r��:dl�dU�be I��i�D6i�|�p�Ν!�̯.���l�x�t/-��fr��(9�� �I�`$�&"a��&�ꗹu�n� dp�t<	����{\�XJ�B~����@��\��Ae�@�������'�2�|Y@J�����m���۱	>L���$���o�.�M͒�����2cBR2`rI%��ߔ���!��}X�$K���J���'�?���@qe��α�3hiQ�s��a�2k��8,�F��m�1��/X��^�^9�_$��r�� �J޶9<��������3�.��E6�4��q�I���壺?d�V���],� ]*���6:���ƉN��*]�y]Q�백r�'P�o���O7�L��ʽmƦ�|d�jS�2aC^�bT��^|MT�B��%�:�>�>X�	K�3N�*`�hT֑=����&�9Th���M���p4�%e���z_q��t�mg?��1�;U,IB��3$��]?��E�H�Z��T�7{�DTE�7k\�laZ��d�{���.��fy�P��j .f��N�6_P6ż̟��/o]�7�7S�&OQc��:�$涡�#N>�� /�\p�j��D�[��U�I��im�8ofǘ�۲B+6�]���yU����7�U��h����4J�B�_y��B����k��ĉ�-�d�ۅ'�i��6��#��2�W�ǰ��i���Q�˳@"�0�Ē.�1�۠]_��N����A~��)c���A����ܾ�K�����&�5c�i���f�A2d\��}�-�=G%���:�^�d�.d<!���e.D�̖/H/�W���5%���D/͡�)*,���a�v e7>��������T�_z��X �Gg�r;�,;��=�>�'��a�g-N J{��.����Պ�r�_�{��M�!a��4��Ã ����x!X����n�.f���[�� �n��a�:��d��\���ֿ7헟���"�+�D�W3�~:�w�B�5A��Hٳǹ� ����Ꝼ�h�L.����
�g��O4�L|.x��VC�p�[]���C)�
Ԑp��_�B�p��Ƃ�H%/�8���^�r@ރ�'�3���V�cˢ))�������n�Ϯ���͙�l>��q���]>��d���RI{�2jx0/�x~65e�%@�R��94��� �2]�a�Lo�'�}1ib �r��&�lI��@~��o��l4�{b����֣�O�=<��N��hL/:�k8:�L�o�x��� F!�Ub̅�ݧ
��#g�(��z�#-P3�2�P��`�$:�iD�zG�K�N^9O�N�yvzB� a<����?�$��I���͢+���:�:�I�,��oį�(b&6]ec �,��j�#�@�2l��5�๫��ia?�݄�Λ�Z�72��2>���d@䓂(U�i�jѲ,#J�Y~e��^/d�眊�äL�#'��(�tIZz�,[Q�C��B@���wP�Y��%[O��a�$H�C<�����%UV
Ec˶��$�&��@����?��+80��v J0l_/o'l�U=i��f�.TB�@���~���K{����'|�)>�p�K�%�|I��W���P)S�#^�zS+s7.Ϋ����4��<�]p�J�z+A�� T�u��̌�����hTD<�&���ko�����rݨTG/	^v`<�C�FV��h_ZVO�CÀp�����m�؎�%����ߨ��B~�Gx��&Տ��&>�Z�ף��ϞҚ�'�X�e�f�1�Q��� ʧ_��[&i!�g%Dr��'Ѻ�E({�G�2�5��#֭��5!Aav����ǜie��s��R�֬������k&K��g;(�_��Kt�,�&����7�_��g�Y�j�����h��6U�����\��Ʊ�ݼ�����Wm�y�m#`]ī�JPLzu.ny`�A��q[y�=(J��i|��4��c4�U�f(U���5�$�v�^��@�����g*����g�j�t�R�e�X���x���Ũh=x�T�C�>��0ً�]EKl1���P�}�	9_!%O���"�Y�q�|[t�;'G�ۛ�$;�h;#N2��CY�j�7�d�p���\��&����OY�z�_�	�z۬��� ��G�=��6kӠ@�I4[���KZou��"Z_����n��xӐAT|�j{*j/�iۜtB͋` �i����8b����e�J1��	��F�S��UkAb }�o��~(B�eh��'M���<��PP+��&�-4�Kg3��h>~\fȆ����rl��5 xӮOB��e���: ��4~;�>ɨJ�݂oxbE�_�hY��_���R^�E>	E���`;�����b�� ��	+�����V�T���6���y�0wc��΅��-�����F�Q���@��6ݙhf�-�H��N�	5�G���Õ�dz�(�G�e��F��6��ͦ8�}���a.S�o]�^���$��M&ea��_ȉ>�ɇ�؍��m�~����6pc9�����r�ϛ��$�p5@s�x��p�^K[��I�^qT�F:��!/ N�>Ja������$�YG_=H�����@nR�D���=�1�Lz��ޘ�oCålj�zpԒ�Y��x���ר��w�Q�{�^x�aP�	��$ׇdH�=�mI��{�jZ���Km_A�����8�����Q�|�ܺ����sb}�J���O�+>%���>�?������E��N�@ڹf���8�#t��������s���L���	��O�6��IU�hZ#G��'dE��cӅ�W�\����G3w�Ʉ�õ�)��~:���
�U��{�hA��IP�	�v3��%�3�|Zc�~��Aў�w��Π.���ǐGO�qa�B^���t욚��y"n��T�Z��c��� s�(�F1�#�W$�Ůq����м���[�;�tП���33���s�I̟��p���^0s�_ӯ�~@�$$��ҹ0Pg`0�~��#���z�[�v����Hi���=�Gy�NL�$f�u�U���s�?DV[�|o��?��v��¨*[�TB���(�\'#IEEyͼ*�%g0`=}����E�m�"Y-��be��?Eӎ��]cH��F�4<Ts_
���c�j)�P�탙^=�w!�',롟�� ���b��)G,T4`5P�+K�K��N�dD��}�nB1eѝ��bZlE��D����_���U�����P,��Nl��me���T�?�ݸ#&!�?GF�Y�s�u4��EL���׫(�|��bF�$Wؿ� ��щ�=-<��$���W�����5�!�m�/�M�v;�[@I[�ҧ�O�m��A*匼�3H��U��<�3!°{z>���L�B=��e���-�Z&� ��+8O���#²�v�ei�2M����^�h7��*�����Q��ö!�&�7��*�Bs�&�a>E|�EdGy8_�uTDM����w4��N���G�^+k^�������Oz��_Q�#I�˛���P�؀u�M������[ˈ�Ȗdƺ6�s��j��EC�̑�q7���^�Pq���ɂy� 5����P��=2�`\��x�oq
�^�p,�8$���E��O���^��f# ���د����Ũ���=r��P/eU'�u{�è�f�(�/�o*4�\�E�2AM��r�p��;z��Q���{�Wh�����w��&%0�ҡ�2~q6UU��\��n��{͟l�HP��i��M�\�F*��S9�(/���k֦��Fj�H=,T}ӲYHƉgU厄=�����ڙM����'���?\ɣ�3�/�`lN�.w�b�g8	�HJ��H/t�"b��SQ7|�y�Did4Ȅy��_l,I(�[�vu��)�O7������G���S'���t&
��=:ײ/Y&Q���;F?A��X�i���:� ��N�0W�n�>��3���8�$ʓ������;�h2�4&u����r�� ��_d�msk4�Hd�Ban��ˬ�~Z��y�4�SG��k��О=�#dƙA<�@��)�9�Cua
�YĲ���á$_1dc Q��x'��L����m�8`���zx r`�r0G6��;���*�6k"bq�f�!��G?��V	��<�pa�<��sp���y��C��͓��_����QwΩ��߾�xxD��[���~�OS���@x� �r����������n��f�232��wk���R�c�D�ƀy���o���I}��	�B�|�P{�,��X\[����_���i�-�`'7�
�QU?+�*��f'y�*�m�#	oB�8,����A�6r�8QZ���iS5-�Z@E�q�Uq�fk� 5�(V���u��������t} �3u�.��r���2�O����)��{k����Ж�ۡԪ�#�ᴷΏZ` F�VD<����R�ϋ��t�K��TN��מ:��Ңo��@��i<i89qW�EQ*�͆Mo{�3���ҥ���*��檣]��9��Z.Z�x_�	GOl�:'ݹ� �PѼ������q�BU����Ű�T�
&��tR�@�BY�h��,گ�BBl��Qa�
�T
�I��lY�C��TX� ��$sӠ�O���1��-
j�������Y�e�jۥ��X��r;I��Bz��gV��H�G������Қ��L��R�tgK5�6 M�K�pp��������y�� @1��k�~L�~����G���E�?kH�r���?6%`�y�60S#�?��y6o��<�u��Z�h%Ni34$UJ0Z�q^N�)V��"TȨd���&d��K6��i�5a��t���ŕ6��|+��Ol�/<�)��+��Uy�56{���,��Q5�����J#^��{(< Q�b�U{��+=�NuJŒ&�B��S4 q�wKPt�㾋Ȅu��7�O&?���п

���Z��`�t�/J�y5)Q�R[�F����%c���^�q�Z�6�z8X�gl>k_%��s�E�e����M,��tt���u�1��=�F��$�R���JD�<x���dF�6�։��q�����&q�zs0�qf+���R�+�%"�t!H%�vcȗT�.1�#@���b�^���~m/Tpی�5���z%�^�(հD1�`�&�C��$0K�������ҥĶ!����a��Ʈ|�<Y�F�9%sȭ�>�U�B�P<��-�d/��	�nc��`(���r۱���4/�&��ݾ��Xs������p��ISKiE-H��dN��hd���|Ocŗ�tݹ#~��F-�s^�W��>Z�5Ci�� 
c���]	�/�f���2!���x��� @�h�r�[�Z���kb�w���~=2Ը����A�k��3�M4F3<���ﮋ�������3:�K�d@�#	��ҙ�:49A�/ծ�$a�Z�=2	���$��������+����қE:�ɉzK��-��f�#��(������=��FM��gوxĕ�$�c?�6�N�k�v&5Ba1.'{#W�������	�>,C�F'�k�{�=X2Y3�bg��2#��H�-�ׯ!�"�#��e��=6���󖰢і�� ����kp�D�HW"��Z��N6���%�������h�&��T�r�E��)����Y�m��E9�/��� ����9��G�_ؕ��7u���<�9-��^�cU#�b�h��Fө�g���=���)��m랾p�F�K3�S�T��Q��45�t-��Kc������=>�8�c�����A��.� ���5<�u��\���HԁT�������i���_U9	hPS�ϖ����S:9&^0o�Q*�7yZ����l�U��e\�2�ȼ-�(��w���bs��9pB<�:����>��C�vBZ5`���� X�:�J���U�u�P�c8C�7
�A�(�R��~$B��ږ)��bPF_��]���t���%Y�����,h�{��7�[���g��~��x�hwl�NS�|q���<��O���Q#�����sf�^:7��g����(�Ǒ<vظ���X(;{�1ݰ�ĝ�_B7f	����@��&�}پ�'z
�E��i�ɶ�(?�n�"�u��;fB�k���
�<�EZ�Hg���Vc]X}��wxb�/�M��P��vMJ��WZצ�| N%�;��7�E�9��)�K�9"&Kޡ�<r&������I�z�T:ϖ������gU���{�J�9W�e%�kljD�a�s傝1��e�پ�=��6OoN��J�S`ݫ%^���7����x�ĀaA��B�4�[HR�#�n�Wj�JV�o�}=BY�4�a��> X�.���uRa�	�E1P�BaU���Fm���V�:�t,�Z]yӶ�./�i��ء�7��3�X����r�ƭ4���{ßkAp�%]5ѯ�C�+\)�v���"���&�5p��!�y�
�����vki�Co468���S�ƐȤ���P��6�}��&����l����&�YV��Ƣ�K!���"�]�g䖦�������cr�C�E[`:��ޓ"A�O��)��Г���P��f�+��g�&U�Z��5���=�hG$����C�yT��������ca<uAW��e�]Ɛ8@�(Ƣ����m�f]�I]C�1��mr+�m���Q��aK�@����j�Q��b$�w%hF1��1��s����hf�ճvG����s�S>$w�����?��PM��эX�-�6��
�w Vke��Y�r�k2W�ݦ%t*:�� �M�C�a^}G�Wqy�úCTY�얢>Ц�1�u;T~���x�,'mc�a	���P��٫����i@ϸ�Qj�hKYQ�P�V��}@@\y�� ^1 xu� 붒���.~Ⴧ�wf��bn�/�a+ֽ�v���dO��94r(�;H�@V��-�GO,X�U��o"�[�`�LP�p�a���`i����h��
3�Qʼ���������(͋��T;>ٌ���(6�Li��� �����H8C�UȊ)���Xa<X���܆iAZ`�JQ�fZ#:�8'Ch-� ��SAW: d҆j;�����P���	!�կ�M18�zZs��uqe�r^@4�Tз�� �>R�R��c�<��*@���{8�<Hw�L������
����������aq>A^��(�H�X���7ig_U���F�N�(��+
�#B��&u���~��k����"G��Z-Hw.���[�/Ж�G�Yt��h�!1�8Y�O��zo$�A�^�pm��Ͳ6Y��&J
�ǲXf)����?낽�;�����'7\���t��n�3/<�'"�[T:�M���e��C�2�����ζ�] ��5�ٰ���S��ʬ�I�Em�\�NYN@{��F��t�j�k�������4�S.֛������w��_ɧ�7iI8ezɑ�cY���D����X��0cSEXݕ��y�ޚ$r��Cʑ�{�1�1�(�"��*�#���2��W#Uio��k�PvkY�1s���AR��񴑕$�o�+��N(����e�0������8��[,qk�F�a��zՋ�$��;wq�~����]��M/T0��[\Ǥ��3�d��ؘ��Aw�?8ۋ�4mf���[�ߠ�DZퟄ��J�46Β��H�٣2Hd�`����0& ��c�Q��/�?�9s����G�Q�,�.����mg�% ����ڥ3���yjKs�Sw�?�b��?oJvR���'���~��)��b
�
2		���HP*�ـ\�<�L�׮3a�$��Qc?��D�%�%��&p�l��6����ޑ��FP#�Ғ�L����e��&��G8�L �rr*\�H�����l6����"�ųǇ�f�c��lO'�e�������[ޝ'�KZ@����M!�������Ѡa>�d*�HɣWe�;���b��G�	P'~���:�	���#��mCw2(�!e4ߩ��p��t�x�/$A��O���y����0)�EQ'���&�#d&2u��%���$<`���>r��Ɗ�E��qe�; o�)A��mx\=ʵ�C^��3��h�N�����:�|0��Z�3�' ^�U�<�"&�_�wb�NR|��SI."";)������aen�����U�ah�iQ�D���ګۚ��V�d�㷥�!�TU�t;�W\���@�_�H0nnfM8|�X푟(+�|���;����=w R\r;`�bVX�?c,���ƌɉ���*D0�.�RD��.�]u�dG��`�hT��6Y�`�72�ﴫ��U�i�:�����؞-�Tx�u���Rd����S�6M2"��;#@�{-���X}Cb�ngb�r��(z�����X[��s/E\�v�˶0�u�˹�
�JBD=�9P�/�)�5�����M�T���r��w���P$E���6i�,�lb�9�p���1(�(]�~����� 3@�J_�&�E��7���J��1"ۦ��)G^yn/�%L�����_������R�����Cn0�y��Ҏ/(��l6�4���㑞�O�<(ԗ��C��$��>"���V���#�⼧���r�f)�M��E�&�2��"��.��:"����!$&�w_�|��������;|J�������6�)�zڵ �}��'m�Ga��(O��{��l�Bi��i>���Y��^�BM�4V�ڢo�w�F!Q���"���͒�΃42ƛ����,��)�����CQ�Q�C�~ϐi����Fd�iQ
��3��Ę�gPȲ���΂�o�jEC�-F@�I�C�tu���;
E1�}B��m�-h٩�D�(��q=E����G���Jٍ���\!Ϻ��* �I���,#�-YL�3A���2k���W��s�������,��Po:���ݕ.�����T]��'z�@�l����I<[Bq@!�ح܅�RouK�?\�fQv2R�&��)�dY�65N��֨~�-��鹜f8�Z���.S�A@�.�j��gvK��߶ܗ"t��6�Ѕ
{y󣀓��X��qZΕ�z�\o� ��j;�%{��={z��恳��UMd�Z;V5�T�v�D3޲g�A��@#�j��6A+T�1������܍62��jC^!��#�_��S$y��� �<���)����ҡ��pt��L�2O8�.�����fa2�2��h9;\����z�"���)��|�L�5�SrYl6r�jæݫ�E�M�u��zS�e�� �e�d���^����YB�bz�AC��o�>��O��0���&��H���V@<v*����K���n�]�Em5���=�=	\*3����l�<pN��n��i`�ܘamȇ[8!�֯� BE'1ȅ~�����"��m^�;U���[�\��vCi��L���;w�h��"Hߔ���$ر`��A4���I09�P�{J��a�'���g<	 ԁ��Mi|� �NH&�n�1�����SDřIZ�;�;@3��V��/�$:��������T�m#��$� ��G`X�)v��.��虋�ϳ"eD�T*�v;�پ�i����F&�y��S����$I� �x{�uɾ��4WaNRKXĴ�̐J�u0Dn^��? J3�e��AY����'�'��i6���E�ɯ-̖1�b��Ki�?��@�3#��VMw)��$�	��'�c��b�]�~���Xh.-�4|���=����-�ف�Pf����D�-T�<��z�ZuP�~�"��� ����l86k�M�G����;�Iq�lƩR*q��a8;dw<�R�M7��g�ӻ'�_�'�:��Hwϊf�'#�`'��-�z�^q��(:��?}+0�z�M����� ��H���T�(K/�VV�w��>�D�p��㥁"N{#p�y!���S�^��(�^��c�ʉ��CD9�6N���
vG�v�|5V�����Ab�1��X���`4�N�:ӋK�]y7$/k^>�>�nh��f�pݺq{�\�.���8j��B��wT}T��hK�9z��urޒ)�����q����/��wCx:v�zs2g����X8�HIe�|&��RMV�Z���[�>�����,�S�U�p�sڮ���z�x��o���9Xc���>#Ō@i_�C�)��`��<`�h�Zz��|8��/%��*�ݴ����՜ʊ�m��J���(5"�NW��	~~o��g��Z
��5�+����^����u�"�@�$�v��$:�Ը��0�!�mmP�%l�Sv[Ue�a���Ζ&��/��نËb������()ȩ�E�~��@:S>��PQeqEe���t���Ɗ�r�5�6�P��?���1<�x/X�up#g��6"ut=,/{ƪ��� ���(�d��V��Nw�s�	`9�:��!��Yp�mt!��T��ԧ9ʦ��i���򮧍r� b��%a�`]�r4(_��.E���̠k�@(�jv#�8��N�L�y���Ry=T,��Q�y2�.{����8�k��B����0l7?=}��b��9\]&ə���c��T-�fXf�:��� ����,��;�0�?}K��+4�x�0a�J�v�{��rq���?b��)��\�����	Ƥ������	��=S��R�2W7�>�#]��Xk�϶��>)��JjCS�v��k������A���!t�Ë�F���#���)̞���XZt��j���u�y�=���������1,R�i�~�W���̥C1�Ո����}Fb�fdm�'�o���+�8mx%,�)�`��f��[O�L�wz�E1œ_iM��u�?���7�l���D��t��t��[�龪���飻E��~��b��꪿�N�eig[�+Ѓ���"�Ks����*l�|D��g�N#bC���l3�Z� �^i��2�cVP;A����)m.�bb-��>����-J��ݝ�N�b2�3���P>lҍR�^�ּ�Չ�y��L4������1�Rc��#���,ԵwKs�SH��[v�W�A��_"���3����0��+6�`��U�0iX"5�&S+uW�F�^�o?�lGTc�������!�����`�-E��<2+��S�k�Z@���P=�V�IVɅ1"�.�CɎ��ˊ0����No��C��#u�1�>���0�����Ў�l��횆_(ֈMf�%=~���p��uv��g\-��;��솬�zr�e,�֞b��dA�l��\{,�'�D63C�G:4�)a-'�N���/�6��pU@H|{���{��徐J:5s���E,�d�|K/M���R�g�WJG�7kQH}��wh=g��4�Sp�(w%�-Y���"��1:tZ�P%��M�� @�����.���[z���6Ru�(�z3�I�&���sml}�������6)�� �~���j���B�R�R��!�yX@0뭱U#�Z��+���&7���O
3��7�ױ[��o}�g��_�uQ�9���/�P�C��Ju����0y �pu���s�o��tA-� 8�t��o���[(�^�	��ވ_e���I��i�6%C�oجY��`�!���zBD���	�7s��аV�k�w�Y�(P��5�/&ѥ_FNm�� d�m�/U}���<N� ����Y�F�*�J��)�Y�~b�W�#gl����Z�q_�B�z�'AD��x�2s�?�:�;��Q4e(���H��Q�9�Ha��	h�8ъ�����_(^��?�O��Ytc'e�l���v�~�űӺ��9]���Qw�S�95�/p�<ӵ׹Z�u��J5}�v�I哅��jb92:�Ӟ�x��g��;7[�U������+��˓�FJgZ�XF�����TC��^��I\c�~Vt�Dp�C��"	V�:4��<�i�,L�~�l��+q#����ַ\��ɟ]���S��� ���c�I�@��Ų�� �w�-�b[̇�	�qXs(�fo��	"�a�' a��zY�v�`���H�P�7��G�J!A�XG���w��"�1K�`F���#��&4�2��-#m�����A���-�F�17������3ڞ5�E��xl���d&DS�r�9i즠����_MX�ZŸ�� [�W�i�+Ӆ�gKj�U�1�J������7*��
C7=)]��j��^|��ZE������"�"�*�F��s�E=Pk�l�L�d��~I��s��0�T�=�8���i��{���k�q+���F�*��� WU�- a���@8��O��Pѫ��u�#ypĲy��X�pW.%P_7_�_��S��N��u�?\�g��0'w�hw�P<W���Z�
z01�����Ɖ���=���w���t����X���Cb�+�)�,��^G��l-߀��;pq�p��̉*"��ΠQ�����<�h#�Z��B&�:������H´�%?���	FE�9sf�,؈A5�rJ��8h�dݯh��M��0�f�o<8K2��=��D٦�P�O;���P�藊�p���4��|�^� ��C{��U~��@���:-����
5�_va��p��∬�^�*h&,��A���Ĕ��h�����{����)�,�=�O���=�Q	�:Ç0d�%0�F߱'�ĸ�N7�{�CwQ(rt�=J+�UjDW�R�8��wu�`tW������*�S�Ob��.5a���kMP��w{>.~����A��%{����.�E!�9��F�Eop��+S1r(K��+}��1n�Z�>�D�{�����T�L�.��v��p䗨�2�+���	�VMk�#�L_0I��ٌo�$�Qխ��Ul?�� 	Y��L��Y_���d�]/0� �Bx5�*�h0�6K&���}V��T�G��2��|�Ե��=6U�Dx`��n�Zҕ��'�b�E�FC$ħ�3:N̕����lcߠI�ė�?2��[M�#�@�i�'{[�`�����$BYw$x!Mڤg�g����!�f���d�T��;�$�D�S=S_M��{j0#��L�E$����{������6a^|k$��� �[|נy�1�ّ��?���j�ۈ�qZ����gǙo�5)5wd��n+6���/BE�B,�sk��H4
�e{��|t8I�B�ۚB�.&Y���a�"կ$Tړ�@�3��r%�'�(�a%%4���#S&���|v{���b�XO������sJr(K
2,�����������M���/��Ǫ�č�-�L4r��5x�j�Jc��IO�{f�^���)'���O��-��>�X�r�I`=�v�˗��4��i����V��06*ET�3�(����Q�u l,O�(v5o=wIY`OA
��bSF���5�T���m�c�t����c�&�tSv�r�4���V%��d��}O���Q�`��?�t���:x�.�;��Eu���4��k�f>O��	�ٶ5o<�L ܖ�8j�s]�O"4��,m7�x���-�<e��!�V��,W0ߛ.B.����\�����v_�""��K�,#�	Κ;�G܋C'��FNz;����r��ygn/���!wdS^�i'Y䢶�KO�"��HG��u�z�:V�?n�f�r���<����@�e|_��#L�S(.�vO�Ė2}y�]c��nfo)7,NЛ�3�wb�@P���D|N�;�ԇ-4JlGz�C;͂�����A]�d�j��RGdG��Č,$�.�2�w�(�(N�\�/�iߙ�I}��me��&a�U.��S�]T����:���F�����4Y�k�BmG0�ö%)���9uo�7�OZ�)6���F�#|L���:�+ j���z���"�DU�~kYYn�|*��|��L��A�E&晹��^�эI�o,V%r.��T`%�z�ڐ5��&B�k�� =�d(����=5�odNk	@ƞ���t��	Q`0'��B�q�����;vǓ�����G��,�k\R
=()�I�T�5��~1�KG���((�l�=���X�M{0U���N�^���fè�~�����,�]���W܃3�&�Y�_+��o� ����:��OD��Ma"���(LS�|�[�rvqu���P�VOEnB�VV^��c�=s���3�Ƥ���c�A� קW��X6�6]����C�(�f}�g�j� 7�� ��<RM�zε%���\P�������/r,������;�bs�P9���8-�gOIt�!��o�ƨ���
@�2Z�!g�_����|{ќ���?�V������$�ʷS����fE��3<�S�Ҟ��c�W[�U���}}G�ؿ�V�?G���0x�����n3��C`hq���H�y�@�[�J�]�?�*JVJo��D��w 8����3�!���1�ȭQ�g2n�)E����5� ����N9���O+�oE��S�8��5��<:�����>E�g��GDM�[��_^^z��{d�sѵ�6�IN8
~����Ѫ���\8��߆����J �v��,Aڤ%5�cĿ���;��
��+�k�P3����ughP3�/�G�g`N������B##���e16n����=��������Q�ޫh�F��O��>�]�m_/�^m��7*
]:�JRn�����{��;7���u���AHWu��xT�$�erL��2݄C�^��ۢ���-zt����׬U�t���TB�v�p�k�����%K�0�_��NL��,��1a�8�m���~��/���.�È��C��V�8�5�рus$��D��j���T�ld����?,c�8�s�V�5Yϵ�)�M��MiW^�]q��t~���՞� .����4�>o�.Oc6w�XŹ�CLP����1���p���pџ�F�hU84�b�@��6Jhn��F�(�s�C�2ܜ^zL&�ߤ����M璦0�`��[��� p���P��I)Q�."۱M��j	�����4Bmj�O�%D�k^E�۶�K�P��YPd/2��/�3���=nӦ"�>L3?m� h�f������:O��[%s��:��SC�U���g����4$\'�#R��n78��9Qу���je8�������A
�'T%99~�s�U���N��B���0˴@��>� +��Z�_��G;k����|�*�Q��� ����Ȯ���2�X�>�gx�T��:(�l�V��2K�e�9{J��bK�+Ȫ�:�@£�S߲�`!�CLu�N��AV�A!�Z���I.nN$��mk��n�������X��6i��̓FfЗ�_�,\��M����D�*u OA��{n�#�t����B�w{.�S*gO�P�����P����zT�+~�6<�m!��\jv��i���N0cm�4�������C�ܶo�֠���o�l�C�� ��~����pT����$TM��Ky&�e	���2�fly�0W03G���0N�m0-k�����z^�t��Ms�)�<d��m�4z��%�sp���]-���f�  ����T]�KB֊ٶm$���*�,�E��!�E�(k�7�1b�7�	�4D�O�X�^�i	mG��@^���20��l���4���wc���h'�������{g��rF?��p�4�7�1�A���S�^}g���TӋ��t~�ų��-��^̳%�؉��4Q�A���uqz;��c���l��Е�װa?^��^$sZE��I���&e᯵�N��6�y4\�C|�H:e]�/Mt��i#S�%&�A���uF9x��PE�&Ρ���^��@�j�"'�]���7�w�1�������9	�u2Ol������3BT�]�`��/�`Ӵv��㬲$
]�� O*�w5*i�A��]痘P(��v������8����-�0�:��lG��G��Qw ��Q��t�٢AӍz*_�\�\�|T�Ec����ofͶ k�%Y9ߡ�Q&i�x�O��
��Ss+U-�
$�_��S�G�߇.yH3�$��6�lˎ���S����պLI�[LT^OmR�W���C�36�fl�r��u���O��\��0�� 7�:�<w?���qC��s�Gk��xJB�����}ʾIG�[��<�}/Z٭Td��Bmp�_�h�Ǻ�T�
3rA(J_��_�+�3o�`Ҳ�}-Jr}�G�Mw�Y�I�Hu�p�)�*j��O��ٮW��GT�Ye`Y-f9&�4����O>~�C��*қ?��0G~�M�E���>r��t� �~4f��Q9�3I�N�>�dAB���D\�hRa����|�h��R�:V�љ���@��J�K����#@���H�\5w����}h����>tV�ɸL>�?M]��X6Rs��[����-�ϖR����7�;K���B����+�I�s�(��&�ؾ�ѭʍ�;-�֨�O��'�<3�o�t�hE���pC����Cf�8�rio~gn6�}N�F�H��\�c3�{�7�<�|Ά�E�'�l����ix ��AZ4��ҁM��&#�/g��|�۸�p4����k)1�+�#�xh-]j{?��������/(�ܞy��m��
��#�����"��=���P�\���Wc;bE?daS�����i��e	Qv
G���R��~P=�1�7�����,�PbP�xTF���TP��&�4���
�	�@11[�~v�D�x�B�ۚ��m��)�G��$�6Y��j�͓V�i�pT�oi�s�W��Bå��)l
Lʬ�'�3�K�]�}��M���0L���Fdu\[�X��*�������j�rl���J��G.o�3��.�L����GS�(�eA�"tGq�+��Nxz3��%匿Pph�V�ꗽg��[���8�P��f�8��#�WB�/D�m�8��G9�|s7�^X�[N��|nuG�A�Bɀ"���9�?�Z?>��HL�_'Mbr��t��p�U�R|b� �-��QM�Itq�����ͅM�u�%XB�g2�2�����r)EUs���L�E������IL���^z_���xɀX�}��T��V�Sb���7C���Y�$�X�p���
}���okvv�����T )_ú���r���*!Lx*F���}�ފ����FP�<�Inь�FO;�Je�>�3[ez�4p��)y�r\~���3���\�� |�/�"���D���z58��TƘC�<�p�)��-�]�~��R�./�՟��U�^���zY8OY�dN� �D�S9��֥���4p�߲���#�ʴ��N�0��޽H��{�l���3�=���j��I��H�l��x$p�D�N���PS�>+�4�6�Q���
P?�>2����do?�&q��7w_0���B�!Rn؎H����\����8l��@Ed�s2���ZE�x��#]�O�������Fg޲պ&e��� �va�W����; 8�����P��Z;�pH�?6�b�,Ԗ�g��6��%� h��r�l� �8��(èע�I�E|o�h�`D �R��]tz��u���\��j�N��辖I�7�4i��⬈ �0�Oa o �0��������4p�t��B ��Jt;��e�*�$�R�j�m�>����I�`����f�w�N���o���΢�0_T��u�궲�Y��g�NZm��=�\VB�]ȤVeʀ��,�v����]�춐��#�־\J�h�﷼D�Un��v� ��Q;OF{���2Cc�r#��Oᯟ�M���[j�2��� �M<�3����L�x9	�^*��F��aBO�3�V�Q0㌅"�.�IX�#��$
}��VepA��?OGgw��B0��kK��	����Z��a68�4^u�d���dO��"K �4��UM�����4��I&�U�p�c��D�y���
7�4���;Ʉ^y��_	�/O\��8lsa�&�ը���ǎ�޿�NxV�J��<�5����Δ�ӗK�V�R���@9�ar�!W�ģ֐��"E?Q >cg�jG��)"9��I<�iXDJ��Z�+`5_�,4<�	�~|W�`X���9��CZ�,U>���Y�x�	I��k黊���Ի���כ�y��'l��g�_y�Vk��%��-G�x
Z�����y��:D<� N��lp�
8�B��1��&���ӎ7�A���9TF�,7��?���H�7q/d.��[����X>b��P`��'���4���1���~uc��	P��Pҧ1�"#��˱��>��|[v4��=��=�>�b=<bS~�I-���ǝ�����S�z�>	5g"�o;3�v����c�V?�(���4E�C)�B��2z��,���E�>���=�*l�^��/���j�����Dv��{��Ԛ������K����/�ba#��&�?�L���;i�HO�(o Z�S�۫���Z~tUY���3l��91�B{ȍKh�nqju���P0Z�$֥#�����
�i�����_z���S�����V�뒕f!P�%I��È�g�tD�>txn)�@�`�)�HE�P����).�C�k���������#��+/���_iTK���Z��˦�J���щ0ӆ��c�Dd�U�+d'��J�7��J���쫹_qv��b Y��|[�݊����]ݧ���A9��g�)�+i��q��쵀��GѺr
	��+� v�H:H���j=��5sݫ;���$��W�Lq��C���>����P�y�{oF���F�j8�:!N&����Y6�2�"�� ~������*�J?�tBm�|-_|�@�i�$E�2��%�j�u[��5o��X�x_�okl�}����-��t(�iT�F)@*�-�����/ �`~E���1�<��N�60�ٸ��+ܢ&���x����rL�1#d�:�D�uԍ+ �fz�x��tR�þ=�j!���N��МH�&�&N&�i3��XKwDWU]E���LHU1�A�Hx��7IT���[��W;���ts!T*�z�;��C�EX�05 �(k��m�:3�ު�m}b�v���/�D�̊%R��@�pA����_�pөQ���|ch}P��@����S����ڵ*y���4&��ax\q����코!t\,Ӛg��w$P)Q�$C�6�a1?�3YA��W�������*�Ģ����m}���?�:d]M��љȗ��@�ɷ���#��;@�����0|���a}GnR�yl��<�}�a�!p�+��k`�@{N_��Ҥ7���<�>2��R��n��J�<��Kt�h/�2�1�#k�l�[74���Nz��
�b���Z��7���X��WPkA%4���2�_���$[���O�	����G���iU-M����K�]i�4Q����gn̚y�s�s���&n*��QdCk\݌o�N��.��=.�</ �����F�2��7��{%�v�o$ĭ�W���y��Y�qY8��J�lm�zQf�M蠔�j��D��p;��v]p��@�Ĩ����[Y+���O��1q����'R��Tf	�w#��81��ʶ[m����Y�~���xT��I>����̠z"���R���xO����5��|(��3�'��.��ma��J��o�$��)�c�/5n�t\[���t�m(�T�sE�0�ٔV*���ǌ\�ؑ�GZ]��3B�@&���KG|��c����}���
�rh1��$�R��URoq키�X����F!�
�v��긝C�ܴ]��']���r,�wDR:u���$�B-�E����F�$����:<�ش��J �S��d�?���**��Q�kî+yL�n�m���P�EX ��F`s�\�I�e��Ċ�����9���>�&LkkӊǨb�3(֤�7 �g�vS����<^ZP�:?��G]n�p���uK]�+����y�f�̼���ev %�=��(i�(�*��S�e���,�s<c�)pxM�*�ȿ�9���O�&y<�|��1��mռ�J,���\E�q(�1SFn�9�,j�c�=� ��%䥌_�f'����xa��$h�7���ia�A���nA�?N%t|�ņM�wg��(ʈ�ڮ_�U��M����n�{U�
b��1R3L��Өȶ�ޝ�f�y]C��)��ms�{��O��J�n���������(�~�t��:�q�j|VٌA��If�A:�<�����͙ܠ+�M���6�S_'%7hX�1
C���M�����0f8���Ҫ�D�L���Ҹu�[Qv��Й�B�G�ɧF�|yX��x�];x����;jF�I=�krU;�a��*�b�X��z$���B�BK�5�3�*�Bs�@����]k����b�����fSh�[�̡ P��F��f?Q��� �(�	2	�f�:�
2�D�V��}��=��KAg�:�(��=;�4���Z`_V�a���J��,�G�q�T�~p.s���?!>8�߻�r) he�ڮ���)��p�˰o���ƨ	0Ԝ��@n?���m���|��Q�~�Gg�f�Q��X�л�Л%Bv�"�X� ^6�H/��'\O>�K%�G�0Cs��MBs�����W�ɀw�3�D3z���㓔tf��|�@�a�$k2fN��4I�i��0���p����s�9��u���H�ug�CWf�m��W9+u]�~����{1�mx��i���Z6#���g���j-T�`�@�|�S�/�e�'��|o���L6���ԏǯ6�ӞN�'����)�ƨ#ĝF�_6�T/�T�B�?Z���\r �b�HƂ��Ij���-gi�_z��+(p��Eo��U7%�e�1�]q=@��?A��B����@���R�C*�$�j��P���_�Qc��"&�6�:{��s��ym�D�7��ZB� G�4,Ò9�`őe&�tt�C⻫�e�G�����:Y���I�3�a��i���O��5�t���N�PV/��$3����mٿ��HCb2��i��͸h|rWꝸ�e]n��T����F<����"��ʀ½$}ڀ��Xp���XOkRdm�]BX��垁(�r�t���hC�㔁RN���~��>K��fC�e�ټ]���q"���m����e�ybL�u�����N��T�:u��K�m�:��Q��A_�ގ��թ��/"WilbVU��*=�\5z	�=�3F��ly��h«���3͒��@$�p��׭�,��=�H�8��q��c��X"��2��S\�(�Os���7I�,w�blV*�8�I�+N�o��L�Q�����mΕ�ׁϵwr��B�f���>��H=��;��0��X�FF�pr�m��n�-B��;ϝ�]��h�-�ONQ8ȵx��cD��7�誆�_OB{R�)f� ��f-�%�n�u����z؉�~a��,�|߹�KʃCGB�`�����A���_�ڲj����Z�B��́�;Ԗ�A�K������2�Y��Oq��M*�BR�;�ɼ+�<	��[�b��Ջ��*���B���ڥ���ɰ(n�O��O��d��I���5[뷁8����s��7���a��e�K=
��<�B����J*�-�ے�DF����jg��Lh�ܟA)CflN3��I;+�=����t��|��}��3 Ӄ{�p�w���l�),ӫW��&6]�����yV���Hf�GTx�a=6�9��vE�7��߈��%eL��'�~f N c��yp�$?�~��l��2�t#���R��C��BR�l�cr��H�^9�IM���|��S X���E��4�I�|2~���g9^޿@�n\��-�ť8�j�mW��%fA2C*^��x4�UrF�>���}#��G���%LZ��c]�Mz{ׯ�����\�ܝ�(ڇ�[��{Wt��ꏥ�mv�[�	]et����}�t�j��K�&�7F����@�S����uq�[��b:���F���:J,���>T�Q���V�x�g݈��m�^":����]V�5P��i�2?W�G�X�cŭ�"��Jc��S߷�o���%�1sY��� Sb!��Jb��e�n?����xڞ���e#�K ��z3�&b�I�"���si#[O�z�7��q�F�p��mjC�DpJhbK���vp%{�� ݐ����V�F�
�ʐs�x����b�zi�NC��Y~�S�����b�,{O����h��4(<���}�M��R:��<� ���6V��#����2�~��/[H0g��=d�|O��̅�m��2�ׯt"�����[���b�%/��K&�K�i-����Ѽ�n��FON���@*�OZ�Ӛ�JS- �6��z����]t�x��Q����}��6´����A�n<j�H����K��o�,Pp��7��<�Y�X۷�eM�f 1���W�9�2��ٷCd3W�@���3&N*IV�]'�Q��S3�)�|s���TTc���O��m�k}��`����>�Ib0�k�3{�*��i�� �Y�(UU�֩�iY�[3��SNYݷ݌���ov��ZK�ߦN9�2 ������7�u9�^�Hh�B��B��W�<cQ���p�} �,�q���C��]��,^�c��pd84����V��iM�p�E����sL����)�/��p�r�fv�����5x�E:�;��eF;OV�t����ZWI$�raLҲVr����4[^���������ȴ��{�bw������6��w�sV�g�E=����8�=�P��y���6%7ΰK�hCՇ-f�6~7�['�<4�^NN5���_�@��w<�%��{l|���0n�>A���aؓ�à�5���\7'�&F��.�%�f>T��ܘ�0I,Bc�_�~�xC���opSɁ��L����i8˲�\��+X�ΐpP��58��\�h����X;�v�A<.����(ۜ��K^��C�9Q��6kD�CH.��g?�������U�$x����p'=��"f1��Ǒ��ΰ�wH9��U�@���"�9�$����>˔�f_��g�!�yCR,~U^F���Q\�b�����3��!��ۇF�c��m�o*贷ڡ;�Y`�P�^P�j|S���],�r��1��� z'���t'55΅�&�2�� EZ��ۯ�u���n�S�-�(]�R�]:{Yz"�����X�l?�Xzw��^L������A1��}�'e�^ځ�������*��8��P��%x��V=4�ӥn�}�c.�_��\��G^��j���vV�8Vz�SDo���q���N��>2�'��Bw�"�Q�� ـ�Hv{^艄�w!���m
�:Ȍ)�V��� $�A!�#�ϳ@�>���-�5��T������5�=�C�ir�J"\��2�w`�d�y	��#�C��98��A�gP�T�7�{��Y��;�şEj�c�t�<${fa�f���(+(&�Xs {�N3>b �|�\��\�X����O#�IPp��wdi�0	������7z���#8�f�F���Y3;b�!m�=W��(M$V57�R�Ȧ�VZ�$�A��8��6�KZO�&(|�D74N@��ih�"��,E�6�_��a�<��i'�qDo��k��C���C�5b]����rXl_yzEE� G�D-�إ��E\���uy�4Tw�d���8�e��_;�F�c�
	/R� �J��3�d�e�?`Z>� m�go�$�����������r��VQ�]И <.+a�i<I���͐��v�*�h��)��7�"�^@���QY��3���ptޗs�������|�;���M@FÀfX�q��Y>�;���ڬ5����@��2���!g ��!b������1��kso���������H�5�aG��M�ud$1�A���A'b�Ff���5Xz*��G�Z!�C�ܾ�-�������ZBzsJ_]u�I	e�8C�h�M��0~#�k�S8�EX�\��I:�b�DW�'��u(e����k��0��������f���1���N@�ʣ����a_�|�$���/h�C��4;�hh6�,�Z����T��^X,��|U'�az'�C;?t�b��h�3��&���a(G��>a�6�2�Mv�'S�uR�Riׇ&"Q󺒶j-�d�n���I�������)EG����m]��6����կ�@�?�`���əBݡ��-b;� �x��Nc��+H2���h��x��E����τ�E.�DH��J��ɵ�sQ�&���~���x��د���1AɈ4���C����Gv�� �`�H@�JQ-�a�.2�x�ø��+�n�z<�Mv�׷��߰�V��0w<#���e�'fbF�,��@D���Z.,�%Ec�,
~5m줳�Ш�ZW�b)Ȟ�2���R;^����0���"[AB�:H3&U����A�9甠h�g{f�x�+���(+B-����'D�{���$fQ\sZǁoJL�9^s�U#dm(�̀vQIC�@y;��K�~���������e�7��5R�"�
L����Y���YD|�x~�x��U��V�U92�~��|%�G��'?A�/�&��oO�^YSe lGjAɏ�IBIhQ.J1��y�c��¿8�_J��gI����J�8��e*��x��NKvAa�݇�2v�ʲ����d����*�=�m���^|ލ�1ϾN�{?@0O�=C�C�r�ቫu��r ��EG����l�%�&��ޣ��1�E{͐�y�l���ӛj���d�>L�ۯ�H��E��l�����melyIY]b4��=I{X��Oɠ��E��T4�#5i��y�-
	��EK�/^�n��f��j>�S9�Ng�"!ݺ�\8D���J[�4�^��c��reWA�!��L��<BU�<�w���v�_���ɰ��cRr�A�!5zH0:��B�V�����Beş�\=F�3/�Zv ��A`6�V2T�VQ0Kz���JAvH��a���KW>��6j�.��׫_#�ϸ��Ͱd��(�GU���;ߛb�AR��o^�[�/d/�箰 ��_6��A���*���C7�$��~�~�r��-���i�-�V3�L[��U�4e ��W�6�?�v��Mh��sP�㴈�' �UskUڢ����f�x�[��O�h���,�q�HoT�I���%�X����V������T�.�T�4���It��'�����a�cy�"�8=����ķj�@�/��))�D:�E� M���_��$E� ̠��0ͬĴ�[ݼ�*�~>�f���v4���[h	�P���Z��.������|GsNv�<� �uR3��*��2�����6/P��57��ea��Ҽ�=k��3�����7+ )XVL	�7ȫ�}����op�A����#�_A'z���T#��jL
E���;/�PGe�K<�0p��<�[�������!�?n�}T�����?���6����Ճ��GU��w�������<l)�L�K$���V�bX�Qp��� ��k5�����bi�@z���ÂQvh�o�,�-z	*'R��B����u�'B��3����)=�sA��Yn�ls�(b��]����� �)�Փ	=x�9N	g����ǚ *��z�Ux��LM��n�
����
u��)b'�є|�1&�g�G�[�B�~I����Le斫-�q�}!�8ͨ%��8r�%�s� ��7��"�^�f���}�l��Y�$�J��)X �z���!��TT�����^�`-Dd	H�{F��	�7g�n��_LT��C�;#���X���I�U˱�#�l~`����mIj��=�?О��Ja�\���Uΐ�Z���ϖ���ȹg=���z�O�ir�GCYџY��V�1U���t�o��`��8&�|�`V�I�s�S(��Lj�pp� R����T��:�@kd�W�-gX?����ɭʕZ�	��7	d 82�!^��~A�%�mN'_��@C\��p��uI��<�J<o��B�)�#�F�	(Q5¨kfZ�/�精@��F��`�搾H �]t�1�6��Fx؍1	I���ډ��yzBn��DY�=�N=�%��&u䃂�wu�/k@�ğ���Ǆå��|��=���P�u����e5��~����c������;i�l@��dK�툮��x����A�c�
<�)���ե�,���E���K�d�p
�߱ ]՘��>�qo�#w#����p����&\�/�8�����k���m[E�C��i�SCݚn�ؙ�o���H[�`�ŷ��>P�I��M`�,s��o���~t�x��0Dn�I8�i��u�w�d /��LG�.>(�n�C5&���oh� V`�I�4�1���{���ӤQ���靂]f/P�-���"M�>H���qҗ��v<'����kֈ&i��~���Bi˓��������H��N��M$�g�F�i�B<��8)�2W��\`���q��ϵs�"�J��q/��\��%��@�3γ�f�3�v,���됬�AQ��~P���H��Υ�-���^_�*UH�=�?�dK�$�n?����0�RS����P���f8���=�e�8�
���3��&ĊK�~�
D�+M"K� ��/��|q�f���V�_�Le���h�g#%���L��[���of��EWQ�l�C2v7�ž��C0T���j��W���,
0#��� ]˵I�X�#�uՖ&����v�ݏ�d�_m�h��M��p0��634_
���7[�Yh� ����I�y�<�ʘ(��0n�䂪bd�S�15+�T����R��	|w�E�Nȿ��R�����Cs������+w��Y��~+������_1=��Ћ���|4��ꄅ�
�)VQM߾�j��t	U�%�p�������El�{Gc*C��@���j�j����S�F�'bڢ�9'Nݫ��S��0s�k+��+ob��}���)�lP���u"K/�7���{`(���U��u�o`?���ێ�� �6$$*��������$=��'���\�s��\�ѵb��4��[AM��U���e��n������s�n���KE��N�s�Q�,�FV�j�	$Y	�eT�Q���q�v#���;�?��7tw�ih^�3^a?���[\Z�ј|�b�'2�}믝Y��2.R�b�yה(�W4�˲��i1� ����8���0lu�q=b�<��f:�f��'��&���0�����&������j�"j��������2"�<:67�0��ttL�ٯ�/��Nie��e7��t�U^�i��g��]��%�; N-4#"@��J��8V�HbU��'"	R!=�=��F�	.�/�g�+J�x4�9���c*S���|b���F���×z�g�¹���n�+��׬�ưI��1��ڇ�am�d�!O� ��*���봬RU��3������'�-X� �N'W���.y�����ԁ�k'���nWFb�����6_U�y��B�(�4�J���mrjӄ.�ھ�׸���#A��L��*��*�kF�Ċ��m8�Uaɦ�EE��ވ����H9�A�A�f�H_8�ﻩa��-,��{Xx�,��fQ��#��ƥ�Ti + �GԾ���op��+��3���|�� �kH���ı��5�Ԅm8T	mʡ�!�@�|f���O�e���ڒ�fs$��#��| `%�z3�e��F�����(>�����	���BwRs����I��x0�pM�7,���۟Z��<�1��9�P�������]35k�j��7�e,,	�o�rv����.�3G"=G]2���4��0������U�FعSȲ�~���(��r���=�^�0����m-�l���0#�iǺ����	FCa�����"o�cǨ�_��G.e�N��L�/��"mFNT�k��}��iNn�H��S\1��3͸h��AkahP�5��Qx����-����G���x��
��R}S��p�֛�5{����كsMH�T���C� �"�T >��x*���k�ǫA��a�{Sl�f$�SgdÑW6�EA33�(�c���D/���@q:�{�0�1�c����5�`�\�!Z~ ny@�+!>�U2���j{yf*|n��S�z�GB�%��W�`�G�L��`�HJ�ѥ���d�p���� �4�#.%bSf��W[Կ�N��A��9�J��fUl�nL&��Fz�D( �Q�����ۈ!�X�a���R���*�p�J/����|p�/�ȹ,vD�!����nv7<�WV*��q2�H~ɋ��I���7�����e<��`"���q�n��|�8��@�*��b�Q1v�dǔ*��&��5�.�WZ���5�Ʉ@ߡ|���K�����g���'��/���hS~aN���������}�
�����h�+��H�
j5��{�r���q)[�3�xc�q�!�j���ŕ��� @|�4Bq�F��Kt��'�*h����@����>�e�a@ֈe��^V��%D�B��!$�䕗;�U��E'U�@���� ���%���?(KF�?߭
�g�ҧ;�[�+�[J�Z���h���/SJ��I��1���0�3�+w���W���ͬ�x�I�۞�A0�v(}��=ZOE<����X!2M9���k�%��m��C��O�� �������a���!�ZL�m�%
����X���H�TZ���A�B�Q�(�v�tJ��9�刯�x�w�Q�v�r��?�	�0�͂���Vޗ[G[?���2� o���E�
������nAЇ��q�앎�;��f���B�VT.v������6]�a��ຩE۷���?�*$��4���7~Z��Y&�ʅ��n��AC����P���p_dx����f�w��^�H��7"9Rڥ��|�B�'��C#�M��h�tț�>�@�������:��x�����ƨUw�Ū�k?�fΑLI��y�
`y"�����	��&>���n>���խ�J�y�ׇ�D���J���=�L��9�.j�uJ���Z1Brc���?<鼞���S*�(9�hO�,���Hm�����ȕOQ~����1�(��`[D���@��,�O z�}�M�|:i$�h��.�XP)Aw�a4b��F��?L�}��.��_���\^2�k�a�I�����r��ѧ��G�_��?���f4�h�%+���Mͱ|'?\"�>�@a�r=a뉴΀û�8�JtOcx�Oȁ!Eu
����WM��ш�-��Ro����b5��ƣ�D%��f8}sW1� ���ObZ����7�ho\���B�G����5ߢĮȒ9
ok
�e{8��,\Δ8�� ����)#7�dA���1�L]���۪�K�ݣ��"��P��P�ڛ���ly���o�v����&_����D��UӤ�CUz�����^�����k��	���9��g����<��`r�N �^i�H��
}�&Fh!��g�w��g��M����W�%?�e񥢱����(~}���z&���}W�Hm�nS7S�^k�S�XL@�K@�L�iTF��5�z��o�QƦs*y[t��D�
�m�J�Iļ�U��a��Y�����+2�b��3ga�� �>U>S����_/�Pa�SJ�R"'���,��[$���xL�d�o'}D�� +�I�r�C}3&��T�G	�2��T��g$@��k�h��[�ww�
���b���8�a�
��VO͎JT�>�>�&G�bR1 �2�*Q@3��#`N�	�V��f	�o��Y 
7,��1��5ݠu���G�S�:��^u@�ʁ�V�m%�������V�#��W(����h�a�ϸ=�ď��I;�aW����o���e̗C�H���5�iB�Pn'������ ���{�"��d)�t�â��w݁ñ@V���S��ͳQMq�}6䆣�:O�����9�.��H%G�b���=�O:'��47��h=Rěi����+2�a������������t�`h*���b;�\v�"�`F{#ɦ�])�?8��x���9������p�,]�������tD{����%(KCQ��=��Ƨ�b6tA��^6��%�@s�4�y��4�_(1�*�[S�TA��Ϧ	<�~Ȳ�?��Wyru�̈́a����eg,�v ���U�m�N��K=�7ˉ0�7��sX\K��N;�ۓ����,�:�n�.#-7�>t[�<���l��t�G\0>Y70O	 nS�*P{��F[p�����W<��e�ࢶ�!�[�!޴7�H����V݋��(-�c<�"��۫��,mٲ[	SX�u�_T��nFkm*�����B-��H�O0vP�F����p�Q��K��~㘧2FOR�_������_C�]�:�W&�̍�-PTyγ\�=�v����\iٯ�����:��>es���97�^�e���Uj�U�����W�f|�B��+a
�R���<*h ���ة�'z�� ^3�h�u��F4����,��ಞQǖ'��.	���B	�b��ce���ew®���x�[[d����\iP�.��9نR�q��Zm���OgH^�<M#R�Q�S��B	�J��i��6I�o���A's�<��?~P����]�z���A��OY$弐=�X��H��H2���4R��',��he�Ә)��/�Q|�-w4��I.������	�'9@I�(��ƞ�oі�Q��+ݟ�uv�t�n�a/��-yF�)��5n{�GЫC#%�i�te����S`4��9�V�������C9;e�yiT^��X��nkQ���k��/����g;�9sp ��զ�h�]�~�@�c��ҍ��C$��MW�Ɏ�4r�G�첟�
\�+^���Rr�H�_�,';f�
99�g��q�"�3NYK������xؖ:�d;?�JTOo3F_�i��(�l%2���Ytґx���H��vT�A�����"��+�1|#���ڷ?�yǩ�����XQ��4�V��9n��p�-� ϝtv�*$����(��7��%�YH!Ʋ�b��:���� �lHđ�?��������0��	�����e��h78 H�г&*o���_��LcJ��ef�T�b͝ ���#.���*� *n%Z��.�N�wZ�$�+��adj�e�^�D1y��F�L|��ĩ�>�$f��Җ^�_|�H�Lߔ�T����9<�t:�>gb�����[���`�9K��:��m(��F��|@�����mҝ�E� ,~NK�~f�$�ᳮ,��g3��#�i�J1O�l1����xA��f�䨞_�x��pPd�%X���G�=����5���P{�.�� LU[OZ��,�cG�0��m�w��d��~и,Fm&��j�MB�,��[��|d��[�0B%ݳ�e&>J�
e���V���E��ճ��qq�MІ5��� ���F��6Xi��Ip����}i��J�M]o��W�Q�RJvXQ��)����|GlP�Q�.E���f���wt!}֔1apvk:�m�z<�#�'��N`J��H����*:2<<��f�^.�R<bQ�d��Ӡ2�sJ�.{K��ӟ�KI�7���t_�ނ��M�|⽋^��7ls�=��u�!��<�	)��n�G��a��d^U
7��(C�
�2�x���e��:�E���c �^=���"@a��l�[l6��k�����2��N쫂׈��/���мc�d�R�~!MIO��U��?�r{Y�h#�<)Ț��� C@_�����x �r��壮�慫?~�֣������~CA����MX~��u~�� ����Z�����ZS��!����8����C�?}
��H�`>J�&J������s�� 5���y@��4�6"K�+�n�b%�^�_�k�lo�)�ha�x�''��k�{���U���w���#NY�`転��l��%��6�� 2vz�\R^Hh��Ӥ�7>ġ��;�8i��S�`/Ajs��Jf�����^�)����[@�!{�������q�Gxs4�_tFHrP:�b�v�'���V���s�6��Ѝ�ɫIl��1DO'�S!}^�$���Q�/b�����D��tW�ڰ�\l�d4��{n�Hߢ�:!���0L˿��]�"�Ԅ�-ܨ�>Y�a/ƹ6b �GEB�1�^���T&�e��"&�E]nF=ݔ��[�JF���\�a��|�JLu�QsXt�������!�D���n�V|c���j����o�>E.�� S؇�EC��n��aq�C���Em�sv8]�]'��t4k���aѐb��T����-�$1l/�7Fڽ%�8˚4�b�/����c$��Ȱ�z�)fv�
���o�i"����>ȓ��$��J� ����R���/��ؓݩ����m��+�K����TP����o��o�+l�j�	f6��Y:�1�{ez������T��T5�s]pGEZ���B"t�y̗M��4~��,W/+C�jsq�bM�zQj(�HGj.H_�7��L����I����˨�]��Dm'�K���	�#2L?�{�N��s��;Ts&,�;����z4���k��bN5���b]CtPt�<;��i�c�Bǜ@,7���c�q�bQ6�9�Cӆ�L}l��~��J�ٽj?H�2/�L�jj�Dڏ��ҡ�}�kIF����S>�Xf0�ª��&�[n�xۅ���}���iA 5E,�a�to�e�����$�A$/>+ư��ɱi��bЩF�1[gIi�O̳����~^;��l��=��~��ι�N�:��5�c��˓
� aEаYQ-����?��`eܪg��<47ݠ�����C�1���=O���x���()?��}��H�M]��r�N\4L2�K�jb�U+�3��U=�a�jY��Ѹ^��׶D��� �<O���1D��u�>�����Ƈr'bj�S6��||<��B�i#\#N��4�*n�B���c��Hv�Q5�1���= �x����D9>�}��tG��$�3A��߇��A�1I��y��j��� �? ��1i0�u���NtS��|�P�g|�X��6C/wJb>z�)��kgʢ�v��["鱊;�����I�S���.4��I�9_}��P��Xkֲ`@��Xb��.~���0r��W�.-0MU[����"�?��v>���~z	�7��v7+V��y)
%1�܎��޻�;>���C�\V��9�N+�r�8�D��N3Dg�MN)�wo�܇����iT���=��yxx����S㫫�}��4,b�R���(�J���0�M��JZA7G�|}�J�������u-�k:�ZN|IJ=/ē
:�,D
A_鶴��Vi`�Q0yF<�(M0�!=�|������ (�Tޏ����ư��4�-�213��������Z�⭨<yI\2VqB/�v}�r���r���WI&D/J�c���N�Wbɠ�?�'�
�$�w9vb���X��|��	ѷ�C�_8Qi�Q�O����P ���b��?*C���j��������5䣚t�T%k����p{! }�S��tE�/�X�p��˪q� ��nc�m���bn�U�P�a���	�t����c&���@�X���5�*LR���[�?���Q�!��<�@D��t�X�rͺ�m?�����^,8#!-Ҫ���G�G��[�a�n����5�r���87R������� �!��?q��V��r��~U>x�jK��>sޮ�"�9���P�.h�	��L�ܜ�Bn%5�	������af�ؒA׌��A��!���_m�;?o�Z��o9ǥ`d��6�(���߱����K�
 �Nthz �B����o�Jd���^'�d��!\NMR�� EW�q��BꄨMI4Q��_������Q�AT�t�f�U4�{Z���� ��:�����5l0�pd~r�[wCC��ʃD��������Iad����Uwo�?B�
)�H1��wٌ�xl��)�����E>���o������� ���%ޜ�g�6����o�ы�.���c����\���D��2���Gt`�ܹ~w����ncΣ�R���F-@�!���'m�YrM;�����������w���{�7�j1��&��ٌ�x��-�Π�� ��b+H��?�u�eMo&|���\��CZ��h�q�4X��ɴ�G���nL>�2��u9����|�=�q���xS;'��iq+B$��s6:�����f�r�ɸ >�����cZ�����6c�ӭĆ��B�o{Z?�iޒ���|�ξ'���thl�
xa�B �#��u�qׁ,e��XW�+��?N9�v�] �>�t�B]��AFd��z�cIa��#@Iq�%f���|��YK�	.n�[>x�$�����{��p�-r_R����S"��zez�9�!eN��	y����H���U�b���h^��qH�ǭû����?��kX�WX�C��h���%u`ɪ�b��~ rva�,r�g�.$��9a!?��u������T�<�u�`n(P��d
,we�a��
Y'cG�yj<s>z3�����y���+]4��R%��ԭz�t��D3aQ�4]�`����结yj�:��3��u|�KP�e�E`����ܟ���h�N��������{ȼ�amuTW)���@�%.�n%M:G� ��p=���3�4���T�}������D��M���$/�v�H^��
H��h�v�±�u
�j��nۢ�*�� �VNw��3�S'vS܎�
'�n$6V:�'{��,;,�����G���":QP�+�ǎ����9@s����w�j/]J2��<� ���b9R"�a�J3�8q�._��W���J{}\0CV����-��H_���R����M~=Ē�r�[�c���rǰgw�_&��������,df��#esE��hۆ,��0<[����λ��:�ܩH�m�:�:4�F�^a����fʫ�P�oaX'6a���c<YB>���G̿��r�p��}��?U\:�m�&�'�5�W���dZ��MNwu������ֲb����WD��j���D�`m##�gl�C		�i��-ܑ ���"o����ٝ ��۫�m!���<+�z1Nz�Ͳ�Tj]fl�:�D!��y�z�i����¿��vpr{����R����]�g#��ޙ?fc	D���m���3d]��߫�b�9]k�R��0G2�f#T!Μ��u��u�yi�Qp��$�X_����f�kJB='��ϻ9}~6Ux�A�f,�{�$�<�N&F�f6�kpe���§ψ���jh�EN�YdZ7?�>����aT�9.ԇ�Z��3K%���<B~,�ޯ(ؤl��VT9�{�d��L��7(�������Fb�5"�)}o#NU��R���=ۃ�mC��f�7�����N�ҙH�W�|��F�̦P_#شh���^ 8c��h�,6�R�?�btDewg"В� ř�I�/���2g��2�d>��jy�����^~l�2��A�_��!��]�/�d�|c�W�l�P���I\]�ZE'�-��������l�k��i8ϕ�m��a
��M��`��V]��> c�����Og]���cn��,:S04W�����~����������H�݌2mJ��ҝi������r'�&�T��6���^$tI�aQ�@�T�̡A�TLOD�=�`C�Շ��?C1��h�f�D���n1�ڜ��j¹�ffa]�t8�8"��]`Y�Zj�'��q��Cwf��8�1 �<�Z�����I�@AY/A[ꑃy�;]�n>��`�,�����9�ZM5�.���1@h���:ʽK՗��Qs2#ӔS�������\Q澧���^�Y��Oe?hF۱բ8 ��6�9/��6�}�L��u�k��+5����Au�S�ȩ|7�	��88���t�S�`���qGH8d�eh[4rc�}B���mh<ue��+0b =&�YqwW�d�(DƯ}�`�C�0h�#c�6*7�}�4tܧ
^���"��M�$ #s�4t�N㎱<ъ ��GX���h���
Z]���X~��T�M��������:��+	%�O���~��B��I�N���=6�f1�����0��CR�;��{��U+��*\v�s݈�xH/� Ԗ���]fMJU��� �y/9�2jCc-)���b��5�5ɭ��� h�g<��M��q,�R�VA%� ��\!���&���WV�;1�Lwhr���s/�eNj��T��5��߸���>�Y��@EW��m�um�w����4jL�b���$!ea��J�Uh6��gB3�{�(�ml�>�g}S�!�Ws���Ϡ�����%)i :�M|�����4V�d���g82kz���;��i�9���)��p�p"�T6�y����J��F�ex��4�,S��LΑ,�B��8.�G{�Oc�M�(u�c=�]\���IOI[F�l�x���(�Ȑc�APE{� ���@���Xm�|X*ù��5w�+i1e���GXS(Li*C� �􄪺����
k�4:3_����t���]����?J�JI;țO0!>�?O��y�6�\�o ���h�V�Z�/}6�gx��^�۰�A!恖t(1���<ݞ9�<Q��'������.�+ٽ�WqWa�A�|�����ߣk9��UaML�sG�5=�R�J_Λ�+`���v�l}��6H|l�g_������kFnE8��v���p���ԭ��쩞iٍBy+���`\{"�������"aw���7��6�0�s�fs,���%W� hf��0g�}
H�en������y�>ϩ�ysUSS�
-Z"S�_`��Y��f�eh���@%:�'/��l���ωȾ�$�h)�[;�An��vjj��ipNy�`��O��Gg�8�]M��ISi�d���2R��G�2��j9p��������:�Z[ΈRJf:K��ȟ��I�I�4?ygZ/Q�9��"�no%������:�ıs+iMȘ��E|�w�����-��b24������3Ց_}F��z�Y)�ĩȭA�˸�Q��OE��5�.��z@�>fB�+(��"I��ԿM����ܱ�פ!�G�V�=6h���P���,�n���'� H��4*mj[,�
iPI�BGtw}�	YX�W�9������I5&����+�R�v,] M��~��n���4|t;��D'�SvZP�WyB��g�;�$���WY����*W� b\Ȳ��m
������#���Y�^��]6��1���da�G����y<�����6jR"�I��~ޤ�Ĭ�"ى;��(��SRW\:���M��;:%�VZ��۝��l����fm2t&s�%�B�����C��#��f��D��)�L��R~�c�ew7ϣR�d3.壏�@)t��\A��e�X��ut��`�E�;Dq��_�^��/��UB��S��PE4|���:�Ɛ\�%��M��5$��۬dY�肢�QU��m�[�U�i4'�F�S�q��1�V��K�'֎��ߢb��5�Y�KK"R��Q���-������D	Z'G�t����֪9V�2m�x�k��&[̒�i���Rs���zM��g1S�P��t�AҸ���^�bh~fq�+��]�w-ԝG�xCИ2�;�aB&�^�S5"��V�$��yB�_|�I�hɽ�d@ e络@i��'��b�,�����cCv����Cg������DnF*6{܄l��"Ϝ/�Gߴ�S�d�"khTx[Tmǝmz����nNV��XVY|�*
ʳxf���Wan������ D��
ܗ�
Qng���
���`��8��Q���^�$�ƭ����mt!����M��0�:ص{���#!r�;Gw�8[c/�]>a"( ��39� #6��5��KfR����:���e"�K��~�:�8`���P��F�y�r�
j*!'D �5U�B���Z���~lA��ECԵ{ܩ`�C@ԭ�;�ȱ���mY�5��S�K����8Y\�ߡ`"�q��8k�-힘�}��ˌMa��M�����[�<+��Yo��6 �S&&�<^B��ۭ�x�d�^��K�+�f�Z��:�#�I�ED t`/�1ѮЛ�S!�e.2a:/����?%�N�Ps:ׅA�����e�0-(���k[����j�7>r�,J�����i��O��p�{�Nb3~��s�kbGMK����6|��O�T^�,�z[ ryKI��5d^���<ܾ
2��R3�ok��m�g{���Pҷo�.l�����<`���?�s�����-f��ݔ�"r��t�Ο��j�K�'��ʕb�/��o=��qL���ٌ�.@w&�|&d�`n^���c���y�(��C�)#�.0���jxX�β���V��R�:�)�ژXy�� XfK�1Q�I��1῾��
�v s1�;:
"�bO��V���Q�xl�~��z��Ѯu���I�2nJ�}�Q=��W{!x^���?�0���f�:gn��$�g��
�\G3�-䡱��\D �!�B;�E����˩���Du���'�%f�nbT�x�C1��Uf�m)��)1�����2np�|^f𻠦�h �������6��j@�1�3���w)IBㆦE����_9`���9N�`ū+���	��3>+�ĹNZ(���[��OX?"?C�)�!aD���J��69��4~Ȍ��J�|�R�����n�����ʋ���6�-��L�:kgA�(Q�h���QR-!�	�ā���dCO� ��ݱ�h�Tq���!��HT�s|�Ͷqi�Ģ!�����y��a���ԟ�lY�+9T��7�,���ѳ7��WDu�(��1�\H-b��G�8�M�bj8!��wh&L�<������;���8V߄����{u2�4$��'�����+�e�l�́+�򐣏���x�d��C��!�T���+-�S��8?�hz��J��РՃ �G�Q�8�y�X�?��i60�i�r*���(N�׷�V6ME쵾���U�1S��K�g�n	ѭ��T���Q���s�FɲJ��=v΍euU���������Iq�m`�t4_����{����|��Os�V����\���
#��������J��#:dJQ�S̉{=�0S�S'���J�ŝḴ<� �V����� �y��@��I1v{�攎�yb{�^c�N��t�Mq��
�"1�n�v�Azx���:{E�J���8�iǄ��rHd������ ?�F/�U7�Tܦ{�]0L � zw��]�n�!p#;�� �<�M_�UBc"*���W�:�B�߻2��-��Tō�O��^I�0LP���۠���̛�(c�q4ϼ�],נ�����n�h�sQ�Ͽg�`��˼Z���a��3������
�N�э��Y��0=����(t�*�$������E����	ցL���OG)*�Ε<;����ѱ	�sZ�D��[\h-��r%6H�Z���O�N��y3�����I5���Aj�Ъ��]e�Ī�}r�h������Wb5&���Ei���Hg��*�PfE �ڢ;�S$�>Ù��&J{�yb���;I�]�Vw��Z͝Gj�i�I�S�l�Eh��^��MJ��(�#�D��kA�wa�A�/�'�Y���*��4ɝ�����O�ӏ����0��S�o?V�O�S��a��t��@���K���N���9� �"�aG����w���(�,l���%���g�`|���3�M���'�Ĭ_�M��d"�a���Z_���)����yz�MP��m�M2�b���2��ڱV�"O���h��K����8�.�P'&������0쉛����v�l��:J�3�AK��0'Y�L�8�Ў/ߥ��U�����-Z)��n��v2����w�g ���0f-`��y�\���S>����iaK�$q#�`7*�H�Le�Y�PQNF���-�މ�� 2�yb�{B���I]���'$�0[����D ��X�����yjT׌���9�R�H)�b*�n�˒�,L0�>�w��-�IY���[7&�	���bH����	*�.l��$i S��h�L�dO��D+�?U��x����J�Q0��SW|W_b~w�Y�4�O~�c�;� �Ӧ����l�3rьDs˲��,�l�I�.ը����I�	3)����`��ҋ����!A�nw�j���<�z�N��"9�|K�M����6�|�!�@#%ɮ3�Q49t�*Tu�c6`�C���͇�$Ř�e5➊5�T"t�׮WY�R��͈/s��� �{Eˣ1��8l]M Sz�Q�v���̽��O~E�J,Dg��|�{w��|ؠ�����a�q�dܺ�ZQ��������7�0>=i(�r"�n~|,�X�����B�M��-������JÏX�8R��Zwݬ�����P���T��sM�u)�{�ݷ��I��(}J�~Ռ0����7�F (0^|�)��ו��MO@��'B~XIu!�aR��⟙ُr}Q;�f��2v�y�H�1͔O1�$�8�Pg�:Z��M�A������
��R	�r�j �/�q�.v��"sVO�K�{�_�h�c�v�#�Ce�тCt4�����x ��낵�n.Gt���8f��M��>�5�Rd>�)�~=@��'ҝf �������� 2��
ZX?�F����L����2R�NV��kؼ*�98Y�_G��'��6��O���%�T����b�6�_bqX�0�3K�G�é�����/�8l�y�	]C�&I�ֿ8^6L�m�f�$���SIG�9�� �#��I�5w��0��GO�Ɠ`��[ܤ�*����$��z��a@�R�>l��^�]&I�E�;gW&t*L�}O�ʕV���i�j12J0��|��*֊۔ �նc�z�p8;B�N$6�τ�W���97�����t�ZYD�O�ÿ�V���`����yo�W��,=�f<g���7Gu�Z�R���t/v89�b`�v�zga�v;�
����hL�PCG\w��Q�	�C��h[~�L��t`Un�VxY�iKK��sSF`j8E��#7��o��<q@����r�Fe�Q.���;��x&1c��KhWU�;@zT;$�&x�)b��/ +"��9�f�'����ꏑAF{��� K�
er����׻�r��LS�Z_��T��+Dձ��g��s� ��;P�z7�o����\^��٧��A#�;_db�V㚍�(��@��A
�Ld#���;_��^��}�H|�|�LL�<9Ն�_�ϖ�5DQYA�:HO�8C�<p��#��Q�}W"�0����5D����Op{�o����FqH��V�� �^�m	�
�2�Δ��r�I�۷�4L�%�s���^/U0�V����y�I�Ƨ��tS�)L�Իޒo�BxM-��b��˴���֘��n�ԒO��l +iQ����V݈бD�M�jK�_j��;%,�sua1���H�΂!(�I%S��B�d���{!Ի�źh[UF+��&S�π��{��{�Sڰ�
���t5��q���	���H�)\n�#c^a�	�������HXu%Ρ˝���j���;��~I�w��!+���MJBrn$��������#�j#����g����v)���^Cr���c��-qQg��T;�T��v3-EA[c�@���K**
ґ���:yF%�(�,@��(�c��IP��蕢mr(F���*&�]���a�I�K�s^"��{�S�A��0����:t�>棰���k�=���r_9��0Mr�!r�L�X�IZ�O~�a�W�h,�u/��F��{�L�d�u@���c��VΨ-(��w��N�!aO� ����A�w</�	O���C1�>8t��d�������q}��H{瘏$IZK��J�l���-�����?�L:𭱆�#N�4��n,ݻ��I���1�9a�U
�	m}-q�W��c�A�/�o�EXJ��u�ļ~�G�#W�-\�Ci�e��Fj�!#���HD�h8b�'ߌ������M���zibr�Q���\!�ɳ	�|FT�2Z#�j΃��R�!΅j	�~	���Ƨ�y�V�IX�q7���\��Eyu	�����JK��	/��]��q*����6^��YV`���1D8����\+���bM�}��g%�Y�cQC��V�?D��2u���}���~g2���K^����|w�E�O�-�4yt��`"���yb)��!j�2uS��7��Ճ(��w�t��L��1�߮X�����Z�hj���z�k�,���3�J�y�"Y>@�9������^v�TA�!"\�����	��Z���P��m��j��]�Bu�8�^Ħ_��>��ͫ�	v�<U��p�
�yh�ݘ��)[�ܸ!6�-
�GV��&aw�����J�,��U _�K�.�5�g����8o����5�"�db3�j2�xN;�Dt�n6��W�x&yѽUj��#N2�5�E��Q�l�$�����Fq�/wE�F�Pw�<"�T��i�؆
���o2#yRK��5>y���.��hy`ʐ�uv�|���,?�(�$�p�ݣ�:��T}������2��Sս�L�^�ڱ��c�*K�K���Y��0I4�M ��$������U3^��j4E'�M�&�CG-�aد�aMh�P�ST�Ph⺚�@{�<e�I��m�-� "��1� ���ދ�`vt��������A�#���>pc��rk����ޗt����)G��re�N��cS�u�fҘ��[���0&mG�[lcہ�@�K!a"�����-�8*�����\R�r��i�Hv���cٛ����0�}������d�DtQvV`�� ������[�>�	��)N=<���)��q�o�tk���TB�߽������̶��E�C��c$t�&5�˼<��S�گ �}����&�-�#��Ú�~B2���̹�=}=��6p�eo��y%=wZ���rD��s��ydwx�B�.ؓ�v���+���sW�S-��Q��\9���O2z�����\R�t�<�v�<x"�)���a��N�|vV�4h8��CB��§���X(i��r)�EE]2�E���W1Ff���1��@�����N5�,��
#���N���O��t_ڎmF��Y������À��ja�6����J~��>�E��E6Ɲ�Q�ف?��Q���ڂ�����2�xik�3l�I����T�:��+0"�o<��_ݪ��i���0���ގuY������.�Jn[M��uVn��8�sU<����O��%%��wQ��ӹX[�i��F�c �+�
��wu#У�<U�h�Q��@u2ҸXv;ă������&&�%x����%e�|?�NQ�l�J�dA��\������ݐ6Dm'�I?��{]~���]%
(	�����2��u,�Pg���{R��U�ZO���5Zӻ���!�.�Ճ�i?��+	?f漄O� 8��`i��7�S�rA/e��O����qo)�vOH����cːBl�緔���6��N���L��x���t����{Y����B�DWa�O�H�^IN�:y�����,����݋��<��Y7����^ڊ� ��XN���R�tR��^,2F\��WTA���Vu��\�n�HAuC'��O�P��Gf��S*�}��6�2'^����QL�_���k����
��3���b��+թ	�^]K~7�x��.
c~.Oǿ��y��C+L��u>HuF}[ٛ���uJf�2���$����ě��+���R�o'�t��3	u��f"�i�'�Ux ~A�vt�4RDu"ꇺ3L��g�N���� �E�M���3���<��7�Ln���QK�ɷ��� �L$�c(ͺ�D ����~��{1y&�JG��܇�4��O\�Y���+G��O�`&���`JDǺ��O+� �ؖ_�B2ݗ����F�l3�������+�����/�-Hc.	Y��}��S'0�pі��}_U�.H$R	�׀��?���i�RO!�0�:7�'�IY<�3/�D�>=:��ݩ,�{��s�u�m��6P��E_�w�TaK؆-Qmob�ȃ��k��[| ��PkO٨��;��x:)�Ch����s��e�`��^�>� ��/j���<�s���������9۽��<M����u!�% ���6�.F]��KtUQ������'� {$������5 zR?E׃35CE�
"beq{�
�C>��ze	�^(˟ a17����@��[jw��t�"���>٧�򻼇����h�	���G���jҦV ��]�	� �U���m��HXb�D�c��CP�C�*���#%�T˨�c�R��!/%��GKظ^���0Hsnj��$4(������. bӬ�f�N��h��-�H[w�x�#g�ר4����s��%\�.�:R�m��HȑE����P	�fHƋ�&jY�����²�ϺR��D/{�{٘��nh]�6J(տxOn�(�UI��&�g�r����┏\��\O�nLp�v/���V�ٿ���@n�82es3A��,2�r�l>N�d1L���Ej(��7_��������,v�,̛R]6�`��k�'���j��3'+8�̸,�f7�%ȫ�/�32 �V92�,ıO���0�Yeb�ݠ�����Ӄz��0?W��ލX��ѽ��v��{�ug�g�P�C�'��S�&�7���
������hLN����(D����z�\|e���$����(�JuB��~�UL(Z��[�jF�$0���"�~=+�/��P�g�PY�7TO3��x��$�v�ei"�ڍ-'I�CS"n�R�O#�xT=���[�#�y
�;�H�n#H�I7d�k���ک��Dl�tnh���m��F�a�6�3�!��7Y�X}�)�)�n��O��Q�d�-a��-�Ќǡ>C�|I�v(6H(���`�a
�ݚO���Ć��9�kjw`�Jy���o��ejܬЕd��������,EHS�V%uq?#�H�g�$�?GTUK���Z���5%ul����\�-��<�	�>I���Ӳ��C��,��nnN�ze���o�K�Ţ�ǹh&xb�W���E	F�O�f��������Av�JrrB���Ji��On��r��KO�݃��Lu����5��X�V�vF� ( ��i wr�*~*���f�1�$׺mh�볡�e���}�ž�2=�&� �c�[&bA��ٕ�I���"����$d>��e��Q�� s��uQ���j�S��h
�e����ښC\��E*����dsST��v��t��p6!���w1Q�t�yX�@���~�53c����H7��E9�H��b�wX@���N���z��M��r3��)�D>�����ɍ'w�2}�P]���1^#R-�z���;���G��X;��,�m�����|р!/�3�p��6Lߺ��<��a��q�/]qo���L���G[�B�'�Y2��,�~��X���4�=	b���5�&��L�`fTZfM[ɲ�T����B��
%϶'�I�S��]*NJo���Gf@�7>;��!kZŶP�}��e�E||�G� ��C=Ҹ���?�����V�?o
ZR�Y��2�G��8K[ �[T{�XGR��'�)��?� �s�oC�<��`Zq�D���%�d~g��R(���׻\��ժ��baCω*>���$�x�\�8Rr_�&��E	��)��0����*��Q@$G1/nA�Te}�����d���uw
�����V��[@�R��Q�6��Y&�༈?�WH<�9-n�%��S}*��o�D릏���\��L�b]�6�n����Z���l��s��@�1��;t�^A�/CH��\��s����YS�je5k�	���Ɍ���Z�2�%�F���|����A"��t�>�#o������&�^jͣ铎T��۸��eZCz�@����hˊ��* �A�K׎k-xV[c���}���Qg��q�_�$T�V6��`He;.S�]%���vDKGګ�Np���\A�:Ґ���$%�V�� $�Mw��)mb�N�5+��UQ���xE�Τ&q�`����~�x��z{��)}�A�-%��)߻G����KX���2>낀�)�ӑZ,e�Q����B㒜G��b�������2-��ˠ??sr�K�V�G_�A!E`�\OX��G�*��U ��#��L���^6�y=,5��.�A� C�E֟���U������ڝi���^��X�Kr��B�e�&�q��PSQ����M�*�L,������גּ�;a�֊��j�2*<���͈o*�0?2�#
�2�c��x��<���!X��|-45{�c�Qe��c�<8��ZoEOم��_E��:ކ���_>��fl�}(�)T������s��U�d�k�kr��M��Ss��>�Tx��ݸ��p+��K���q� Er(Qt��?Lh =e�����w WvO������vX�]�o+GN�VB}Ň�QmSn�#������$���l�W��K�W���fq�=��;�������N-�����/C�~E/X�6'j?Ͻ ��=�-kZB��]/�������'}6T��",��;������ϭv�6bN+b�*�/��,`��N������ہ�y�������|Y�E}O��O�� ��U��S�7%��Rv��]�\��A>��/]5���1�J-���I��[�d#��Bj��MK�A]���������������떌��E����
�r�9q_a��#�Mp6�\�56G�s��e8��wj�����MU��j�J'��Bb\>T�u1�MOn|D_0|K^�t�~Z(��^������K��+L�؂n�ਠ�uVŒ~�n�pY>uH�K� O=�Ѣ��	�\�c���T�\�^��E(^F���i�#}ݙ��׼꒝�ޏ�֬��v^�b�J����M�X9o�qwMP4h5�YXfpf G�� ���^y�Q:���{f�]l����Ek�>�	���i}�X�F%e9���uׁ"s�w+���*���wz����P�y����D頪Ȁð ��,�[ix�0>���rAd����W�O�W1�>�Cͺ�}\ ���Z���G�ni��+h��s�v:00�F�k��l{�q���"�^v
�Vd����J4[��7�`��I�4)���KD�=����`��@Fwѓ�W��"�Կ��
)L~���-n*ta7Rb�%��!1�[�7R3
��ȉe�Ⱦ���[ ����-i�[�c��%�f�߇�|`=��Z�K/R+7�{���b���5ˣ�5Y�NH�X�I��R2���&�[&vI�_�S�n�"����i!2o1T�}�̵O���)P�R��w��7�--�Q*@͔=P�8�8k��s�̎t�Fh�tAqv�I�e�V��	S�������LE�'>y	��Yk���Z��s�3"�S��O�i�=y=@=��mI�
�f� W�D�vك�k�#���<,G�G+��[��k��vj�
L����_�K~��	�'����}U���C���[8� ,v�m��yAz�pri�cl���l�y�0J�r��a���&~�`g��:H_u��+髚���l;�8acn.�{����c9������$��-�Dl(bf9S�xa�W�$�0��y�K%�����Ɵ�!>fB�qa���{�f�*t�t��̗��A�����j����`X�&��o�D�@���K�V��R
n�i�t�^��B|o^o�Ǒ�m�^k�MH�S��;�Q �d������yJ���V<	1�͵�e�s�*����RyƩ�]'�ڌ�'�ᴴ��dskɟy��F&���=l�F��+>�:e0��������籤�oiYL(��H�cR�in�L�*����b ����/J�d5璖�qZ�ggNT�9��:���ז���:��wL�⇦������
%����	s�R`�r`\�-�2��A�F{T�Y����N݋��e�G�/;�E=x2�^�ظ������	�,�D���
}�߶P�1��V{"��_�glZP��Tչ����R�����Ά��ڄʗ �$R�^�x��V��~|Yc����̯@��S�P��ubS���&P�7���F$�̪Ɣ��"����к�SX�^� �ͫ0;���hj��=����N��-��w������D�Pb���#�̂��xvUM��,+�w9pDi��&|I�3m3�=}�EC����v���d�	�(��E�bv�io���&��ћ`"D��fu=4���L�g�ґͳ�V�6��CQ	{Y�����c��Ũ �R���&�1��� N�Q������;Zzٴ��7����,G��������B2=N�-�,���`�}�xcrJ�HK�5�Z����|�����FR]{sR1J#Sʚw���Ѝ]����}1ԒgЗ-.�v>[�'�g��<p�g �c��}b:&>�/&܎���@*�g�~ݽ�/h�@a��!D�����7M��Oj�J�J/�/��\��/V�:��G����2Q�����Bgw��
e{��87J�
�l�p�����:h��W���,��-��%����ʇ�!�T���7���fR�՚��?�C�_KBLhWhTY�@-9LF����mk�����&����O���e&���e<�u�ZW �9�}iw��# oø2F�<�h
6�(wCU�0���$�䊎q�\��#�ߞ��m��TO�5��Sw?Al��S��6v�v���'i^f�g	%l�@b'�%Kr�M���o7x�rֵ��F��B���' ���wX�� ;�m̎��q(]oT"�Y����e2�De����N����!��4�G�ԭOG��(��Ƿ;��=�&w�y[��>`��w�۠�kw?�d4����1Y�ו$�iD��I��g�ڋ��l�#�rn��4�6�bL�0�"&?m��C#!$�>x���#�1�#�ksZ+��bM��&
\��E\B�ປe}'?�<c�YY_p��Z�0�޻��X�X�s>7�Ҭ��d)2�Q�����_���
�A�?�Դ�M��1��'��`גx����>}-f�O�S.�-ƕ�0��8KD����/�7��z��Zƺ	���Wl��|RVh�h^��\b�R��s�g	VK�a�*"�$����c^EЪ�G.��
R�~���O���"��Oq�
�:��ը��<nvG�D5p����
v0Z�n�����8����W��\*b�<8fmXYHd'ƪ]E�}ZL�ج~M�v|��8֤�����"�����p�|�ȶW4O*�w؇�hEBv2$17�*+�A��JG��C��!�߅tʙ2FA��SZo9�\ya��c�l�������l94-���-r��R�K������9p䬮��U>�]	H���19��ق��lGeo��?~���鑖#��,��%;R� Ì����"��ហu��,M����lP�`T<��(��d�RUy�Jnu��X0'"���B�O@�2!j��R�R����8�H�	��br��"�x�K����D���oR��Q��Sj�W\ؘ=�q�����_����7	/L�V�'u�+H�B���b���L*W�i��?&�ཏ���Gd9����:,�u~H#�,`0�ּ�8A"�v_]\��<1�l+kKk^�)�7��-�#�Fd�	��'m[����b�,�/
"s�R�Dn�HvD�1o�����QOQK�ܢ`|lR�L�|'�]���w�!��M��x2z�
����K�Sx�Ԉ���1?��k�ihN��j@<*���]jo�_����@X���U��BT�̥)1�r3���g�NdR$� �.l.m`N��)9���nf/�gڳ4:�u5,�J5�m�sI�q�%�j8\��n�: �Mi�j�����YQ�t��]Ζ������p<�ÿWPrS���݃�.�L��9�8z�ǒ��!��f3`��@��iZt�h���Y�t�vߺx�>�Zb}�1�������/��$"߬ ����G�.
v�X�C�B�S]+?:9�m�!�%��<Wj�l������X��]�J�
�e�ሣ����9&&�@F��=�ThF��.�QD�G���,�z2zEG���7÷/�mw�8��t��M�$���T�Wqk\��!�Pep3��@y2���]"I{��&�t�����t�;��xJm��5��u]�wYru? EIРs!Z�އ��s� S൐g�A1�c6��f�>J��-ߞҕ��"'[�%��m�wYQ�ڠ�K�������֦^@��?b��f�������K�Z���Rt.!j1���ut��O���="��/l+��mڝW� s7V��2����u��<�p$f�C�6B���.��Ns��g.!��vR�\3ӱ�|�̍V͑�y7O�@?���rrݗu�����Y�=Ƽ�d�JM���`�b�df��
:(]�6�·z�-�0��?������B��\I���Heh�I�e��=2:�	P�e
���(k�C�>�t�r���2���~Hj���_LR��T�
�5�Kփ��JHA��rW�vjE�q����Z�Au+&9IB��\F��M���^�]�\�0xi|I�dL�B,H
ü�/ �s�<�\���A���	Zs���M�G�5_��tI�Tb��r�������f�FnM�	��(h0cSBi?)B��~֮�7�Ӊ�f]�|S/;�P�{�H��%v0�!�������'v���2�v1-�i:H{��_E���.��)�d���ou�V�GR�l��)��B�o��b9��5��2!E�۽�M~�Cj�*����0�t��>E*U��X�i�(u���q���k�4���Q�f�Y:�&'$��x�ca�;P:I�#��տ5\�JL���r�O�8�9�$�����1O6�Б���t��!==�w@���l��v��/8����en��0�ze"[ߨSj"�����s�Mz~��"7T���:9=*����1 �R�t<� )]}�5��F����oW�M06)Ji�=&��c�팺������z���a��e����N{�L�M�!#�'q�%5������>�EĶI	��Ѝ��ǒD�S@�ad#i�����u�$JΏ��Γo]�e�+ڛ�!ғɺ�#D������!�0��~)�<_��ɱ8U� ������Q�91�"��$o���<ةm@s�ahU�Vx]�ۀ+���Y(���L0�ƛ65X���ҞtLb��H�!r��zS� Ҫ�&K<#�I��0��@�ko*٤�\ݶ��+|�4�'��U�|��@��w�svʟ�b�s�,�!�J=$����>��ş������Rf͙���䨀M_��}3��/�@�_��:_G9�u�t�C��n��p�x��`uof��EZ���I�B���X���p����Ȃ{�8'��T��Xjq���׍�2ZV0q���V2q���[\�$���=4����Ɲ"��n
�;��ߧ�����_]��ȶ�V��S������gso�����_f�|�ROi�3��t<0~WZ
U^>|S�y:�ɔ��{���%.\	)��~z�w0�X�<��1���D�
��'���t�s^<9$��Ýhtn�L�m�pG�W�t�&�辨�W��b��7�q��CR����Ct	�hJ5j���
h$�B��$t����]7y�|]�cJ��&ߑF@�x^�t�\\���s4��}��#�N�f�?�4�Xm"0X��.d��Qӌ�e���@U��`��)�b�x�\�򕫨U@�=0cE�]�$9{�[2`�f�ǟd�$����!��c��zUԝ�XG[_	 �,�4���e��f����|��\��C���G�cKP6�G�:�~��=���Z����ຐ�F������ϰ$03��K��gn ���nj�(�v��B߱! �R⩎��M�!Ѭd�8���|"��՞�|���&�
*�O�;:��x��.6�1�"t�Zj�
�����8�{d��5�|zz�w��9��.����S7���7գ4��������1U�ԍu�a��G�l!�mZB*8?D_%Ѐ\Ʒ �(q���][�#-����"�֡�*Iۏ�}L�m���-�eZ����1}ϞWE�^���v�?z'x����ݪ��?ꤲ ƨH�j/�7�I>l����-;�����5��7�%a|��%8o�1�ĥ�]}�S�3#�f�]Ѭ3��
�t-�9�<n~Sɜ8���܈�mkk��禉�:l_�zP�@�j�C�
GX0ϐ6
7+��P�
��>����vu�	��+<bʹ�ܝ춥�Y�B�,7x�q�$�����	ڦ��KU���kgj��
����D0���x~�|]z3=��Tr��&�BC1�� x�(�K��v0n����:�154��yZ�Q��V�����?�:H1o��NI?al�)~��d��ea�E���pw�����O�Q�o�P�Jñ�9�n?��3kC��v�w�lj|�KSg\0�K(奦�NLP���ǋ�?������F �}'��I�Țn˿%ۍ=d�i��HѮ5f�0mN�����!1�*�����n����No1�YI@��hm?��V6�b����x�\�e�2�%$I�k\�G�A��	�'�6 &O�E�YC9��W��K���4��61��d��WSo�K��8Q d�qp��#^�Zn��>&��R7;k��ĀY0^ԟ.�KÕ�9��,j&#�cZ��b]����2�:�S��	���c9�
E��]��=5�G�G�%�YCc�$IyY(G�w����)�8K�j(��5~v��/�ȝ5.:��!_�x�2�OJ�q�utB��#ˠ�*����h甤g3���K�B����	�q�8
�"y:��l��X]f��b�-�ٷ �Qe �ar������]�K���[�}�n��H�y�/Hջ���Ý5�~��rP����Z�����K��M\��	u{5��h� �U*��b�c־��������B��V�0q�����
HK�}�ԫ��0�(�&6^Q!+�� ���K�F3ZRe}��ra�ug�T�^ ���M^�;��k���Cֹ4��ԩ�T��"�va����
�l�Qc7s7�-���$g���A���I�>Ю��7�y���w�|�َ#LHo��_A�R���k]������>euQ�>7���=�b��s @��]��� L�e��D���d���>�0L�EH\��f�ן�3?R��x�w`ni�5;j��kea���;le16G�2�ϼ�Fu=�a��6z��`�!�_Q�-�nvׄ!���Fqv-�3�"^��0���U@�m��Y�Q�.���F�A���-w͒og��Ĉ��1k�O��C�$v�/V�d!o5ˀ�P�VڸG�5�4���ϟȤ�	��<9�����7LVp
�5���!��8ߢ��X�C�??�E��!5c��������:���R	h��ć
�tX���XI��l���Re7-!~�=�/�8�|�wQ��^<$����'M,��5w2LV�8��-���K���F%�E=���(���jB-:^/4��Y����Oņ#X�S��| �h𣲄�sF�) nt��$��wDx�NWCe�|#�m�L. �Bӻ`�yɓ�i���ʟu�P��s)EW��'v7����/{D����e�i:0:�`)�)�
4?_��l�ߑ�'�(���&Ki�u����WP������fDő��g�e����,�K�L�#�yc{ei�΁��v�c�u�[`�XY���\Nz!g=�:�xP� ��51��-�`��8^3�0�B��N%�)�#yQK+X6y�I��iH@��]^(.qa�*����վ�@x�4��|���@��&�7���G��i��؜z��w(���� �505+��3�>k;�H�~����r��������r��V��}e68�i鶯�'�ȽϢ�v'ħ�L囑t;!"&ٶ����[��!��<��%���z�)n.H��[4�	�!X䐯����sB�.�Ŵٞ�t�KK����N��hp�H�j N)�\�y؏��R}'(��#&{�B^�f�J�h5eTh�Z��AYw�6��E����Øn���81�%�c�`�����d�?䬳Du�'=�5�@�)U�R��\�����'�$��V�?��Ď���s$�S�?0"Z|>P�DG��z%�̪WD�q���;]r��f5ЕD�ڤ������Z�TsF�h��9Tj�^V�&��ER [�|��$Cq�tݫ��x���
��c^GoHU.	aQ��NX�������\z���ȣ�Y�����j��술"�� n]/|r~����|y�Ǵ�k#�]\F4]�4��{���jO�j�cT2���	a�JL:�R�r ��2��&�I=�6e�Au�6�ف\�mW[�}�l`ol�X��v��a�!5�@N`		���5����l���Ҳ�Η��Pp�����p�Y���fGӲ������:�zc��	W�6�҄X���!�S�7�y]����Z�-2	�hze1�8�4�/��ո��ֆ����±P�^�R`ǭg���X�����Q���n�'����=��E�+ޘ�F�U_� nP�݄$5����䤲�v��51�,�x�2㪪�7�qZej0XQ��M�<���{c��ǱȮ��b�g����p���#��:��~�
�q7E�@�LdS��
Ѿ��B)�^�p���I��mY�FrO{�	�.��M��~uQ�%�"������u|�=e�ӆ��(6�%!:B#����yH�j"O�2��!P�N��%%���-�-�tg�D��/���%*ÞW��/~�'�#����[ZeO��z�>��Q����T�I�n���V3���\�3.�Z%�cd8����0����d��'w�2��#A�����	��/~�Қo]�(3-��;�`�U|���gk4�֙v��a��I�Z0��GF� �s_���Y�%O/�����'�?��*�K&H����|ę~�%l�G�����$����ޜ����˾S�����+�L0�ޢ���Z��R�G�`��y�����,�)�4�8��{�4,�^�O����L*o�^�va!�J�o�ȉ���Y���c[�W�� 4|�r�R}ٱ�_6�K�=�"d?�uҋ�zZ�v[I���vR�`�s�ox�4%��`�= ��3R�9��W�t��4T�CҦ�.�Mc�,X[ho�,��j����й�G��T ;��Q9l�4n�dQٴA�q���6Ӣ1�	�ˆ؝���a�uF��4-C#�V	�KҞ5���tu�*��	 �܏4q���<QS9�
�������+��/��t��_ڻ�IJ�B�|�#��M��y�4�� �(�kciq�����\95��� ���xYy����M|��tԜ��b�~3�3VnD�4�>�,}.Q��Eq�mH<pz�P��8�pV($���E$7��8�gkC!.=�D�J�2K��X"��	���Ǵa3v���S�p�7ou����S�VN�ʆ+i��tB��J��G@��)9\�D�_9�d��V�YQ���8B������DP�U�FB�\�-:
 ��a	����̚3���^@]F{w��Y�G��N�Ԥ_�m��v�䗜|�\�l��r��JTyL��&j��R��������Y5�a�\�S�������$ᧂ��Z��Ȓ�`{���lٔ�k��S��ۢ;E[���C����]�SZ�$kB�����ώl.|�$�*�������G�[�Rǐ��ENTF�m<��r�Ol��T��w��:�����Z�x�IW���@�7�Itą�������i�i��wH嫗� ~�IZr?��=��M��+��I36?5~����)�7��(�o��~�
��`��ꔡu�(P
��l��@�;������Ѣ��%_�#�K�I6�I9�%6�hb�v�����c��e�F{ �l*�h"(�~c�[��ԴȈ�͗C�< ݳ�>�ݜ����7uE򦲛�����1m��#�{]v�n�S��C5,�Ê@3Sh�(K	d"�jk2\֍�"������9f�c� *�4��Dt�U�փ_���0�6�,�A4{�6�ǘ)�{}`I$[�F"�-���0֐��>㝠I�p��G�����^S�x"�#]��ð��@_ýA7?��u���t0w�flWgwF�������Ui�t�\P���&NE�;�#�����},W�u1�q|�3�U��z�r�V�����٭�l�{A�vi�ѮLc��<7�4����K�e]����.�aX\���u��&��;?�4�-4,�����,9�](�N6�����t��b�^pW��('GFyb k�Ǒ�Ib ���އ�0q]6��z�V��6�����:���׵
��x+��P���.L̙~�d!����@h��UR;s�3�f���]C�a���<Zj.,�i�s
���I
&�a[�	\.�l��[���@���G=M�}*~�
���:���T	Q���F�B6*��n2�e��ѝ�C�i^����mw`��WAuQ�d�Z�&�+�$j���X�}^q��^��u~Fd�t�����D N��f�7�8�����
�KW�Z��?g��џc���8�_#�]o��*��m����eAp�6w��*� XR�gd����l���+`�e�?��$��)�K��Ȑ5O�� :���5R��f|��v�`_�-�FX�Ft�R�o����K��ր�kC�?�j���2,� E�ܺ*�|{.���?F��]B�d)��� V[B��Qz���x3�:��MԤa��z�좦:�s?��L��'�ȉ0.�d�=�S�bQ n�-��*菎Rg 3h�.�c@qa��`Twj��Р�o)=ٶD�-�����r�a���SGg�����|�߻���%�ttO�D�iY'�{�R_n5!KoS���.G
|�#���q�؛t�4޻j�*��� _�寮e�LC$���k���ʴ�^��H\��gِ{Oˠ�x���N�Q�@~���պ���b�q~��J�_Pg)Rw�Nɀ�$�-���Bb�B�WK#��1j��Yd)�LT^P ��1�������
�w r
N�Ƌd��͗���ymK�YQ�}��q�=��5��@�)�ۢO���ⴊ�k�HX�Г�+�˫u�m6�C5�]�>
]�LKl=�[J���C�^6a/�.?��
X"W`?�� ]�[�7��X2I������Sn�Ƶ@������j�H��r%�u5�.Ym͜�̴�5�z�}���Z����Mh���>0&:z���.���i��;��m�i��B��!��L�)��Z��tʫ5n���W고�-#��*������l�2[?�t����^�����/����խ%��� ����B�v�lĄzE*�i���j��*�G�J�9��^ZCD����,` ؊
�)�H𮕳�m-��WE�<�EY�߀���0Zp������4��w�i��ף^��μ���T��̑H�q�Mr���q����?$v�y �y�]��k v�M���V"N��,##��p;��C$\��Y�2'P�~4٪�t��޵����Ͽ|��4]�L�̎s���=�m��z�T� OU��N�A �O�����I�/<yˬpR���#��������n��'�p%s��`�Y��1SiE�����r��ƪ��c%Z 80��#�B�&ш�݉��s�$�,��<E�nr�a���Epɶ�lmerQP��`2?\��A���P\��6�a��DDA�G*��) �%P*��0��f���d,?R��$^}�_2����qe�W~a� �5:���b�5�8e�v&���7��a��|y1�����a�
*߮=�4�����>��{����_��A[(�vDn#?�B����de0�kGygA|U��t������5,ۣE����3�,1z�]-ajw���H)�%�/]B�J����ǌS'dsj#����y���@�<y��,�1A(n�J���`ϬH �i�V�!�U˞�냴Wqt�ݕw�A[��xx{ƍ�[�LڵQ���?[ӼB<��c��T85¯��?�45A��]m	{��G.eS��yhPW[������3�e�1����T���vq�;�/k(��+>�\��M���7A� ��WhO�*���b����X��&��JZBE\�â�_<ǔ��
=��R�f�=-.��o-���b�j��gi��tCM�I��S�A������였.aa��63��v���\D-��o[y��)�()J���>z]��T��>��X5WQ��1> �ӑ���fJ����w�*�(��;�:�ř��7�G����{V�[^XU	���GkZa�u�4�y_�lu�/>P3	��&��ir����,]�h�)�g��~��TXJ�|�&��0B�*�1�҉(�T�9 �'+���~��	�u�nC�,%���,Ô9T�S2�ހ	�0�՞aĻ��o�M��s4 ���`�e����|��dL~(���0 �;�39�;$�^9˓慬��� �W����(��b�Q���"��SӋR�I����#z6ʕ%���� ň���w��U"�Z��Jd~���,K-x���Z
O�&���)�/>sjV��d��EW�!�xs��c�8�� �,�2�9���6��y45Π�����g�x%X���*.�� �#�$$�ݸ�`�3�E6+���УV�Z�"�?1@��Щ��A,�ծ�˸�<��q��`��xh�L�b���-�Ꞩ�E���g��9�NǰB�?Ϸ�.Om+?�ю|͖S\����+2��n�)P�K�1`!Ί0<��%�1&n�FE�b�u�@(�YYh�;�Sm��Q�ᅄJ~��~�.Yvk�q��$k�L�T�&9B&�h煨3lM;e���k��y�$��<���jv(ؼ7&E�V�1��t���5�Z;�8���is't�8�Ոf�e����\y��緍��.��&0ٴ0��m��L�b�Y�k�hk�ALe_���jD��2��-Y��<�>�]��.�:z	�|��P�e�i��[�Nn�)B}H6���CL�
��x�	��3�}���P̜��G��f,��nGtM͛.sD�W���z2-7���egv9a%N�}�p���ą�l�G�+�@ �5��=;�Ѧ�/V���<{���*��=��p���<۳��e���y�G;�2�Ǧ�X���Z���M�������X�j�4�C�<�jF����+��ޮFM��P���d68����U�����s�~�AHz|t�*C�ne�$�g��4����)��'�o�Y!3����욓pi��g�Xe��l�)��VR�B�ӡ�o �� �:9
�>�:S7 +?�l�.s�Ǜ�F?칵�qkO{TN7��d�1��`�d��.ٺ]�w˴���P��8ϳ���%�'����Vٗ�v鉔�U��>�lh|7!4^��8�9��{-RGN#��&7�%[u�3�9��������݆�b��	�P%�@dF
w�3�4<T��8�p�Qt������j���#���]���PT�!�ui�F͗vR�|�˼��12��\0�uA�Xd��MWCS[�ayl��K
nu(��h��I��2"�=�H�acB��(�{��>S�Ӛu�f�?/��J$ �4�Q���\Ō��0W���O!�y�۳|.�9x-��>D�P���8d��l�%RPC�Yڻ������ϼ4^��o�y/婜~-��s��K����t[K9�3��;
r !
LTfCO�Y���tea�c��Qm��7#?�ҩ�[�{ծ_�ꏍ���E�S����&RQ���2K뱀��&f-8֯ă�f+i}r�Й����Z�]�*�Sx���*�&Os����83� ����ni��}2��Z2�o�5>��m�9��q���m�%�큆k�.�6��
/� ��m� �Y���;˴s�<@��1R3����3��7kx��F쓼^����x��ʲ	|;�~�|)V�	��[NUz$�(�4-\�	�W��i�6$*d�qG		TG֞Gh/s_O�<��1��h/�9��������;�;���y뒅��^�K�	n��k�����Bc���1�I��nTx.$4"�����#�l��y�g�=c�$��}Gu��s)�a�,Q[�Gu%�\�U՟�F�"�f��΢���2��h��ٔ]��9�7F��sMԋ�z�G�=�Y�|��s�?h�ȏ���W�6
�h]�����f�0��m!�f���D��ֽ�oc���<G��j4/V]|dc�@�'dJ�+|��~A.m��g��*^��yPjzM�̊Bſ�&S-�9+��3á5���[}V�RZ�O����wd�)Y uWa�aq�������ju�[/��&O��
9��wU�W2��U�q�^{	��ۨ&ٸ�㧙����T"����O�v��T�G�Ȳ��Z`;��3.oN�wN���/��S�'0����jQ�O�]d�?z��:ۚ�%�?�	�_�ԛ�q��_X-�_�P���.k�U�w{�q.�$�VB���H�d����$3f�p���l$WJ�� Xz��*g{0*��/Np{af��H�>k���,Ge@v�W�g|z���0CyB�����Sx�����̬�^�ͣ_j��V}�!q�"cxfX�@m�w$�P����pfϛ��|���+��,M������a���J:0�BX��?�Q�z���v��� ��u��zMzN	Y���R1z�]�d��*|Kd�H�]-�I�鹭5�=׺_��6)?�oJgh�S����(����z����6��{k�Fqs�A���p�aWs���xW���i4'H��f@���YQκ��ö��\ȿ� ��$�熞��
-�0�\�5�YoͶC���V	Qk:���i �˙=[T"��+!_� �&���`�Uc���L{-;�9�W/K�9��X>Z�ÄY�G�Y��H�Z��%#'�0��;��Yb�ʃM��{�G� ��5����F�����vp�1@�U=�W%6,����	�Ig'ל
���m�v6f$�N� ��$C7$�W���0�%9��{p<u'������4ûJ��x����b�ږg�bǾ���'��i?�.VN�E�Ifå&k�Ip�]����pG��xw�\VWxa��1/g���ʚz��{�	���0�ti�a#�>�$H-%�Pk?�[f�>z(��q�r^��`�xo�*��Dy�]T���h^���Qt�����ːV���G�Qf9��Ѫ��8#�u�- �ҏNQ���E�>z�ږe�vNe	��FRfF+�P�v��]�� �G�0���=��s���z��뤉oJw��{�9c?N�$v�"��t�Ɒ���ܗ�E.b�ON£� ͫ� &tw��v:�~�W�E��K=tK�5&r]�Z%1�뮤GX�]7s�Ql��a`�YG۪P���9��F���CwY�����H�ȹ@��@�a)&T�o{8��p��<���c�����٪K��*�V�P�?���o�~伖N��U6��I��|��Y�E�'�oP3#��_r�G�o�w�\�tʣ��bH�9�O��f�=b��0!�P>u����J���J�%�\��	c&>��	���^�萸�����>�B��]���� ˠ�x�8�w��^���m
?����T���D��$.u%eǪO�,�嶡�v*���b:��璐�Y�ʊ-���;�-z�$PI���ƛ ��.��NW�On�b����P�'K���o�����+]E���W��9J��U,�����$K���@,��[�W����#��|�P�o$���I6��G��Hdd��B'r������`�+J�o��yk	"I���V�/��%O��	<IY���L��"jE,�NKn�aE�Ϭ�Н�&���Y*�%.��k�m-�߲a�/M��oX^�y�ྨ�c�=��/KT=_���{��0���P�̩ŀM^��S	;��7@ʷQץ��X�x�#?%��S3ŸZܳC������Ջ����',O*V�D�˧ד�����H�?C��e�˕mrCBn�I���秉I�zgZ�@��0�Fn�:���-*��%��j�rn�i�U�V���R�R�UXq`2�]I���Ȯ1(���n�砅����]7t��/���r.�ZV��|[�aRS�7��v�At]+:_�5�B&��Q�PZ�4�X�Л����>. k������[ĭ��U����J�۬E�ÔD
Ė_�n��S,�I�s��Cp�=p�k�ٴ�w �7x3�4�vs�a֥����;��a��8?������h0U�d��!pt;ټ
�g�PÊ�cרɤ��&c/2SmT�s�����ꛄ^��AecAJ?��/�,�X]��B���{l�
mZn?��Z��9<��ං<��@����|�㭇���^��6k�� O�������<7�uպ�����>w/��t�v����&�|���sZ��G�᮵�*��Ȯ���.+*(^�CB�X� ��<n�_�yM$6骉<qd��:�@>yv�u��Qo�b�\�w"J.�2[#kG�B�;p���}�OU�h�5w�V�},��!�s�;st�`�|r:�ˆ=
?�h�M����:��];���|���k"����a�L���/m�@�������ng�0\U�oKg� �������wooUv�b��锢1�5j�-:(G|΍�'���$|��K\@N�#�/\W�u��î�UO	E��At��H��]���?}�<��|����l��Hε�б
�Չԋ'������D�r����+��]�}F�1t��+�:hr4�ڹ�0�
ǰ�rd�Z�tă�6{	�)>V��|d�q���v���Z5p��:���+�r�1�q49���=��1S�T팯`RD��ۦ��L,�o�Wy6��HʕQ̸<��:V ;?��J�|���bT�ſ�Vv&6�e!��7�V®��L
���q8}@ K�M�.	hC��I�z(-��=�e�^���(dlP`*���[N>`�K�����Xa�Xi�db4z!jww�����;�O0�aLI
��Ï��RG��0)y��A�s?�b��7�f�ƕ�PT��ZH6������i���5��+���N�s|����� �mn����e���Щh���m&a�9A��œ"�f�ST���DW�aD|���Բ̚�a@��&�OB�JH��=a�!�hX���Eۘ��b�*;`�� �v����S����'R��"���+�Ҫ2Q0%!��Dz�k'?���o`'�!��,��U��T<P�S�U8u�J�m�����40�vGYƉ��ҁ�����zbb4P�ɷ���ْ�]Yem�����f�&~t���$�C��`N�@X�1o�:�yB��(w����i���f�r���6��ïu�X�%C:�����ۆ��w*�d_��U��Un	NJ��E`C��n:�N�6����춠>d:wP���O����(�;�v��i/p�˧�[H���@E�/H��	�H�W}̅Y�p�(d�zj���	-�jg�j/i$��@`���hIhf`����ϛ�޹(o�����Qn*�E���<[̥�~��B�8���C3�����G�V����7��#XM=`|�]��Pu��h�
�	�\"NVt�&#�p� ��:"9ZS��v�~Qg�����4n�d	V���M-�*�`󤏅���u�%Y�>� ٵ�F��I�b�i�t8_���������A/��f�ʪ��YZN%����@��[����8�ڭ)�U~�n�(��cA3m?�H{�tR=7A��E�nX|&��U6y��(a�j��/���z���8Tڅ�B}��S�*fVW�۰@�`6D�˩8=U��	��.+��^Ak�	�R�(�\x�u�P�m�1o��{�rn�ES*ʇ
�Hn���0?��v4J(pv4��65&f�{�)|	ʷ�V��(���OJiI��ڄ�q�&��C��vT` ���jM���lº,�'uv�(5M]m�)������A6g��Ǌ�cbs��I�TB0b��Z��N��d��`�
^w�l��s����M�U8�\#iz��%S�|���n�*Y�\#cj��;F>ɳ�����-Q]�@�h��$�@�AFo������@�.[@Ywf�e����Ng�7h���%؄~�?�q[���;�Ҡ�[+���p��>�!���܁���S��D��"ޯƸ�������"��4�#�c�s��7 ����{���рh����8;|�9��NO��.%b�3���Lk�����CUpEJ��~N�eJR���v�?��_ʎӉ@џ@Ʌk1!}��[#�a��o���z�������,�4����U��օ}@x�i�,T�03���P�a�-w�]X���d*��'9pi���8<��tw�&�\�
*F)<�+pӹ��}�`�����jM��	X}�&o���y?�9��\�_��H�]!�'Q�'k�J���W�דnݒG�}K��.
g񋁣XPJhd�]X�4{�n��-����yc�Eg�i!6V��I)�h[�̚K�]DƵ_*ClD�~BN1��ݎ
��l�i�0��.}��j=�q[��L�K�d���&���r��p\���6RW^���֬K�K�ugtG�=nU�;H_��2<�BNO�8��Mp���������/HqCc���}�~�K�o��N$�EcFc M�:�&�� A��}N'3��'EUm�����@\�~��*< �~���|ůCZǭ02��hŮi&ݎ�_�[q��q���Z��#Ħ�nr����=^Nql�=�cW�`��_���h�О�.���]�e�~yO`�H9��D��`�x+:�ה>7W�,��E���⫉�L8��\ϐy�*%/��_Q|��j��c��l�M�Q��1
!`B ?hA�Cm���SKE`:��|k\�)4T���G�5�Bv_�_ �V0��������U�h4��^̜Sp�RSx��t������z���j�C�c���&x��IEbP��;0���ZU�B�_J�o�%_$eɻS����X���7�.Yp�ZBĕd���}6+����o��t�X�;/(�O�%�,�<��~.�!�bt��߮߆hq:���
��tϲ��(+�`+-"��dz=.�8׬y�!�fNf�t��rrgp����*�/+�ʖ#	'�#%qI\����,�_�x�vQF?�>�kFKc���uC��y��v��/d9Qcy���y��������]ķ��Ȳ+����U�g|��jh�?L��=Tp�n�4k(+W��PM�M���� DI�/��0{��o��\nbu	��d�mU��	p�pF)��.�:Д����,b��O�PX��?	�!�>���Z�E��"2�:1��R�L�[t:	l�l9�����T��e�|m�GqX�,�W��^'�N���)�)�&N��f1	��d��\+���0���g7��O���qG���4���_���x���Z5TvX�>5o��lO��K�d�s�p��Z]��L��q�j'DP�r���rd��[����54�A�6Y�q\�+x��$�\�^s�G\a�.�&,�#���4!j/�����󌓖�[W�����a�W�� �ɝQu8�0G����p:��RI��$zoԼ�|�G:�[?\�%U~�L}�@7�ںS�Ȗ����������g��A���@֫Y�Leh��5���MS5ma�yl�o�'�t�xa���I�"��[�V����v��)�C��z?�+c�|�����k^ґo�	o _��ɭx�,�!�����Ts�a��5��z������,��ݟ�qP��w�� bрń,�I���m�,D(�B(��>=���I�2�{à�#3q5h��%����w���P�wĝ"�y%�0��L6�~Cj��pth�Q#R�Vd�����@�U��:W�hNݰ�� �M��1�-����փ����Ӣ|���,ʪ�7����=��8�~��}�p`�k�-%*����?b�`w�3$�.�$�~�v��KIF�)�%����5k��y�^W�B6��>a�}�� Q�NU/�Et2iux�YB�ѝ"e��\
�����J;��9�����wL�mP`������Հ {�R�X�5d=�'%Hm�x7�z2s�>pO���\2*f,�ed]���v	A'�[4�����O�����z�E��u~c�*�C��=�CG;�?X6p{%��P�5q��5j� ��׌/�(	��N1�ZH@���UNj�1gJ^�&��F�4���.�`�R��cUګ��SI�@�:Ǿ��g3TGȰt�.�Vm�L�]��	V��GR�L��z��{��Ͱ=ص_�nH�u�%�y�ق�� �b����Ƚ_g-��JR$�=P>���W���)���St��m��9\�����!�n��F�@Kf�͘A׆à�0:�z��RJi��*×�^2��-��p��C:�{�䗘�I-qI��we7{���ژha�@�.'���5�{{Ku�g��d���`�R$���]U�q�h��|ۡhʥ�)D1�a9#ej�C���`D[ݤ�tVG?`����F���DkEܥ�4����.)����Ѷ���{IA�G��v���6_������2b/;W@��E���|������o�G���շ󠘑��{�����ML��9T���+5����J_��O#��~�Z��l�ȹP�l#�Pn.� �x�AC����n����k7��*��ڀ��hf���J`n"��'��G��-,�Kv�K�sp�B���!�wW@+�]L;����e�KA1˶�r_t���W;�s�C�lO�/;�qO8��i�_��>9�r��#�y�^�����Ҿ)5^ή�%�J���� �y�~�	���j)Ů����j�3�1�C��k�.���E��8��侲U���k�}p"`?i�g��H���[�����~�@���zp�&]�����$�����r~���46^�]uG�絘?a���L~�#�ݺ`R�k/�O$+���$�b'�����ߺ7h��Fb�8G4@.m��Eh��D�R�&_�\O�P���v��4�#!��g����J�^�ҋz)��:�-
.��*�{�p�Rp��Hf�����VN�	ɼ9���Vz��棇An�5"������!hDc����ԇ��R��8��a���UE"���/�*��|ؿg|;α|�+5��ANp�0�Fb���JOj"�
�.AWf'*�]�n���6�~GM���>��t���p\��떇�V�#*�F҄�~�I4!7g�|�s�W��E��j1v���*D�1�Pa�҃��}�� �A����>��:�R �i&���
n�Ɔ�zQ���'��L�5��w�6��]gk�&c�Q��-���$`ǅ��#'�Q�L����ӧ5|�VB�H��� k�t	]�J�MZ'v�h�|�6���u!k�/�{/���<����a��ˡ25���9�z�d�Rz��v��%���ER\�kO��������+�cp���I��}�G�k���UJ��!ћ�@!�>��D_9]�c�njAh���{�A��v�c�zכ�d�r���R#v���� i����v��<$	� ��/�voؐ�����S���{j��s�۷X�`��n��wN�s<r���m^�Bl��lb~��=�hF������q|qY1q7+_l�$8����	���0L��y?�5�;��!n>ʼ�y���B
>�T��a�#��F��TZ0�������ڱ�?1�#�G5'%�l�e,��J�X�������"�;[P1�$hY����Ҕ1
-�,��/6:6������W��Qc�iM���N��>��g�,������j�
uQ,��/^��Q��.J��_t�q��"�T�gV'��0���K��W�H�W奔����)�1īXN�lF;�^�e�����u\��V.����4�\��n��j�i��A�9��E��_���^PERK�+�?�E0�o���U��-l��x��+�:o=;�u�?${�PH~��0�\�-y`�7�h�
7��ʻ�
5'Ҷ6AԨ�DU�Y�2���ra�1E��Z�_��7�
�#�em�BM��f�\����?�����jG����F(�f����I៣ƻv<y�[�j��uf����(��!Ė�p	}ʵ����#`�hRn�+��s�z(����
Ϭ�\~!��A�A�{�8�Jڢ'�T;����!F&eR4k{�o_�E�����͑Ñ��o�*���ɮa�邈���8�pE�QY %�GpG¶��?nX=�������:�:F�{p����a:u�=6߼��>+MAF�g1��j�oEK&��ee�d2alK�~�tBzh.m�+0��X�7�IL�jS|	⡎��f	j�5q�����F��-+��u��͞�(	Ăޑ]�j��v�O�n�\�z���K�����l�Y�-�"۸BaLf?��`sk6N�;����b�Ò؛:�e������+�p��<����b����J�y�f�uk�tfb-R������^4��C)��Q&��_I��x'K�aM!�� ����?�39\0���1�|�}ZTGW�2?���0J:�
�0�o{��P1�7��ݮ�G/��x�9�6Hȍ�dpT�Έcpl[�1NEDz��|�[��U[p�����4�O�E�V=�`gDZP����F"����E�%�j�I0��ك��ݽ�5��3K3]�z?dXD	�En����vg���xÙ�ND
}�t���ƫ����젆a��帇�	�6��0�mX�[!��(�#�
8�i�Ȓb	/h��}*q�G�̀Ts�=N�#h?7
~f��Y�sj�g_� |껊5#�=<��qŌP�$��`�[S��Nӟ�|����ր�x��y	-��b9�,���L���{�y���ׇm7���-��/Y5biљh��Ӕ)��4@���Ki+�֪��q��1�X����! Nom"�{�����ܝ��`3[]�mɴ��Y����7od��I8���|�Y��/��q���&��8�{�� ��>�'�c�t¦���aU���u��w\�::�V��}A���?>.��ŏK#
��K��á���Qc��]�Y$��.Ո�ц&�u
'��##�d�U��v�6v�FvFN{�6)�5�Ɲ[��٤/�x�5[6���@p�=tM���bڝ�8c�>����H����fy�� �u�2�?X��Jͦ��C��`�F���uu�/(�W�e��� ��o����V+{C���u�7��˶�m�xg�f%yX�\�X�{1���BNV$���Nv�P�2��֢�>Q��f�~QC�䛌g��a��[M��i/sU`��6&��X��]L$�\ 7<��I�h*C�$¦ ����J�T=��%^�6�[l�4Rh�<�'��?���6������M�޷߉��=5�&�]�/W{Hu����>���S������l媩�a����")l�:�+�	���Ô1g�q�k����31�W�5�Ji�����!��!��7&�s�8��)�1nylT-�� �[e&f�5�y�׷뽽��B�O1A��\h��E��e�t�	������T�}ծ�N=+�W\#��@}��E�V,mL�T!J��	�l���iD��i�����z�+����P���>9���G���BD�1��V�I���\9{�~�����k��Ԁ�	�F?u;���p��ұ�,�K|����}$c��&�/J ���?��~7�h���|(Y��D���l�� /DA�ȩ2uː��>(胻hѾ��0$�QA�H�a�<�4��jf)�B��rX���gY��ǝ� nh�g �Z����F�ٳ�:,���f�!��(�߉�m����Ny�;�$I�/��,�`i�8���al��_|%v��إ�6���ϋ�����L*~@�˫���7] '�=�?2%�ʫ!��1��]�&�D��#�-�Q-�P��C���'5C�H.�,���^·r����\�!��_��p5f�<)���6�=�{���E���Q�D�n�\��Xt��)�l �a�Sٜ��ե�}��C�{���(����[Mp�1�Q��ĿP�E�:�iOԞh)w�C�9/�MS��p��n��u:��"M�r��p��*��S��m����M��_��������+�r��!
��4��j"1j�ب�A#��_��DDg%GB�Z#Ŀ�������3	��6oU�>Pqz`n���"}�7������&�]q|b�;sDs��� n,._���p3�H}�q��b߻�Q]A��#SF�$���~y�UiR��P��Up~Mw���V��wv;.��Ժ�{�e�W*�e�"�AW���9�վ�
+�� �H��T-^��@�t�F�B�@=�k�SO�JJ��|Ԃr����J'�RB^��r1�:ki8bs(�n���B9�R`��י�P�(��M��<��Y�c:�B�K����F����ɫ6�C�M�W������~T-ϯF|q�(P@2�b���4ϕ��.EcZD�qjڎ �N�h;p�!�vC$�#��Kv�XA�"6����h�?^䊟JɌ�jR��@sT�;M�E�#�VX�zx�n\��������2��5b��[U\V���=�@N�؟�|�-�p���Zc	+|��n���Y��9�1��}N�J:$W��Nkq<Ӱ|�Y/Ɉͅ-!:���{���Ө� �m3UIj�];:"��\<���X�˰G]�u� �����:i6�'z��>�̽�n�+��b�S�^=������:e0B�u|?��g��ŷ���W[��!��VSh�&�>����e�;��F'f��IRy���y͠�)���{���w��B�	��h�v��o���	�q�v��}H��zQBϛ�!G�I!nDTPJI+Z���ޝ�
��#�$�[�pٞ|�zR�*&�>k<�uy}�1���3�'��E�(��@{�Í�85�ٺXbM��f�#^��;���W���
im*A�+u��6n�!�����W���Cc�t���ew���yQH�7��v�ɩŲP8_���7y����,mű��o[ x%�" �	�^�o(�|�B����'2����7�QY��d��h��O���b~�N�Nq��#�ڲmD�X�㘶Y�:�t��Ђ�mr1�بB��w�%�]�s���L�w����ˏG�d�Ě�H`��=��: _@���>�VX�N�OjЎv�Ӧ�X���?ĳ�`� ��M����H�C��zM:�\/|���t�o0�h���v�93Z�Ug��� ���4r�����}����!3M�<;�:�q�A9D�s��tڮ�P���y�w��3N��_u��8���5r��)02�U�8B_\%1M	&1�*��O������'�Ֆ���}�i򭘓qI��d�]�}��h���q��Z�3*�B�������ɘ�ϴ/�$s;��Hk��!���K��	N�qC΍��P�rԁ��U���BKo^���6	q��~߯3������3�	#_6߱*R�K�Hk�+�S)��s�JOX*�[��IJ3J�2�"0+O_?���g,�Z'�*��r;R.M�twы(�L���W�	_ C=��j8"㠈W���x�G�V	>o7�
:�¦x����qB!R�o��� �W?���[w�(�@�&�q!�ډU
c;� ]�t�:�{��2@=��DB8>��g�s������Gv���&���ޥ�0��d��2}�i��*�b�<I�Ԇ�:�ON��.���.���غ�ōv5�u[�ܢ�������w	���vgq���X�Zyd�Uv��|@{�Tg��]k3L+�#J�E�� a�N]7fxm$��a�tq5�_}?�^`X��ZHx����0�}�t��	�<�H��z��%%�Y	*�����2�2���o熯��q���U��)F����-7��B�pOFYuh״T�ï�МLם܎���<^R�3��fB@t�z�"�l�6��Y�!��y���(7tq�[�!{�9V ���	�C'z�D��-D�?�C%�T�Zs3ąN�Sn������/s�q8��<Bz��U�eA�(����[O��k�BF
E��Nh�_�/U�ؽ�>��V?RY�+G���D2�ʀ������e��k����T�Ci��
��~��"�����f�t i���1��{FЕZ�a�G�	-�0lI�)nE��Kz>߅'����xD��3�����u��I�߳U�@���ڷ��fL����[�~[IRm�$��X�-�ILj��Ӆ��G�~W�>�G��(��K�6�q��R���?�`��<���_hǛ�hy����Ԇ�z��Qi5V	���Z��B(�h��)$!-�����Ơ�l�qU-�\Ȳ��ރW�:]r���i:��F�ܥ�W��PVO��iCm���Ix�i�)�J������ �TP' 	���=��C��^�Z���բR|�⛖ǻ^Rٷ6##QEH��g	^�ڮa͔a�{Z�]���	�W ��1�*�֯��U�}�%4]�	z���������#��m4|��MU��� J���h�3������W�q{jT8Xs`6��0���$���>�z�TʩT���\���+'�,���%W-=@�ޯ�qQ��Zh��UϼK�v	8�ޕ'�O�e^����4�Ԋߔ5�S�����Ch>ȼ�����yW��<��f�o󯤢$'B��"f*~/���!����a;|�zĺ�E�tl���!�6���B`�~Q��*�?��~Ҵ��p��j/|��w8��q�j~�_�Խă���lͤ~j�>�qh�Ot��5{��η��#>�<?/��]}vk���5r�n�)K�G��UQr�S�k��kd�f�{bS����uΞ�vI���MT86=Eb�yT�7*Lx+k��/�m�����z*��g��Pw�M�ف �T�h̤�9K4'��x^w}�m��g�2��r�\O�]�'�X�����|{�F�AǷ#�ߛQp,m��Kۤ�L��8�d�e{%ћX��/!
���T��ym��++�wn�H�z����J�T��?VA��ثe�T��wr(@�x(;�U�N�EǊ`�V-$�/R�ɝP6N鶣'�$��MTYK`#�$g��LG��v�;j�`m������tLU���4+}��>ߒw(x�"7����Gڑ.��_����:�? ����d�0;X!�sh�hc��l4�ư��#�W5,��/Y��ˢ*����Mļ�+�_y��fkQ�rf��iq�h��]�Z}lm [A;PZӸ�J}^��'�B���??+�M��1�2�dt7k�jT��Ў�cb���YR���Rk5P�f�n�CY��r���<th�Q�+���٣l�������p}�n������}���P�*�W5��haju�i�~�-��N��ƏL�"����$��t��Q%׫��;�;w��P��)��i���Q�_�!,�����ݽ��I$N��<ZJ�-/k�붷��l�fR-�A���U�;
+
�ڟ��L=�%�I�1{
��*�¥�J��8)R	`�{%��)I�#�ė�)Yѩ���V�B��L%<�'G3c̭�v��M�g񶷔PQ�U|Pӗ��%�f�U8�>��������	9��B+|z�-LHn>_����z��<7;��)�2��Kr�]H�[6�}�2��S9�ר�[a��0�	�d�#)�\X���������1�v�#��S����-�<}�E�;�u�=kpJ�ڑձ��h�����r�y���9�a{��-��U�>��r8���ډ�^�7��AF���E͘� ���@�\(P�/޶)J-��m��yA��=mbM!��#0�@��p�.<}�>�ív�0�۫�6��S�k];�=�� NO�b/X����'�{Y���B��1��t�N�{L��p���}f�)1E@a��H]o�������BԐr>����_�8PU��������O�[�2T����N��$d�7�5?����k�U�W݊�61~�$�?�@�%�}(�+���d9�T��c[�t���,NO�1��*��a�,	��7��k�UU��Ӟ'�B��dP���f�5'=]��E�&�N%��]] �V4ܸ
cЉ-l�{���&U��t�(���~�b����Z ���;2�܍:������٪4-c�����6�C@}df]�PR�����p�ǌ��\�V����lCP8T,��3i����h�L�Vm��P+!��OQ����	��c4����m���}5���'��^J,��K��0�9�l����<�s��bEc0L6��f�՞��t�)e�o����ѝ�^�A�r�n`Ls��n���̮/��b+���v��2���7��ZD
�"�X]t����R����>q[i���]������I���+N%���Ԭ"(+�Z%\mS��g3Sc��q� D��$.Y�n��"v��G]A`F��T����aE;o��#o���l��'3R����%nn����Oׄ~��&(�rRD��I1������Hu?�;A���ldO'wX�&7�z���_`��-�S[�v��GW���1�ȁ���iB�����Y�˶��o<�SGs�`�/�g���|���{�8�2��H�$B
Ƥ	?�mN��BE6`��չ�yǫ���rD*u�hϓ��-Pd"6��尲���@�]�������J�,?z>�o�)*;/X�՜KXXǄ�;�Jd�j�M�R, j�LǮFXK, _�aufpo*�zQ�>��v}! �v���>=����XU���5��(Pv4k��"}t�[���l���>��Ӌ6T�i����0�&�1^\6��:��^��{��*��1�D���Ktvv�/�7�i�~8��LZ����{�Im�׺�ԯ[!$�p���k��6aG���Gޣ���p#,)Y�!��"zV�RC\C|.lP�l�J��!�>��+��l?wӸVeO��?�b5��c�6DB�&�����͵����?��
��hV��$���˨3�L:U�P=��I[���}�y보}�38�-��3��"-׊Q�Y_��c����`Q��������̦s)$սBr��ϟ<l�tUU+*�ӪtY)�0�c��p��t��38|�G2��>�wd�4�L�R��h8j��d���Vj���Jz#�'�l�Օ��3�ƌ�T�s��)9�R�k4-��L�~�m��O�K~��m%��u����8ۊ3�����L���&��$(���]��M6�Y�7�F/:Fk�wW�,�����5l�Dz}��_�<pD�c�g����V��'�᠎|O�1�8�a6�����~Xr�.?����І-��F���� �E(�!-��h8�63��ZN�}���i ��Y��0���HGb�G)=ǈи蓬����8��";�nۘ{s�4_�5�����H���Y�_��3nS t�����Ζ�2_h����xb������-����^�Ҁ�9y�QqD�!�"g2O��K���Z��mc�3D�^�'���`2E9���+�q#�]\���Z������s�s��W�7�	�;����m�ч �h�*U��F5�-���O�e��vnPS�vgPl�B{��ʳ��̌�K���s$�li��/ʭG�=�M�аct��.$���:��w��:���/��T?;���l�g��`��P��vs�
����̼�/���T:���7#�nDv?$!�P։�(�FL�^�ܐo&M��
��;�tL�k�,�� z����/f��	��`����fB�N^����_��5J��u�D���L�����|�%����{� ʆ��!���&v@P5��GAN��E��<z4!��E9%^�t����`��Y�F�Ұ��V��L�W�hn��H`x޹��p	[]�rM���q�>Q��ʝ�A֯�?�����FZ��p\�
V�����H���؝�4�Ik�Y����_�k���6�*����X��D��nMKs�5Z~5R�����<W�'ˌX==$�r5��
ƍ/�h���R��k��RC����S���~��ɾ^Edn����`e>g�(}vS�2��
H��ƝL�A5I&�#g ��W�\:���6��)��e���ڞY�W����TH.���VD�l�oU��*����h{��\�k�c���M ��T\���"PỮ�on)l�7r^J��]�#N%Fj�u�u��i�D���ˠ��~%��%� 	��p��-�!Й�Y-�G��7LUZ�j.���O�P¼WZ�,a$o���guy�z�����H`p��}�X���P�f�Y�J|CTl���\��71���
hbCjV�8��� �V���&��tq@`[�v��Hu#�1  Ni��� #>]W��z̪}�\9��J��w�&�w#�e�o��-h�0S .��'r�|Y��	N��N��� ��n�\�����J�0�{m�-ֈ�Q~�iN�2�.�`ñ�<�Xd�C��i-���چT3g���Z��7��ɬk�qu�٘(�+* Ugi�Gj��ԣ�1����e�Cl�KOM7���Kz��.���k�޽�V0��%gNNK�_�A��h�ST���i�@�pA��xF��ؔ^:�ݬ<��ka.1%�|�nm�/.��l;�A�1��ݟI�0c�ۑ��x��C4Z�gW��{��)���u���}7�O���;�e�)���Z��N�4,L��;t]�c�H�����WrE��$�9LN�=I����!l��h�Z8-�,�p���WL�[ܡ��جe��|�f@�`BG/�� ��ظ�.t���4~�lޘK���By
.qr���#��L�|�m�-W�%&�KkjXj�8��ف%�R?���`kf�sɡ��Go8�Q��GGG?#�D?&��Ə�F,��U����}Y�3�[���r��2k	f��4���Pf��2�?¾�U_����Bʂ�_dW�q�hx	�U��,�K%
M�9�����{h�Y���\\�S�"�#�P��\T1���
�ȳtc&��u��ZS"~�Գan�d�~(��6�h�l,4��+� ���(#w�G�~�
�{�i��h��?��D�#� �Ӥ�?j�+�w���U ���V�#��Է��cz���KY�V߬��5��qF��N1���r(��<�н�)�������ji�8V����TC�F���y��t7Pp��v�-���UJ�5a�[{ͧ�D��-�D���t�6N���֑*�n�L�{J��x����B��4�v�T(�ȆGY]o8�!2�`���e�6�ú�3�螒]�B�N�+x��t�7@��ԃˮ�wY@ޕ�*+�����<���/*XOF�(_WZ��u��E4)�%D�����B��N�R�.��~��Єt�&AEk�ٮ(y'ˉ��"��ӡ�/A�.�K�,FS�UAg����go��D^Y�y����;�Z�݌�"/�|�f��c���Y�5=%���,]�ll,�"˲^��D��]�&���%�\Sj�Բi�Lª�b�����ɏb����4�ʦ�=Ic��.%2�s�f��]�7M�R���q����I��� X���t�0eTAu.�ÏG7�t�HHBt{�e =�'�dcΜ�z#pũ�Ov�� /�Xh.h��<
'�Ȩ	�%;,\��E4��P�K�'=$�~-�[����{}_�ښ���i�Q�N3-iQ2NQ�F�.���B�#�j`u3�Q�W$k��C �&�vL	��ē�ֽet�_pD�N��A_==_Qz&��p����b��^������t���ηfSm�����$B	�U&�^]�@+�킳`������s<D?2Q}��Q^��(ڄ���f��Z�4q��9����4�
Q�e�p�.�����V�O�1��Vߗ����&�� �3pGM��2�s��V>���I�AB�\	VS��zuAtY�5��cx��a�.ZU��7Z�
�c	n7��k���:\�hb���|���JH|���Uۃ?{���vQo�����ÿu�A(��S���]~�33��d����.w�P�D���3Z"p #�=���,Ͳ�y
�z��^c�}@��km^v~J�q�(�a=#V��N�W����"��1͎DБ��93Ĉ+��i�_6�0L���[�h�
2FT���Z�W�Z���x��LE�Ӟ��F���}�|B��Z��vo 02)�]�K1��j�q�~�ʁM<Wa2�s��S#�	`��"]Ag��E+�P��ב���H�Jd�=�)�
Pc��	��tHv���=�v-|.tc�w-k2ů�	�w*\����8�mY��L]Nh"���HBp	��[�ۈfL����Q8�k,r1[	�]����������J�Sz��%a�5ŝ`�/4!,��5̺$~/�Sʈ'�e%�3Z� oXR_:�ٗ�h�� ��	+�'�Ξ�e->˔%���Jr�����'9�c!��^.c�f�
�\Rb������)e����X!	�|1t��GxV���'"9 �ϒ)��
G<,(RM�C���fg(�n��m�§x@W��VS�H�{��}f#v� k�`��¬i��?����� }[����چ��ضX�KDF���d��� ����AwQ�-x��֔\E� Z/`�[r��D��>����?�Şy��}�,��mċH��9ht���m�^�0�J����כ��=FmТ	!6(��8�\f�ju�Fed������G:H�'o��������x;�PWO��gd�7�`��2B_(` �Թ�Zk�B{�BL@+���8��4���qZT�tD{��8P=���O�j��;Bf��C�9|4�t��T�.c$8"84l�#S�{�A#�mP����lԜe�X��S �j�x��Ō���s|��A��!��*���'�c��L��Bso M|0�cjz/�������M~hy��2��w�@Z��;�t�#$�i���(^�����2��D��-��N�8��p%o��*oF����I`�R�;A�z���)[�o�HJ���(��^^���wo��G��#���ɵ��Y�ħҨ�AĂ�t�M+R�����W�Q�O>�NG�*.ʾ`�V/w>� m�5$������aO��:w�����=܇�ܟ���mA�8�(��ȟ�x�e�$�"�b���G�5e��`����P�;�f:8Ŏ�z>˒AH��V������\X��󙨱�(���P")NM��� G �[�5=+9�Ηp��)	��svx�z1��t��|ٺي��-�mL�KW�u�"��r}�d�����OÕ��g���	����'¢3���k�'Qq��:b
糤���F�����B���ϕ8��2�c.�p]Cr�!߮,�d�.r�^�;��^���Β΂p�'���?c���Ƒ-��6[��AWy�%\��+�|u�LQ(��4?q�l;��=;�)5��q@:�m �����o����II�Ө`�I�=���d���!&�TPY�Ii!,��el�z&�9�����u���=�����#�,S���:��@��{V1�����`�iL�0`_� u��-�os+W�KȲ�O[B�Aj���C�v#qm)T���͆dP��#N���)5�=��2�,%��뗄�'X;����"��T���R��D�Y�k92��AL���j����+�9sו���rHde��B"����%	y-�x9���&0Sd��_�䦊8��@4��מ���%�"��/;�~~�o!*q��D計���McY*�Ͼ���?/n6�,·@RnS��O}1�A��~z���%C������z�`���?	4ݙ�E�`��\Z-A�郯&K�5�ቜ����c�jM�誅�$��G3g�hUڀ�~V�V�؝�=�6G�
� ^u?a>%Z��G^�[���
lk�_��fz3w�U���k.u�_$6#�m!�ehw�H�p�]ZK=��v�+���.�nX�19�Y$�J2U17g�;�k���L��~�u�jTk�g�!_I�jY���r�J��h�(�^8�_L5�iY+�Ʈ�O{�����N�� C�ߏ;�u����Ύ�kO8^pUw��ڢ�ۓ��)s��6���7郅�#�z�͇�H�i���k��؀���1x�,$,d��niN8����D��vU���)ބ��<7N�D(aW���}V�#�f�+��-e�@�]�_S`%ǻ�����;:J^�H��>��	1����Lq<����q��k�DB�v<̴��p�.�x�[���5��ji��v_d�-�_Q ��[;xk7��K�7�u����֛-҆J*ȵn8�C�넑i_2�Xrm�\�a�6�FSI�Ļ�J&��]���MaCux�0��. "�)j_�����N�ľ�e�,�Ո�P�p��;�O�[�m\��O�hA(X�-ǪD �{/��|f�d*T֑��	����l���/���k��QMt�l�"��?��'���Z(*����ul�a�� <��D��!�c�
�eT���hw�y�iw�bI���A���
K)]�`S<��c6�mR��=L�؜n��3].���&�ں��B�F
XSJ��d���-�)ؕ�+;:�_YӁ]
��;"78�5c(K�J���`7VStV9fV��Ok����b`;�|(�=*vO#��|m}�]���tܑ�؀���e�,AQ�|ƌc$�>�S+��O�Ř<a���8���o�=�n�t
t�M[o3���_��t�~�z����+�B�=����ss��{�W�	�N_�F���\��7��C��ʅ�xscge���0��Z��9j��@P!`R\�a�3�	��,O=y��K����E���§�˟܎�!V{��Og��Y�-�����Vsqx�9(��.��^K�Z>w�0]�%��[�y=�����z�Y9�|�h7+�4�������:��@4��#���D^��a�Hb���hi�ޓl��#cD ����(�H� @�+�S�E�7ŌZGT9���\�"jSF!�Ǖ�>̗���ϚX�m��vaK=�OR#�쐫(��˾x�<����ͪ���bV9v�!���С�|�G�w��X+� ���4K��׺����\�u�:O���@�"�ο�@cU+���������Z�Ni�1�pmG,�����(�}Ы'Jx�6�ǁ�U�F���=@ �f��0
S�W��Eq�~5�-%�����{�P��>� ܬ@1�ut��+׫� �;���O�\��F5�����ښ"�/�d^ 7�ֳ=KcU�ۀ[(u�:���{����Q �!�Sp����+�	�>{���'l����&q>'���5�C"�?Q8����%�]=,
�iM��|��}�2��R��&�ZR�kW�<n�?{'��ĩ%�<���� O�VL���<۴t��i+�
�Z}e�-y
���Y7��W��3!3��v�<#N�/�K�4��H[E���4����Sr!5Y�e~?zd=3hm�m���[~1J!������]FXD@ˎ��O$�ʜ�B���r��V�#��aD��d�g66~�s���=/e��v��G��(a0��v%"�K���'-�WX���B�7Sl��{0����F�!��3]�����\��\�[�vg�*Ս���$*���黣ݴ�������!�D+����f�1W\S,
i�=*����h�1`�hnXj�f�v��rL^|��p{=r�2�\_M|#[=#�@����U=M�n�W�=�Ӧ��C�u�z��C>�A�J�x�{�"5������:����X�o�Ζ����:���6g�\�Y}�C(1T
��`'�|�DZn}��1\�LC��fu愉,���@c�����]4���g��Ä�y/�g[.�ZZ��x����D�B��Ev��6�g:���rw�@�(��A\GM��m!ܗD I�����2�R��=p[�1U���gJ�WX�B��E�"L���e���6$P�씤�g1@b�3�U2����b���k��XX�����ڙ��X�B�)xK�������!���l� u��L�����07�.?0N,��2jG\�fu�m� 谖.��p7�wպO��+�;l/Q��o^�w'�䠓�չM��ɯ�~�a6�ޏ�QG^X3]���4�J���C�8���������=7�7v#�?z.�p˅��2F��UL�5�g��������Ǯ�?.�k2����֜�_d�@�/p��Bk��s�|mN��L��ע� ��-�I�=$f
�)Y��r(�_���i>U*L�:�(�91�[�E���4�II�%EY�L��j���tg�縉�UA琦mp���v�r���v�M��?�]���p�HN�U�Jha�*W�T�p܍-�cY�XfK����>T>�-8och�8p$�����p1��PH�G�Wp��x���̛;��o�ޅ��/Mʽ|D�ЏY ���.	<)Y�2������(WcϩRId��j��+\C���f�'�A�w���u�H�3�Á�nU�H��z�Zn<��٬�D����,Wd���I�%�k�#cC���� C��G_E�H³��A#�2�5k�]\`�4I�/�#*	��|�/F$',���:���<�]�Cp�@�D��b��i�O0��q�s�K��6^�`�cnQ��`EP;>̅�:��5��MS��7J�sU�%ל�'a���8_L��:�#����QsA9DD}�>��1(8s8��g %��ݰX���/� i]w	p�h���gOE�e�:�1�Q�R�^OFI[�l�B�B]�,�Һd�D����V/I��rR��I.�'�4ȨܵB����uR��;�ޮ�,Z)'���)�G���H�����lM�6)�u�%�M���A�.��&���i�,��3�"Q>m&����k�Pzt�w�(��V�하+_NE��ݕ���u�e�|�톯5#J��1B3K�iOM. A�x�2<�mU+D�:���\�h�^<����6�q�'��z���W4R�*|��ʘ��<𳾰��6��cC�<����e(��2��3}�1t�\�D9DQ��ӽ��-r�,��c��d�|G0xu}�l4�"���B���� 舄(�Ӗ�pH:����F�;���<Z��������L�1
~��&{l(1.����g��FQ���1k���2���x�����"�����M$�$�Zojq��!�j��n�-LNrs[�ݛ��\�R����z�V�iRB"�S�Nr�^���$�KՂ��=I���3_�L<R����jZ5*�i�Ƙs�3�g��"L��v��z��̀j8���mp%�����*D����'4c���}3xߝ�����DD�zt=�� SJ�|��A�J�^^�L��8YO���J��E���zV�
�=k�-1vJ��B���"� ����;����~0}�km�`}�A��;`A�5��ـ�'�ʺH����q�Y5���f:������=���EIY7Q�s'Ci'�O�.�ļ-=��˕Y�p��X8�PɤN�#�^fe�1��zu(��*�R���}_wN�R�/�ޚ��Q��Ĺ��'�<T�}QS�����@2Dd_�J����jx��7ķU�r�����jg)���dAT�wYd�;�����4TZS#�� ��i����q�r��(\���飧���,�F��[��-��%��	�>l�6���L�^%�^�Q��G�e̸��'�_��P
�b3#I�j��akq��5�MZy�[�ƕ�6����rB�M]Nr��!���Ē�{���6*�F��_��Ї=q�%{��`3vl��1.����؉���y��_1�3����K�*�����Y����O=is�d�i1G�֨�5��3���Hh���uA�i]��c\a������-Ә�L����A�5�\���o���pq3��<m�!k�u7�(�����.��nyi���<QTK?���MA�gX��z�Z-����ڹ����>��(B�*�:�A`�x`-h���Z�1�pa���0��>� 9T�b���d۫E �Q(�%=�S��0���k�'�MSl6-�ŉ�t�:�8�ONnu�����������	��(@�)�����W�F3����s��v�����s�ĩq_}h���:�0 ��$ �TrZ��P������I�}p���Sm>|��}
�U������w�I�ї%�d�Cx$�A��b�/u�?j��Rj-ʖY��V�:/~e�u�Pxa�ĥw'�������/�{c����\Wh�į��8��@'V�F^'TӻTM䶏Y<g#���=�=����':1�����7,��o ߶�V��9n�U�c����x ��J/�%иҒt�]#�%=^�px���s�S},M$���J/r�=y�hUN��r�'kN����&SΣ����䪐ӹZ+���p5�u�ؚU�� �Æ�8Х��M���{��S,~�	Z����鵰xLmE�g���=L
�eX�������hmMM��=q~`����]��Ѳ�Ɵr-�(cf���^�;���ɺ]����=r8�O]���3A�-::���q nga� II��� ���7�I�����2/��<������8ɨ�;�ݾ��A e����*�)�[C��{�АM��o(�� ��C9���Bi�WH���;��gl�	;3�U&�mX�_(����jm��kq�R�� ٝkjѧrj3W��)^pbx.\�}�*���t�a�Je�Q�؛���2�$��@��0vM_z/���R���T�CX}l2:7��/~j���p�g5�g��<C��R��F�f�j�'� "m�0�x�0�b�s ���l��혇�=�s.P�4�z��K��%�j���m:8�6��T9!I��[��G���k2�|JsZ�J�v�1:Tyh����1ه�����y���ҷ�7� �/Z�}��w��j��ńw@J+A�F�dُ�~5[������#�sݞ)�&�
Ϙ���o(���c�`S�����r!ӫKgTP/_�rCa�7�*UKۀ\�ڟɠ�Jr�z-��w|�<�pbwc�tb��/�X>E������4bqu"da̭�_3�}��Af�̢��^��l��{1��5>~�.|ڈ�b\��_g!R0�)�!I����Gۘ�i<{�b�*��WX��[q{�Z�M���M�^��E�W�7�V���$���}Q�Lu���R�s�i|}�G�䲴P�)�qv$֦��<T"�_��gW��,���u�������"��-��䛩A�&�� �~}Ϣ��/6�>	�)��r���+�\�;�:tz�aW��]v*(�O��Sl{��GJ���0Y��(:֤7o�}ݖ#2��g�i���?��_M����P9-���ªa��i���GВpf,EĤ�U���6k]� ����g��Z-�l�e�(��=F&6
`ÎR4��Y�����#�̳�j��l��F�~���ח����ڤ�����/�%�bT&���<	aѬl<�1Y����7�����,ؘ�I�<��8]&�G�]�y#N<�}8�%�E�����2�=�q�}�ۥ���-���`н^���6
����G�D&DJ
6�;�䢟3��O�?4 �7L/<a~��Bx�ϕ-�S8H�IR��O��k^y����8�I�	n��/!̲�5T0�9����dr������ONDq'�f��}�4"��n�����VZ8h��o�Z���
%�Ԑ�,YF���4�'�Y
��_�|s�8�	-�߂���wh�3aS�����������sR�~�}zu��]�a�v����J���R^v�"I�7нR|jN�sW�n��oiVB S�{G��5�T��A�Г��T"��Ӽ_'fE3��#w� ��wM����OO�r˜
��]�S���3Q	�*��]�|��"������A��������,�u+���S���V��  ��Y�t0��}�e	��k|Y���<[ghC�a"�ͳ�����V�ش�9X�����be��h+4���F��x�dOQ�U��&LL�}��Y������\5N_�G����e��ͭ4�x��w�:�$����.��7��+��������6US��<O��/u�]�{I�<���pP9#a!�=�lnh�<���h��r��8{�{�5�d��tF��>4O�@�B><�(p�#�'�k�%Mk�PG[�ǣ�{�̪� ;����cL�fЄg�@���g�5��E�3��N�����Sҩ Zo��n�쿴�7��E4k� �/�ب��F5�JM�45.q���{��CM<�q���t���!0�O3�9N ��+��1���hCR�Uɷɵ\�]7n�FS��HH�F_xw���9��76�e��0��~�9ĉ����S��$C���v{�o@�A���� ��v�2��<�������b8�m���Z�6zc�w?�z�s�%+�� P�w�i��l�ɸf0�A�|܉Ooک��r�%p��w���I��]�М�Fެ�NxD�CW�N@�A�)�Rv�Ad�F�TBnR�'Z�憷�h��n!TV���^4w���yp�Sm����A�$T���Z��d
�����[O��<f��!'$e�T�CA���|�F�I�1ph�V
��d���a&�u�>'���Xױ�'��))����]+w
:���I;�"�_b�,�S)�ր%�6t����4��^�Q�uz
��Q�@~J���Z�N %P���q���cq�c7߹�0�]��E��y�M����虗.j�E�ﹴ�܂�@�>����g�Y 4�~�p����O�k`B�ғ�{�
K��0���*�[�>��%��qp�B�a�Y�����BO�{X:d}d����z�L�Y�?��q�v�']h�f�#�}b*ι{�5�p�$�Rق#�=]���F��+�ƕ�J+d���ۭ�%7omx�э0S�0 �|��"�+D�L�kL±�x��;f�����Kލ_��[aC#�k�syx��6�m�2���i*�W� ����--��(�!Nc�FE�h�<��,�Wm�`��ԗ���S��:�nZo��h����c�� �l%�a��Q��*���˙hw��a@lRAom��L�r�?W>d=&�a-Gj�^fcFPh5U(��?�|�Z#@��M�	$f\k R���]5����M��<�Iu���d�2g-9�Ј�'/#��q.�/@�8���� �.��p�iL��h�〰�9�2sπ��	�� qrx�N�e��L�v�#v��2Dj���I:�<~���.> wf@��MC���?q,nZ��9}F3Ǉ��߫�$L�XS�E��|��fq��rC)� ���^�À����GJq8JԤtl���r�t����t���-9���k��7�%&jyb�o�_ ��[�"�az�~1�|�9��K�8[����TJ��P����x��!���
�l�1�`�\�R[�ԙi�O<D(y8�r_tU�W�߾>��c��Vf�ڑP�OYH(�C�+]�	�=�CA�Q���������c��u�ad��U�8��i�Hk�#u(�}��Zn�iL�bFΗ��Y"��`�N��{�N�8������%�+���0�/#V���|8h�D``{��CQ�� r��z
&/If��z�M%a��X�����
x��G��r�f4�¸h:�v��ͤ���oI�J�&_%��(�,J�7<��*[S��{g�{�{���:�&nm��)��o9��D^1��y���� �]�o��]�\���X�3��3���Xi�My.ӫ/�-萖�B��yk�%�3�$+`�tH�b,��[��(=��&��	��� ����,�+Z��Yǋ�Ȋ�e�2!�Dg�U*��kN=Ňi���~�w�SSPG��}�W���I��ˌ�����I�_���8:��r6�|[jk�2��3������h��,E���I�Kr�٘@���3^2��zʎ�]q�h�� �����x���=�i�4A���{JOd�p@ǱG�G�m!ѧ(�f�w��n����K �X����,!U��9���Ѻi�b����hKD^i\�1���Q�4��Y���q#q���j+n 4Ԡ��n/>M�SI��	�֔kfn�<j���?��B t�������xz�?;7�/��
�>���8=�'� .���~��Ƥ�q�j�U�^Yѡ*���.e���"����9����O�`��,Z��)l" !O,g?��w�k7	�K>CtC?9	;�ǒ�E*�YB�V���$���0^c�8�$ψC�J��K�3����1*}�!�-o(HH��E��Y|�Jj�0��(^����O[Zϕ�+5FfT&�җ�*r�A��Z` ;A��Djf`�0i^a�Dzx.Hn��q�X�M�Z���vp"K�#�Qy�6��.ŖGf�ˋk4I��!��(\E����?���{L�l�ʬ$C4a�C�o7?qo+�J|��Ը��?��,�9�?z,x�;慩)�������?|g�?:�<�wy5*�~A���n#����j�M�c�e�@�)�K��[XylEB�ˏb?��	��9�?˯��zdH�(r͖kL��.�z��a�G4�a�i���:����+��u@�F���
UG.aa�5���Ij���,��?�����$Z��ߗ��4g���G�Vd�
Z��w��3(�A����X>)*�:To#!���� ;m'��A0�o�d�T>�*�,mN/ax�C5�@�V�,}�4k�wǮT0K���&�ǫp;�l��uY5��:��c1�3������O ��|��eަ��
݂ڢ�\�hRPr?r� l��Z�Ӝb˪]BQ�a��w�h:*��]X�x�@��V|2�<����aO�)��3���}ɯ�Ji�6��YR�}�:z�g���:��Ȼ'[?|3c�dMX]2:)�ȹ�K�;���u��|"��cOȋ����,�W�j�y��_�����43� �I���g�%Qt�ݟ$>�_�'.�R�Y)2ɜ��2�k��a`1��	��gBs?n��\*K�ߩ�<�+�I��l5�7s��9�l�"g�!P�?TG����F/�󷾌r=�!.��g�:����*��s8L�Pz�����2Y`@Xq�B]S��k�QϤ�S@�ⷉ.�B�;P[<�J�z����k�Rpԯ؉�K�\b ����8F�O
�����fd��Ğ�c_:-i� D8�<�����H@�Z�K[�d;�&�[�z��GJo<��*S�jg�B棊�lN�U������i�T�x:=H�]��f%� �Y�?��>�(��5�b�u���XL����<��w�#
ʘ�q�p� A��A�"���z�p	�a�����7g�k�~q�|��La܅<$Zݦ+�]�v�T( h�7���Dm�%�VjЈ4-o����tE��<p���}�2����b�lc��4z�=�c\��۟	�+���o�K��Ըu�k-��+;,�=�x��?�����W����@��f����h
�	�
��o�jn��ZqKYX�e�f�s	3!8�OF�9Xa��0��@c��ٵ���|H!;�`S�LJR"6ǖ��,�a�?U>��d���n�Vء�!#��kw��1���"�3�1�%�!.���	q3��t
����f�H���o��������O�p�
4��MM�-�d_�G����y�gH%Xwl#"@L�����7����zQ,*<�����y:M���
�=yS��: ����p䘪���t��kX'� ^��i�^���c%g��eR�rӄ�AQysj�0B�����I��GWg�625���3��I�(�mJhl/WO�= 4��U쀇Z��]�{�s�+��V��;�P�5P"��w�m�����lHH�hk��Y"��Ȅ?(6b��֌��ħ�IM����d�-�:5TМX�a���h�Ɓ����_61�r�_]�����S��.IϚ"(�=}Q3��IɋLk/1=T����B 1��ɣ#�cN���6ՠ|o�H��A��v�Zު�?�`���_��֣�A�g}M/7���v��4�E��l�ȧ��9��.��{M8�&:<�_�7坌��6����Yްq9 V�v`�(��N7��;�,aWr-͜N}�կd�<i)CЛE��<~���2>���e�gNt��i9��I�8O��l{'��(,�MeE|NG01A�� �μ2��%�G/�k��\�C�9�ʹ%�]ۋ7���4���* TU*\;1�:6L����+W��bo+m:�M�Fn�{�4F�bR��[H��j��K��9���Bɲ�ˤ���h�K�"yKH�\1�Q��u����T�eS��\�l�{ܽ$��C�Mjۇ�}�c���P���X�<���QwjO0wj�rep��,��O�>]� �2'Ǿ�Y��o$���z���؍����{p¨J0�Nֻ��^	���<����U�w��s������V.]�-Q�F[�2:G��ǜ�����EY_dY�Q��վ3��*u����m�]��!G���\��[�Q1e���ng>�v3A_��C���7�E9��-����Sq���	��.��,߰���X���=��Lp؂>2�UW�:$l2l�f��#9�37�'�UD4?��* ��H(���Yu���
����{�r8��j�~�L�]E����·�������*m_*Q�LvQ�a�]P�I���qvT�^
Z3۷\����{�۵i�Q�T�A�á��Q�-�7�j��Zt����\������ u�+U��aE�룠z�ơ�t�q5R�`VQ�Ң�K@l��҃�\k�hj#L�R�*�Ng���|����~GyT�C6����6���w���̂����ͪ�����k�F�)J#�J�q��mu(��C���	���c5��+�6����]�#wQ��{�ͯ?�^�5i��_�:�G,=W�q�HX�`%�tf{�1�w��1oУ���|���{6�`�{o~��3,rK��˷�fKlE��y81H� �*W��I����3Λ�i@��� ��ؠ�^a��B��~�I�tBP�3�딞�j���;�ldx;@�n9m+j>ٽ ��Y��<�c��q�	RQ�[���_����j��t
��@�@_����c���7#u��a���:�k��`�
9��N�Qe����,��-���{���s�
�4&�>���(�E�����^��؟�-ÈUTT����w�8��&e�P�LZ- �'N�h���ǜ�b?uH_M�!�CY���)�3�l���ޟ:I�j zG
|���㯵4�-�"��V�^0jp�iWAK�(�S�h�[�S	'
2�ޒ��7ґ�e}1J&����*�N7�wr�5�(��0�(���F0�g��(/���qȍ�΅���B���sh7�?��B�M�=l#���{kٙ���D{(����F�ؕ,�2�]9�j�\��Q�{�g���q��BV�/-�2�Z�R�K�j�QY![�!��a.@
TN�l~co!��C�(�^�CnD�v���' ����'8yy���ֹ��+���ҥ���ҩ��p�18'tt��쏍;�Gb����7.Qd��I�.h�&[3J�{��X���)sum�h�KH��I?N��,�4�Z����_��l����`���>C4�g��q<eL<$�����X������� O
��~z�2��lc�"M�4L�9��x2�pk��nJ�C�3���� J��q��P�����5l����(���>l� �x:-�R��I������C�9Ń�7��I��j�W��[:L�Ğ;�MD�B1�2��1)�-�b*����|�������<*���;Y�v��+�vP<���� ����4R��~�אc{�{�>�7��ҹEA>�&M�qG�~�wQ���Dp������@O�C��f]E��aN� �\N�YH���#�W���e�[^Ӫ�%�@]d��P�hԃ�DFu	g���O�U^5J�M�'59��q���� ��k���[x���p��P��t��ajBf�0;6��{�dq�����^�BTmfb=������ʚ��B�-�M �j�N���l�"�}uˢ\���{fq�4�.�nq�?���/�CJs7I�[wQ��u��Vc3g4\�p4�Ϩ�jO����Q�9�a���35��X��R�����%[�G��>.T1mʀ�Gzݪ9+�\j+ �^rPIKSN4��U�b���pj"���H�E�������I#_ă�g���
�����3�$�9�V5�����[˕R�╺^��Z�6;)�h0+��v�0r:�iC��H��zv�I��,2`�O:�ֹu�7ŵ���"��˃%�1#Ŝ(k;!/�u�Ɋ�rZ�q̞�.��f��~��|Z,K���1Fwp.GP-�L������X�v� j���?�?Q,�W�.�#~���:�ds8��e���XC���(bɄ�w.�EދL/�h4+�������)+��w�[Ѐ��,�G̰<��Yz0QC�yVؔ4��[H��Y���?�O���:1;����&2�0"6����8��mc�{�
~ٻ���C��o��mZ'Ľo��'цH���X 0�a�>�GL�4��a�Jv@4��^���P�?|I�	��"=��Z��%w"ʯ��*�~Ќ�h��@^��tk���(��u2ꆀ��_��1���W�\`��9����W��t��U�[��?h.��:}� PeZpl��b
�D�����Xz�@��@��)m��X�m% ��"X|o�~�����պ�@����lH�I�.@�8�}u���~�?�h��p�f�±���Ix��N���Wȅj5gr����$���'d���@�%�댎���C��T��xg�Q�$H�����Ѫ1�+�����'Ԗ$����h���cnS��a
�e7/����k����qn��
��M$�v�i�IlS� �v�*��v:�L���-G�I��uO���'�4gvr4����Tȇ�.���A��j��
u���@�ʐl`2�[
�l�{%{�����a7��G��0��9�"��a	�������ݘ�^Y_�]�&��9�cOa`塨 V],�W�h��R%n��Y�A�s���^P��el��BY�$7dn����}��)�?���}�'����-���� ���U|�P�VS .��GΏ ��y�R&	G᯹�,�;[��3��ʐ�1e�#"����H14=f(.l(\��m��
�ȿ�=��6qG6�2Y���#�m���-��Oښ^+�1�G������!M	2vb��B��t��y����1c��v��]2&wz�#ʤ��&O���h��1�j5�H�1�d�	��hP�:Ƭ���,5�~mH�^>�H:B��ӄ�ʈSZ�.b�Ns���IwR�HD�᧣���a���zF0�c;j�'�uYP��b�C����ϑ���";�(*����[�$�����5AH�=*oоWZ���p����������������Lɷd�Ս@,њ3~>*1�GWB�U��/�qB�����b��H6�ނv��Sy���`���9#�06��C�=�:����s}�&�4����E��#��\��DL�K��t?i9�D�n�C�Գ��r\qRGT�M+�5��']�^}#�F�����+*�}�R���D��W:6;�{0�Ա�*T�#��i��As�Z�Џf���@+X1�?Aǐ�i�w-AC��O���O���lI� 	�)�y�)���Q��JON�gyE�w
j��6+U:�㬶�=�I*���eO��jx�Aϛ3�����`ܴ���e��S�uiTɍnzӐ�F��A���wCF2��� *2��/�ƌ�H�ct��D�C��8a�����
�^�I w,����p��0`|ҞlϏ�d�l�e��Ἐwܯ��£ϭ��)�5�9��pW�'�V�~!�D}H�)�<�P��opQ�d��.�Z���YW�KȻV�4=G�(,�8���x�ⱞ��0N"�1�>Ţ7�)~؀mUO�,��8ČI�`sz�k�V��{2b�%����,�V���'��J�m=~ĸ���q5�݊�[��UϢ�qYZ��k���If���q��`#�3���1����n�\�Mq���/;8��3s�>61��jܹ��J��o �`�-b�)�
C������s�@���b3��n�T�Edǭ\ V����4���k�Ἧ�s�{�a�4������=��f�����ண1|��#�~��`��c���d�c׭-�C��.b�5�B=e�����ЮZ�9���Q�V�,�m���V:�k^�|�T��AE�-������	�Lj�)�x �����WXy��u��޽P�'��9dVYq�g��4�bN�U�����"���w?��W;��f��py@,��dg"@��+���4��G�Wt�L·5Hg>u��c���Ծ�=��/�� ���j4��{a{�eY�(����,���!ha\�1�""o�@K�pwӥf�C�v`ǧ��M��&.�M�;�yW.��7�-�)&?X"8f�Y����z����F)sa�T��9Ҽٻu��h�Eo��X���G$Y>���wXj3Dq�$�R�i��2Z���ܭ�@������ dQ��%�T����f�^��=^���##��Σ�\=Y&�*\�NTy��K�@�u����%�[M�I�I��hr.ÁS�2D>��jf���XD�މ|機�F��q���4{�Gx3���
>���득��<��� ��*	Ħ��,�ƅ۷�����q���-���Ot���:�>9Ka������@�
��XX�$�}�EJ�ٷ<�Q����5�\�mcVL^�+�B$v��ڂo&��Yu&��'�B�wР�B/2��O������:nN0h!H(ձXn�R�n�)�PZ��;r������!w�m�����ۻ�Ys�e/D~'�Q�~�q}ꊞw�#��-_8Z����������墊<p�ʏHs��T�٘{3��/��Ȟo�Wt��ǋ��/I�PJ9���0U�G����>���1g	��N���
p!�:[��# q����u��s��&��%���}�P��4qVN�c:$%��d=փ�*�Њ�+j`4��l,jGQ(����^i<b���:L�߀E���ں3��r����l��/���Z5�di��P��3N��(u�a��h��4$��9l��M<�]\1�������������{���nz���Hyx�ZM�!�.�&����uIKd��ld���Uq-$�Rf2��X����"G{ěD=!}���M��{��P�}O\�`&̀���`;��+����o�VD�k~�)j�`�����V+-�bL"CG�Ew�s�<����n!�I�N'����&&Vg��v"���'\'9�ĩ.l}�V�Y���$�"`��y{��`�_ջt���gͅm0R�~�"z	�:����b�G) �ɭj\�IJSډ�h������ͿG|$g�o�:�!(�r�2�����$�oՋح���F������/�2�����y��� ̯�i).0I���1�Zt���Q�gUfF��ʘ��Ԯ$2�Ʊ�	��fu$�@{�Ɛ��xA �4�h��$��`�K���,��q��cGL�I����a�#]}�DI�e��%�Q���F���JE�.�'�]O���I��������E2��A�ѓ !{���@Wr����+"��}���J@8������}+����5�Yi8�hv��W��
�>�,�U��I�c�n_�5ꛣ�p��������GW�x&�6�c�szU�B׼��[����tE���I��D�����5�#��B9�u���w ݯf�yݬdm��)�^��-T��pk.��]��n�����]�?�wg+gKrHx'M)
�c�Jv�S��܍O��Y�!�D�����B�sCɏ�I��h�%u~���G�� ����h_�F��x�Ǹ7��? ��\B�R�fZ�[��[�:���Q��$hUvOam6 �-���GifuL��`t��w�G�*%�Y¬����-=��0�
�E�
Ǩ�kXǻ8t�Q�? 0Ńu����z��.���x��#L�g4uH�4^f�l�o/˩�o��K���kʈ�� ����A���R]��#����>�TZ��������_v^[.~������b���x�Å�����Ѻ���5����k'��0���%y�9I*J'V�� q�Q�	���\�R�N$�-dJ9���D'�������N?���o�E�6���NϞg}���
��1Q�A�[F�ln��u���3�m���\���w�li��L��%�!]S�{���T�#"Ʊ3�f����Y
�j�9� Χ����顏����ך��:9S�K���&����(�ޜ�2��)����N%�16`���8Is���+��XS<����d�8*X����&GKhi�x�����r��*�hOڣJa9n>}5���ۃ�K��������{7�+�D{��k�oʤ3~��Zni%|�_�������V���ܟ95W���29_��0��z���+���}g�A�������$����k
lHlFx0K���r�U����	�q\�\�{��67�#��m<�z����e��ת�!3HA`���Tr)�����ϲ6��<T:�pP �X�kv�i����o�"���@)T�PKc���9���C7ʨ�{5�����h�q(b�Y�Ύ���8ĿJ�g�K��'�h˨�+s�eY0X�[��!�����F��ި,�l�w�F�	 P��6$�O���:!X���[!���ܿ��s�L��ΉL�3�Yz����7�0@MP0%�DpXˋ�:�>'����j�$^�_.s��&�n�/�:ݗ��ǈ�sd�z){Q�7��t��+1�c���X������(�$���s{LF�J���L;:n����y�jv8{)(��6�]��V��e������s��g���R"�Ǿ+hR+����E_�H��ګ��^��*�'�n��D,�<�������� �B�k=s6����ID9���)��oʣc��YfD�`�Me��(���g��u���H�:���.1K�XDn�f��ǳ��'\q^�m�"!�h�B�Ï�v�}'w���D+�P|[
I*��|��1���t�����G#0XM�<Pm��E"vIs5����#�Y����r�WcSv�W���4ߖ�W�}�@e#SO?����p��]ٱ�蔉�Q�_��P��.�h�Os�%;�uwh�
����?jP!Źa����X���u[u�\��~%8`r�G��"� 4l/Г�Ƅ,s/���M���z��6YY�,��7�|%F�&mȗ09u�0���u�0��Vͻ���Kl����6� W�kp��5��i'���|X��mᾏ�3g\�?�4D.A��0���,�m.��̵�[�.3�aX�z*>eb�R�i��/ȗ�+����
�!/����s?��#~x�_��?AJ-#��x-܅�k��L�^1�_r�;T,�u�u���op^��礖e�Nr2F�/��q���$IX��;|6�'5a�@Z��D0H�1j"�J����¹�o�/ ӷ���qA8�Z<� ��c�o�UZQ������u�F���كR�t̞�ذSę�U�H��{L�s�^ԲSp�E�j]슜����QU���Y������pQ����^C��3��Vpn�	��@wYR�dЍ��*-ТJ�IQt��6	�W
�� ��g�n�/���$%��$�Pp?f�����$�Uw���1c ���7���`*yc��s��hBH�~U��	eh�\a ��iv�C~�~[ٮ�Dq���ܫ������I��%J�i�s#l�$�Ю�-=r��,� i�r�����{*T�U�-��vL�EJ���~�l���皓�����䫅�Hȏ��?0�Y,����<sj(����f���~�	�^���bHJ���J_�Oi�=qW���k78N�g��WH��Cc��d8�ژ�c�u�n!""�ֿ��>�s�\�=�Ȭ�����}��F������Ƿ�N�F�����x�f����9�zeU-���l�W4�H�d����2$��`��P�{ ��?�{����<��(ə�S��ND4@U���2Ƨ���J�r^��e��^(؍���4���0f&�j��/ �B8j0����q�I&�)�'0�]���K[x@<Y�Ï��s�ǥr4N�j$���������"!��?z� 滯� ��\�V��n��z�>ϒGe��Y�"�M
f� g�Ԭs��;�䐪�Y�2�2�]��˒�6W(e{���L�*Ȕ��E�N>5�5H�G���2�G��%;�-N��I���';�2�$F��5��*�o�U2�]�L6'�`�26�%;	f(k ���*��c���]!=��|sq�dGG���[ �n�e���/D�1$_�������ipT~��b4ƻ��RL>��TR�~׌�`P�@�	����������-R�]��*���~���]Z;�jv�s�me'���bE�E��DÔ5��$ukЙ��=�����aN��RR���њ�?dFxk X���
�tVcLO��E�iB�گ#�@`�3
�O/B��������E�8!����+�IΔ���%e"|^L/mv���N�~��0^���Fe�/�������f�2��Ϯ���>�zg�`�r�[�,W����w�֭���}����f��D7�o��hwCz��@��{b������5p���1�C���j�t����������ҥP��&T�x�!v?ia��k_0��Ɔ1�t�^\�b�eu��>�C���2��'���ڗ�M�����WD_,>L��06/XEK��6��S���L�U�0����oN�kT�!@�7+�4�j��x���z;G�#������IFK�bڼ^�xoJAt��oi"�V]�m���jq���!���knI�.�����נ}C�hE�Р����f�w��k��sJ-��/��)Cpo@�-j`���C�B���{��R#��В3 ����3�v%��9�q���,�)�GQ��{�X�ÅZ^ûp�������,�q�D{�����'�ƀ�3le�r�n g_����l�E�������wfr��s°�遢ڒ�� �z�"A5���TS���Z� o�,U������=!o}���h�M?F�K|i�`�}ۣf��=M����D�~TˢMn��^ۂU$q
]�a�S�h�@=�^�)�@�ޘؚ-�͕��٬ը����@���>�n�<nY�m;����a+]<�fG� �#��y�7ɪ���?Ѵ��x�wM����x����Y�bd�d�#i.��o> �YC�{�M�����wQ<��<̊B��#�`p���p;۱t����B����tw�s�J�	���Yh��p��?'(�r@/��eM#�є��I���`3��C�Cn6+��SI�\}�AU (g��zrr(2�~��P�MƋ�D7����i<�oAT,��W�k.�@U֗���N���E� ���
�{�TJU4�0�4�d�1����^&Y���`S
P�J���N���5=�P� ��Ƅ;�G�1�Bn TM.�?����x�h����wE��I��]%9��Olk���mK��0�|��o^�T��=�!�Od�o�[�Aμ��Ja�1���v��U-�1ʇ�n�X�h�7.��
/��	��x�l��bҜ��k��Mͳ�>: �f��aɵE�ع���K�Z=j7�ĩ��#�0<([|,����R������ug�J�p�D� G�kv=`�3���p�/�R�7	�2�s���*�HRɊ����u��.���d@��ͨ�Np��E�B�c�0���Fe/�e���z�U޴���B�#�4&
� ƕx2����=[�n�d��'�b��ed�p�`��9�����Z��)٩4����@�m�~2_�a{!?�����U�5�Ϣ�C�"5#d��`}��6��j;���hN�� @F�+�@�tXIG�N�-���g핾�zQ��
���K>O��A�m���R<&��j���`�c�͆ŦN#
��n�W?`�g[)�'�d�h�^p/O�vB��]��&h��O{ ht�%�����J���ہ���	G'm���11���czvI|�2�$Lo��nd1�	��Af��i<�=�B��z���O�?$��h���aಛ�o?��آsN�*�;������/)��n��-�c &�t�V�V<G;����?oP�D��>V��Z9]����w�{y�3`��e��b��:�Bc����F����wФ��5P�w�_j� -��3ϓ�4V�
�8�4��1��m��`6=�)�Qyً�G�*�fi�'BY;��J�JZ��0�]B<�IT��R�Od��J��d��5{;g�+JΌچyO^}�f���l�j�-��$�[B��8G�q^�01�֤
�PM7��?�I��2
?ch���O{3T_5������M��^6�"�y��,}/�ɁxxlmHWZ�g�A���������v���jh���q���D���z��)�����s�vW��5�K[��E���a��(��,]�z��45�i+șr�H�����C�:ʧ�E1�E�.��b���@��g���0-�g��ه�3��xy���yR�s���D�Qa�W����+X�����t��E��(w݌��3��/���@��0�E��o����0\ơ���L�:�D�;�yxքU�� 2��̏�P�����p����N\��z���3�\��7W1c�p�8�hș;����=�� �,傢2
���<qa�(�eݞXr����sEG(_�P� ,rޚ���5��Lf���7��7��E�k�zK�����`�kS�k�+?,֙�o���xb�?�
Q�47�4S���Z�ߣ�����n̆��+��S!�'K�G$C�2����s���s6�qM���@47P���{4����pwnK������a7ȃ�1|-�0N���W��s�SJAG�V��`�&����
 ل��+<q�0�?�*[�����ܳ����=���"�����F���5��׏1s�MZ�f�$���|��z*��y?�B19� �-)��ޚN�w�M��j��T8!+p���	��+�R/��I��B������$D)��*%��Nh?��?$���9Q����Ny�� �����.��-}X���SP���]n�f�:�j�y�L��RK88w�v���F���si��(V���]9 ��g}{;�hs�t[5e�U���c>k7/�8��0��?����t�y|:/�y�[�Mq���{G�r�1Pp�*�tDC�l�^5��l�|�^� ���R�Xm��I�\�e� �
ҙ��zMƷ�_���^��p}e|����ͳ��v�d,���z,w���J�����{��)�y��rS���+����*-a�k�7�2f��
?5��5��m�mYy8���~	(Zd�Y���,��{��"x��P���8�h���y1J&�}y(�%����ɪ�#��~#S��h��@Jl؎�$��_���B�Pf�y0n�lԲ��������]��4�]+�a�Ը�'&H%�B����d��A�ˌ�J�M� szDyx��J�a�A�p�#���=m)�/�64��}��U�`���#n��q��#�y����
�h�*�a�i��H|� ��_��\��k*�Ws������Z�|����^��7d ���^���>E}�c��X��}���'Y���"~p����z��������8k��2���!nN�����rnhD]Hf��b�X`�����^!�j{����k�Q�rɨg��
<���I�oIN匉Qŧb�;�I1�:��;}W(ʞ�>��Hd��l��v�C��ł�뮠!���Iݭ`�6�F�C��<>\�b:�B@{�	*�6���Dw���K�O��{�b�9x5|�J~s��n�\\�Nt]�;\�g]]u���@��O����T]���.�`���vs4n�ŮP���m���߂�-�Ӟ\�|9*� )�\�wI1$��M���8�#y�':��Tb�Y>Ԣ8�j���fǸ����E�|���,X>��9Q(�-��}��v?Qr���d���j�u�lՑ4��ʺp��a���*���<�5
�#�`\4��tK%X�)IUT�q���"bL�W��.��s;	�Q��gL�#��Z?Il��Ċ�s/Ӂ��RZ���dqՁ�]�[MY�A.QF�s��$	�`WU����$�?��O �,wkm�9zR���jU���9'�/�@6�dK&�ב>S��)��j�`j�ASu��C�3������r�-�ٱ�ls
��L����\��'�(%$�T��͡����
�:&�#�@q�v�gO?��U�R�!{�d���CH�P/�/��ɛ��R��#�O�uG��K��J,W��H\x	k��2�5�b9��e�̺�a���Xs�5w
	�xP�.e��K$�m��n�M;E��M����aY�[) �5�z�� lP�~�Y��e[��E�D���"?gFl�{�e9��_�3H*�Yf�Vl�#~�i�'�<<|�+nk�����T�s��s/(Au��>�/�g��4��G�K�8��\��*x����Ӭ�Y��r�zk����V�T����>Nɲ ӱ�ix? �� ��ٰ�=VrL��Z�3��W'��>��^�={$cޒz}9*[�a����v9̲�J_�2��݌���NLk7R�0=@���+�.��ΦyA��4z^�]���tF}��_:�	7i卜�=�f��N9�@���9\��k�Ɯ���4��<�8��
��������$��N�K�n/Z�H@���_���6L���b�]X�n����P�}^�p������"uCe��+�+�6�i�Įr8C=��Œgj����*�$���o1`�]r� ��ɣ3��#�\��vt� ͳ�2�f��n��0�:7F��!�m�Z.\�Q+�6�P�ȑ�#�,���D2�2{t]3!$�Jl�b�����BkxR�\]� ��g��$UMhytb㶲�K��\,j>.V��AD��q@�W;�M,�g������ �Ei�~���16lqQ{dL�i������	�e.��1�_�s�'���3/���� SaϿ]���WrMBM����������*�*��L�X*�4��Ǥ��"�Ѿ�����Z�Wr����V�>x�_/Dh(�`c�e���xEr��߾#��!�
�%8�7"���a�2����E,Y���V�}.D��iW��|���ެm�~*ob��v�ڴ�5w󔨨�.%�^�e4[!�����N�b��}y�A-�����f��VR��qi7�ؑ�4Y��&4/��`��K������%�xt��'��v�J��[kźa���+����Ze=���"�if.ɑ�#j�������o�#3�qz�wØn�B�̣�{�@��*���8@�aSX�;k��C]c	��2��%'��7���6+o�U�q���ϫ{��p����AKf���t�H煱���c<m]4�"� ��y�/V1�H�C�e�2)�=���ҽC^lL�Q�NFO2�oWi��'��EN�� C�'�\���ER�1߱J���5_`[6o�ѽY�;��9w�E�E���b<%/r��^屸<�Q$QQ��"6'%�q�^m{�C���F"M�p6�A��K��2dQ�3�Ɂp�FS�Q�]�<}���&�R�Խ=+ƴ�`9M�WX��!�XE4���Je!���y.�dс�x�t�K�ix�m6�n�3 �2$�L�́�����
�[r\$N ?��)h�F;�������e��	8�\.`��K�d&˵�Հ�Jg��fz�fi:����?��
����X
�Er~���`R��$�y��7��׸�����Vg�
M�܍��!��')V�+�%ɤ�X�7���=Ԅ�=%Z0�_O�X� T�ٺ��=�ֆ����;
7�Q�:�Muh�Z�J�#��7{	,@]��\�q�5jUM[x����-�| �� �578g����o����
�?֟Q�GT��O�MW�t�LD]�P�ݡ!��b�A�i��%��aO�4���5	i�̛~qi����G����9w(��9Q�):��-`�>Dߔ��aW�A�g�[�HV{F�@�43�/��(��[���pX1�#�8�;W����ƥnX�dew`ͳp���MY��-�s�*:�^��F�_rD��?��[�A�!��<���kD��.�4�<q?IZ��9f]3S��I@���8���3��R[1*�/���A�1R��U�����ͤ�JA�k��H���$�qIs��3��*q�>�2H�فW�I=K�S�'j9"����*u�s䇏��p��MP�.���(6x{�����f�͈�e�_��w�w�>%�DO�����ʨ�=�A��Ơ�ᘵ�	xj��3���S��kzVC�100Z�]G�щ����kxa#�U�c�ub��|����3��@�L����1�v��:P��!M-�	��S,�@��{�3T���t��>�u4p]����z8�6a�y�����sAU�k�{�?`O���+ɉP>�|�pq<�ݼ]w �1;H�� f�{�i�|c��J]2A��M59�`��mVqB� ����PW�ņ	�uZ�/*��1�F)��S�l b���h�;�Z7��@�3�1*�!��A*ٽ&U��iY/�u��V�}@�o1�|yf!�a7;�^(Dh��r���y$
y�p�S��
A����i�+Xd�Ȥrpk���-�����d�|摋�FN���t�p+�fG��tVf�06G�m<�S��$�d���$���sO���NeMo�*Q��&3�b�W�f���hb��4�MmDm��
Z(Ҽ��y���R��Q���ʼ3�A�����O.	��I'�pT���| <Q U�)5�wr�M�m�T�P�}�L�Ѥq�l�yx����'&^,w�Hb���٣,`�6N����gȌ	E?%�U@C��c�X�{$�u���#���#�2��$(�^����[&�N�F�BY��W!S�v�r�jX����nw����rʆ�7GS�g)<4�r������>�+�ʛ*��(����6�ޖ���E�גL���Q���c����DJ�̅�h���^�I�W�D�{�#kަ4r+��>ET�[ϕq�,���:���� ,Yu��qWeh'��uOƺ���(�Z�\#�3ZuwT���jQ�t�|L�j���z�o"L���a�#�:5���:W��uHDz)����*fMg)�+�2r�Ĵ�,:��ށfYS�E���ƝT���H	VF>�w�8a~��`A5�� )����C�;aQ���Q<pӂ�?�N��9`	��� �1�EsE?OR����ZgX�)]������?��i��,���q�1�M�#X]����fz��P��`�M�@�"��0�}c�Dg���H�0$w���*�[o�K=�8�]4��lC�m[آk�mt;��M��(eM�m�:������%���^��x,~^`��%�D}�<�3TJw��:.0M:Ɩ������ʫ���A{	�sK��@��8 �o:�O����7����D4Ut걐��㐒,en���3c0G�������]��:��R�|]ěux�v�,����(2�skX.�g������I�B1�JYk'�k�Ce�$$;�k���x�`����; �y����I�{Yڛ�)?T��)"�!,"iD�uY[iҒbG����)z��TP�*��������1��6��b�j\{�8� ����b�h�k����M��tC�� F����(����"t 6��mEl8��bЕ2�h;�w�V�����6NH��J�1D�[w;�p����ɚ���8��36�-��]M�(�TÌ��;��� ͸�����0�dvr@�u�h���)u��潚bf��i�/\�n
�Qt����Xw���`��/)u.q"�-�~�N��*���.��0����|o8
�7���E���/��nt�,ׁs�{���HQ&>�W^��th�0;�_�W#�b%�h�*6e3Ucc�'z���:,���3�kE�y����䃹8�)����gsu��f�Rg�}�p ��o�O�s�cw38ߔo�l{3�d���*��,��6�~uq�X�s��!fvK�?T�I�c�a� ��]����]��6V�=��1` �&��Ȧ�����&@&�NL��IU^��o��7�-z�?��}R~��Q8���ϯmj����X�_c�.1Ѓ >"�H���6��J��HI���}̶�u��Lǖ���h��:Ba����a	�n�s�<���^(�Z���!����tPd�ElP.۶�dm����ث!8Sbg;���p���� �3���S���=;���V=��r��י	A��s`���G����3^2�x��H��N?���-v�(��E��gn����^\�^Fl�߂q�@kާ�$�{\���NC��[��^C`�9	X�ܦ�ɖE�9��8pƗAH���r�q���4F��P}��Ż���)"Y����ZR�n���\�2o�����k�v>2���a����B��V�.�Yj"C�L��6nC��f��x�	������_@�J��� �]Ś*K�4�az�\�r���D�^�J4Zh������LP#������M!��D&��ٷ�wՙ��F�_�r%�[N+�lf�,[Drv�$� �t�?-�A���21��2�����sZ��*g�
/:{�9��"�ĭ	�E�yCu:j�3}f�`�7�r�5Gz���q���Ҵ���)�4$c��O�C�Kn�R�����`Q�?��?0Ko��s��tN��)/5�j�P�2�«��qz4{�;J��,%w��]��v����_'_v>ѕ=����E��疯l�>|ٗ��1�$���,����x *)e�����z���ݜO�y�$��N�w������)M�*���eN��#��F�t;b%ƕ������57K�m��ի�=U�Ux저~�%��U��?�
�&7Oǽ?�rb��&�F�d���i�7,�M �%���(yG���:�Qr�h�'�$�Ի�sּG���N�\_$m��m�kŸA���Z
?�S��CCN�6�t��p�������#/T��ɰ��0�pA[���M�r~���ա�0^证F8��
bK����s\.�n΅�����1�q]��
ٞ6�vA�#<]�=羇ᏭVVX��+��Jz["�"���|�S|s_�6!3��`%z�|PQ��Ú�D��h~����A	���w�T���!2y~��yR�1�:������Q|F{@`�Y��O���r`��,�P���/R��|�@��[��+K��*I�iq�ҽ�>��EkE����!��H���7�S�A�,Τ?�}�K _A;+��ľ=�#t�?�]�D��Ē�Iqګ��5R�p�2yw?�¾�x>	���%�NL��>�7�
�}�@���X%�N*���i�X��{�jѧ%m�Ӆ����wE�Kգ4�4����O#k�}Te���OΪB�~��Nd�Z�:M���'E�Z�ͥ�i���ˑX�2ѢI	��7�����m�VXl��'bf���j�> �"!��B&�I�bVi������ɻ�ǻ W�tJ=��?tI�hC���l�f����q���-��Pϼ L�u�hD@��������k��zc˪{lZz]��kI~�҂���{��ID:�cI��j��a��Y|/��5/�Y>�I5wL��0�>��[	1�C'c�꿃7��Va�yr�� ?�F6�S��ȼ�����r���M����Vu����\��_Ė�nsh'U�&��3�����_Kz(�tl��q�R�r��ys�Rⲛ�*�T����t0ǲ���k��g��))3Ԇ��& �U��a FǑg �������Z΅YU�X!�!��<�{4��#�|5 \rsy���opz����6�?�<��<�9�����×9�/�1f��K�!Ty}��6��{n|�m^����q#���G*���r����N;�2��ޱ^ˊZE���"A���eNK�x*�Z{xޭ��\�������m�P���\�lR��Vz���C8���`������h�Ϩ����Y�JU��ێ-p"N���H��z7�	f�>^���˛vL屫H���9�B%��3b�*��#��[�������X�m
"�|ڃ�<iHQt�/�0���'h>,��.�|[���Bw�}�D�ޯ�u�97T�il
�Nxǥ��zgҴ�`-w�c_~>�1���:"�s���0;��\YO3z�������	��+D�2�iGI�0QAK:��s�t�Şf��[��Fsh�-�{��'��!���]�n1�{_A��w���]��������M����X����e)$�3��>�|�)�P��3:�H�_���l�4��O�ӥ���'�=��"��r��xx�"�I�ȉ}c��qTH'�}V�@��^һSTǜ��.��f�y5�/�$c6ce� �R�o�>| ($����Ne�8>-���`E0���'�9� t����3KHݹ%lO2�-���w��O�$ϲnw��v��|�%e�F��9>�"gvM��jA�>,!fU��X�e�����Ҩ�2S��Ms70�e�(���y5��K ����f��n6��%T� \��ؒ1��LNFe�7y�7�*�4������	"@o%�k��Pl]' ���#��E�@Dv�L�d�߅��R�v�"���hA�� �����}3ި��
���7��r��D��[���������ς=�½z�KI���h'C��,"Rpm�j�WT[�����h�y���]<�DQ�[�c�0l��r6b-�BéT�Z���F�'�qS�^KVEzS�njgK�Yr3���$g,���S�]X_�>�R��t��vP�r\ ��(Ač��������V ������a�ɞ���H�g�;�Q�e�)z��7:
>[�:�dꑾ5R@`|�"��-el��?ڪ��y����\uYD�T�/�A����K��1�;�JO2��wFAJb����2#0�:��"�F
@���uk�zh�[q��G��3@h����d�E]���MW?60${`lR��U𕃬K��-C�y�9���g����8bN�>e����/ߋ3�
D��*,;֍M��A��}�<j�!l�,�ɚL��8�� ^�}YUw�5�+�ʄ!'`��)X��:j�cWR��H62�&+�8��\B�����bt�ט<�Q}���(4k@�s݉gY?�B �nM���Ù��mC���*�:�D�����Q�D��s?��Q�d�]�m��:���Q������E�ھlp���&iz��|+��̭,�0�x�1��Z���|T�lwk] D��rh�;��|��J�����:�عr;9�X�z��ofI$��f�'�/�n�S��2�
.�[�8��*Q	-Y�;�,dP ����Z�T0�b���P~:�9��bpYSu�[��v
���'�{i�� ��O2,����6�*��^!t_Q�_d�q��g�@tr*{�o~��8�?�ʊ��8m�Uv|i�;Wy�=ۦ��.�H
�`��U�����}��V�_��Cti�M��J����a�)/�P�Ԡ��Ҽ
Q�a�.�쌡���Wת(�p�.��6q�bP�l�L�V��T/zi&.������|]>\��1fq�ڷ�����P6Oʄ��,,^`��!='8 ��`�zQf������0)n� LC�a���<M�u�������
h#B�����9L۞.�iѪ�S�}Y�$��e�iTYxcn��_hE&�(}�&��-b	�4�T~�#r��S��iY�H�=<���>���V*,��6nQ1<B�=��P"J�NO
����l��Y�s�gB�u �b0x|����V\b|��Z�~`
#H0��3��w�T�`�S]-�.�:�ڤ��S���̿�e�q�.�nR�`�7O����ۙ���5p\2�+����rK��fk@�5�����~=��A�T���87s{h7�M��uh�y��&�3o�C�\�]�Y�8�i���:�D��G�шoE�F�끀n��䮇�J�^.t^�Ց�^=���0����I�OΛ����'��X �=q����F��y�bc�44�� &�qH� ţ�Dknh]|�s����Y�ҁ/�:7�ٖ�����5ż$F�x�7�T=�ZF�"M[��@u?	��D~o��Z��G���m�bw\P%C�� nD�;�[� B�Y\�(	y�4i�#�9��AD���U|
�=2�Fn4�G'���L�
�m��4��U�d�~,M�m��we��ܛK�*���u�<�|h�Q�NJ�y���j�T�Ĩ�}`�C/���m���! ���7�9���n��-��d�>��xmJ.���2|�����k�"}�����=@09��[-�K1^h�&�I��}]۬);��ܧ9@DQ��B�3V�����H�~bEg7I֝�pȑ���� D�%Vk�3Q��Zx�
9K����3[�9��R^S a]�C\z�������+�W~NQc�č@^�]@?<9��mkj(0ع�~�A��R�؟t1���
�>2��S�������m6�|T�tV��~�0�`�c�-�Y�K՜�-��/����JxtZ�¶df����N6PLPl���*pFI�Q�lY]A}[$U�}�Q+Ԍ�*�G��y�]���5
n���YV�
�	ɺ����B�p����rȨ�Toݒ�p�2�<W�6+��$�>�����j�3M[��)o�hP����&!���{���E�̙�z�>ϻK���2!�$����4�=x~=	E�y%m�D��a�\olAO�Ƃ;�0/��:V��C�L�d_"�g�����P�h@H0e��_K���>�e�,�_�u|A�ۈn1��4�Mu~�(�Pfml�49cK�͟������0�O���wzb�]P� �hIǞ������o!�0�+T��4��nO��7UV����N�<��H!��X ��!pP�9��B�<'z�M�y��e�n
�[A���cq�޽���]�����9��8SS�e��=7
�Ӎ'�[�:R�V��~4�k�LE��Xn��C�9�((!�DӘ �@74BB-`�l3�}� ������Ϸ\�<*���>�sSC&������a�P�u��KTl�םɃ��`��@��#oT�a{;��-��r<B4�3ߎB�/���ϋ�m�¹%$9MM�u�%ǆ�WT7���b������
��>J�%�̅G�f��� �3�@w�ѱNV$������]�Nf�o�-v.��.r���|�+��k�c�ƏGp�Y�b��H�oFVm��#��k=�b�h�ǟ�Z�+J�E"��s���I\(^m$��c��h�U�ݎ�b������+p���z���0���r	B��d����B
��&G�k2RM/�>�K�e:Pw^u���*�cb�=���-�X���B;��ӭ�ۮš�N��Y�q�C
8���c%��lZ��q�X�Q��� �1���7���g�!��*v䚙O�$��K,�P�=�G\\�,|�6��o/i��^�Ŀ
S�)7�N��4�VhF�f5!���%���"�7X;_�i��\`�SY~�t�K7
��o�z^���,�ɡҞ}�!�Z�U�����!�Z-$��PqhKR�۹�y����Ә �,r���?t?D�?���c�VXۑqχI֑֜�-\���gq�3��D������`1��?���Z�j����O��������rB�=�,5��@�"<-�B�F�%i�	|������a��Ѵ�`i��(e��5Cq%Z~��$P�o���Ў�=xL��C�W��{���~EY�F�����߬�n���|߈! ��L���T�^_�cwM�, �Fտ��Ӡ�K�'�_�h�V����V�zRf������*�@=�x�k���]n�`������]&�*B>㾔����E���M�e`NaW�B>A���b�D�S<���!%gl+삱̧{�����o2b�⢍A[���1i��ڋ4����Z-&o�~y���r�X�U�>=1Z�f. "��d���V��� m[�����񀳞c���y�5����Kbǽ����C�;Ma ,�x���F��VD8p�*���i�D:�O*������_�If-@⎻��{�#�W�)i�D;�0hb��k9�,�O: q9*l�izZK�.Z���u3>q���M`o�j�, ���?�ջ��?X�y�.����ؒ��,[��gvU���G�`q����Wji��Og�S0����S��I�J�́$��Iؒ�J�rv�y6��L����gGߧ�}�r��n��4gjTjT��x���W�׾N������cx�,9�S�O�T��]�&�~�) -��e�z���O-S6lҚi���(�轮��8,���V�G+�7�o�Չ��]R�����cׇ�c�T��N���,)D`��wL!\��Ԟ�Q��eL3�1F<��Vsc6b�<KC{���Pc�o�x�L��i?B�{?o�y.�_]��LR��7b@Q��v-�sw�.��XD]/Wh�bk?r��j�ˆ�4C���7�ݍ�8��|� ñʘ�\�y|���)��'l�d�?�����?֩q/�q	��Ǯ2����e� �Ƕ*�0Mc)'A"\�ѷ�����-�ہ���2�h?��)<73͖���DH<U�������'��.|��8�?8�^x�z�����0�d�U��
� ߱o̱i��?	���e�?-��qn����y6]A�䆁eHt��I�y(��M�����'����S��ّ4�<��͟.�v��[t�CK���R��+�B�グ�trk��p��>��jU����D(L�/�.�5*Rf|$�fF�;@kQ����Y#8����P�\���Z�f�d�L㬾B2V�N�}��VE�%�V1�l�e)㺑��M�������!}?��J�����`@� �N}�_\���<�v��wN�J��! �Bd�������MK�S��K�,7|F]r#%��"�t���$�GԷ_p�L��/�����(�]d�OҦ#{�����I�`����CT�9z��9=��:#i��z'o���`��M��AlD�@c���"���ٽq$3��K�����l��H�d�$aۺ���M�ja2>�1C�wz˝�e���n����*�#�	)lj�u��Ա?��G��l��d���}G�h �D �]q�$��V�xۇ/t�wz���%*\t�<�݄��*}����m`p)m2�(��`G��כȧ[s>�:����S��߾��u�>a'6T��P̨w>�dPdu�)�_-qbR�͐�<}tƒ���	��&�_R�����$���ZM5���>n?�3K1�� 3��Ș�1�Q�ͬ�xn9�4�Ò�I��	3���v{�$|�_��Co���<����@�����������o���
e�X���.�B2j��Ů�J
�I-�A�`ZT�	1�%9�^?'��6~F������ǌ�����q��
7��U�d �ۃ�|�D��X)���<D��L��t��.��k�7���O�Ȝ�M�����u#Cr\1����0 )�B@#�m9���2��F���c����I%𵊨=�h�Ab�)P~8�r����{�é֔�zb,Q=�֌gm��ݻ
K�sXᜠ��g�vQ7�Zqw:�_�9`V���ر�����9�}L�<�%����%��u�2�B��s��n�6�$hjԕY(�eT ��7���]}dխ�S%yc(�r��E%,Xգ����Eį����-H�Y�?bS�ߠ�pS&�����B��\&��ih&��Gʽ�/�O���O�o�<�:;�[$��K߹s����K�`\����b��,?Č���Xt�rt��p�h��b�B��DwvX��)�̙#���R���_�%��"c��$��M���:ĕ�
I����<������z2�_M��~��ـ�͈'	�0�8"��1����EGK:&��_��6d����THp��P2���ݶ4���[ ��ʿK@�SX��td�T]n�aj�>��Ē�����Ț�J�6q��������(���%n��e�\�6a����LA�{�5�$�y'j.5YZx������`D ���]ɼ��"��H�b�bW
U�W	��t���37�����	n���"=�C@�y���!/�K!�v�ߘ���e�H���ɭ��.���؆)�G�p�2t��Ŵ��@�3$��gx��C,�R$�:$#z;L���s�ꆼ�,�8�z����Z�l�g'�`�́&��v�|�p���y���r"� �d-J����Q�����L%eN«O��6���_v�\���\��@�z�����5�R��x��Q�1�x�B$AH�;2�;���u�I����և�j�^ק�[D��6|LO)wp]��D}�E:OR��HD�!���y9�J<p8{}C�*��cq��3�R�S�$X|o;hJ�'?���
��q������!bn�E����ys�ޞ3x���>Q�B(���K9�19F�[y&<�g��(5�f�HB�qXw�B�䗇����
����OU%ʧ���P�C5�:%!���l�'��'�/(�s��涯��pS�9Q�n��J�cD�1 �u�
d�#�fޡ���z^\gX9h�'��= ȴRUt�2��,@>��k�_,]<�T��ۙ(b3�2�PM�16�ϔ~n����6�$��p�ii�������*0�sk��Ar�/�C��oo��e��+��"�_��W��!,�&������4^��4ׅ@��s'"??W��|�S5�8X�i#º���&�H��7����.Н�_2����>����cJ�3A諄��R>K�]R�;0^����k8W�<�����1�ǭ�p�t��O�n��׼r�kVb��ӐS0�����Ws����6F���g [y�9A�s� ޘ<-8jH&�l9�:�H���q�0����F
Gw�ğ����壯t�t�#���tC��{l���'�D>�\O&	���Vr!4ܣ�br����zu��8��he�UCGdwR�]��P;�)�T�|z��tL��^k؅m�{��k�M ��В�S/q�M��Eǥy�� Y�#�II����C3��c�:�i֣;�F��p�� 5-ڎ�E<I����ǈ��@xd�Hሢ�-K2\�@!��E`�QB���Z΅���0���%W�b�e?�#|��']B
�p̫B+�]1��bp�N��/Ҝ�,��ȷ>H�L}%d�7�~�q+�bH0�̴�z�1�����B��ű@�򬴧%�@ �[����!H��ߵV�-���e�@�[Oe�@*��63�{�H���$�s���1,c�*��t����k'ӵ�"�{X���_V����@�3��L���k��3��X��D�B3����JT���ݨ@xC�U�����7�=���x5^��'�>Ќ�b2n�z(@�-u��p�"�y���-����xw��:�H�>�	�_s������6lB�0��,s�\C�]#�8ڋ;�I�G�A�2�W����(F�Y�ނ�ڡ�s��Δ��	Tzn�0�A�#D��늲y�L�P��6��w���й<R� '�����^ H��^�Q�Ym�}���JH��l��'� q^�P!��%�p�	̹t1��b���kW���F	X��֦�;�&X�\����xINYy1���oq��*�\ԃ���)_&>��uD16������;!����/3 �wA���[ĭ�Ѽ���d�9�2�Sra&\�4�k��T6-�ܽ�� �4;IN����n��၍Atu\����!9��&�{T��[���7l��D��表���3=��6�y�JE�����4
�X]�$�.�����@D?=�MQ�8��t^f��ʆŻNR~:�[��`xf	�e:`5LG^���'{�]�kq� �#�����j��J���Ԉ�c&� �tKE��k��w��A��#�<�Wj̩�=(G����]Ȋ\4�ަyr�Ԩ�P�r�ԝ�r�VE�0��>(x�����Í�j�s��X�Zy�T@O�L�fZ�3+����*���`��5���N�b��Z)q�6�So�1�4��hۉ fXk��`�Ʈ+����/�P�o9�����|??��n���Ȣ�ʪ�껬Bhf��%�\.�˽_�o�T� 
ja%�|@�7�����H���?.�����_���_ ��Di����C�cp
1���}�Uf�����NϺs��1ĬT����Y�����'�i(��<�7��Pi����l����o~!��it<���t2?dp��8;�>B�ˎZ��co�����dl���~�T�M�\�rb��%mGM��y���%pV)Im���ϒT�#����ad]Iǩ�i�ď9�>.�V=�u�kmv�~E}E��ujxg���R �_CU	)L� B�Q�a�J|������-)���!	6�W���ù_�*��@zY�ذ݃��*f��U@�;]'y��N{��L�c����/��꠷}��;�5}�;�tf�B���1
��c-��� ���l�����t��:V��^���}�~��r��	F�a?�`��g�M$�X�p�X"/i����Y$?�@=� tt"$w�C���r�n.�KB�����MY!�E�t������-u�����1`��F�dK��A9k	�������?˘��J8�B���T��+1��Jj��X���x�����_a���Z��>��7g[�<�f5�$X��(g��0������AYODX�͹:,kT��`&1m��o��$⋘�f���י�W!r6U)��S�[)�ፄ.�Bu��
���_��������JaN�J*��Q��]��j=x#�$%+�&���R���F_{���P��9�����2�=�,˰��C�u��^� �>u\=���J��5c
+��cꖮ��˽Y)'KA/�,�4�� �e�t�X��29,�gxתVB�*.�E�]�n�Ѝ� N�b��*<e��1�{b0Q���Z�o2Ѓ{*�у�P�����(�Td�{	�4d��7n�͞�X^rF�@`d
�YR��6~�[6n#���ע0?C�ܷ`?�"�4�2��F��Sd��^I
wr]�W��Z�C:j��
�Z}�	���w�ڢI��%9�9��1+a긴��+�[�K{_l12gX;e�t����{��2�ń^��E��u��Fg�lVB}�T��+1km�h:��f�Aa`2�Ҿ�R���8ʠ�g�f�*u�%��{%N�Yc5=���:L	1������.�TEKN����*V8N�	�5v���lD�~�s���v��2'���+��� �1Y}bϪ����X͕I�@.m}�;�7c�Xjo]����-15Ibʰ���S��]��wh˼Qܡ&kj��+�������a�~���V���v��\�%}��Z��yB�N��EE>C:��8�o�H��_WC@I
�bY:=l6a��/��E�zI���K��'}���O2=]�p���	o�@�⦠�bhfM�xdm�um;ß����FUe}�,�>V�g����s�����^�9WF<��=@ft|v�-�ѝ��Z@����ū���WC�D�Rk�L�(_k�o2��|ߑ\��ek��d�[,y���Vu�`t��\ݬ2�R2%�3N�*⺎�[�������S��	�-c&lT<k��ԓ��UF��x�8]��*e������h�W���ShA�oԁ�#�8����[���OR���ä�hn�bЧ�z���!�hV�1��F$O��'�����(GE�����.�>$ыǴ~5����A9¸'<����y��Ep�É͙�����\'���|�F� G3 �C/��G��G�W�ݣ����XI��6bNJ��<����Sdiu�Ċ�`��*|�֭�µ�u 5�T�.��U��"���OGE`��[S��K��֩������,�Nc�z4f��^-�7�`5��2e�P��F��FvUh��e�T1̮��τ��۽�^՗b>,q��:<DK��� �� ����,c�U�%Nޏx��w�L����m�?:�?V���>����|�/�������������(t+ 9E0f�+���9�%"�ik��CR�����Zg��.�GH���97o|z�F�4���B�^\�8�	-dL}�}Ԗ|h��j���F&�FV��������Q[���L�"8����b�ֹ|�5��ﻔ����+�Z�����4!��g��im����׵
�{�p]�V����.A2�WP$88�Ew9��_�uІ=n\&^EV�)�*h�eҙ�D��.k}HK�eM
Y�h�y�����/5�W!��w�QDɎ���!��K<��w|G�E�	���Z#��g��-9�LrC�ň*U]�?�wkӻ�&�n�K��[�TfUB�Q?�H�Qv!�1@7S��μ��v���(&��T5���4 C�Un�|K��RDȧ��O	G��2�k���AdeЋW���'8��35Jn)�.䈟=Yˤ��)���p��y��`.�n�]���*ŋ"4Ek�/5;��bt~���z,���W�4Eq��.�xԇ�C"!D��cƝ�ܙ�����<b���W[R�v I����#����f��H��hP����މ>uϧ\�`���4t~�o/�Ǻ�0V8�1��+���,������-l��� �����s8����?�8)�~q��}�K \��y��P�ڣ��� ���z�7���r�K~�^�	�2k�ң��coϪw�|Q��և醕�؀�;(�bO��M~R0.��[P�\��%��3�lb��	��"+f���� 
ԡ��Z)e)F��W�{LY�g�_M�0S[�C=9�q����s��`Z���ŕ����5H;&�����a�T��)�I�DfG3z����k�l��n���(���0�9p��pK���L��	z���w�[o� kǸ�?�����JE�C�$�r��2�`�����Q�q�^]�n�|����G���wW������r8P6~#�,m:�����^o���xt/_�������o<lx)I޳e!�?@d�>�l�}z�&S��I���^����)�����Y�/!�X�X�q}�I�$�B�0 >�ר��@JrW�DC�2��;�y����5��#kY �A~^��̦�zOPq#�k<Ɲ�
8l�d�a�C*�#��{C%��d�:k�.��1Jn����@eLp��r˗:������ͨ[?PlF�Tt`J~��Ѐ��k
0���
F�޽���*p"��`�*�Jႌ�����'ϡ���"�_t ��䟉Ě�߳��O�R�SU�T�V�V*%�;�����pL`Y�����{��_5r�ʑ�j�1al��_]���0m�d�㼱�J<ђ>[hu����g/��\�t��q�D|zLyeg՛PL=��Y^�~φ�E��0+G�h�9vW+�fexm(LeQ3E`nLok�A��R���]�U�L�"�]���68A~K:Q�nO?�Q"8�b��@��1��H*:Q�O{|�Q���X�۹�}}8"1|�P��o�'�ȷ�^�������8��(�?���N�� ��K�Z�}�C܆|�v't�6��">���oH^�� X���߬C<��=����M@V�m<X�,���?Bf\6!��=�����02y���O��(T73�����C�T���,%��M��h�}�<]O��|G���I�{���B�>{��'��h�2�k�<�!���*��H�O�_��rL�����&�L���4e��:�D�,(�o_�}ﬖN{���k����5ȳ9j
�����@>�=��	)��U0h�����m�W�n��\�K�#|�[�Ekͷ�u�����K�D�@�\C�}:2�\{�;C.��~Pj�k4b"�K�>�B��}�/�1%��T��ވ�>�e�Y�to~f�K�`;*z�F�$�O>ً�'\�މz�7&��*���#�v�=�&���Xx~�`;������A[�Fk�`_�d[��q�K��z*��i{��)d8�ȇ 2�֖��F��'w3d�>�_�����u=�6�r
�5�)�_�8��'�k�]}�TE�V��`U��+W�^�d��n��5�o��aI�/�p?��k>�O��<D����y�$[W�4j8)2���5�<����8�W>�P)��Է�`�3e���\����V�V@L��94L��e*��S�X�G)���%:a�0�����Z6���p#0+��o/�dP�c�8aѧ0�J�K�̺�G?*�u����rU�@��7�[X�plŖ�Z�.K���Y�_�o��X+ĭ'h�s����S�\��zK��nQ��:�����xsgY�.	�~Hx��G�W~�Q�d3"�-����T�Jf��#Gxy��, �D��:-�0@J_�5��֊��l�[ʘO"����Ա=2��	����Y�܍ �.���������a�Ka��\��N��~�~�k�����w������i��D�:�ⴱ�^}�U��W�F'6w�>Q=���'�w�#������@�˜�6�˱5�|�@l�.+0��A��[k��A��r��#�y�J��M�9v@D���c�O�-ә�b��2���zDϻ�kJ��\�u�KZ�,)��g�[�������]���4�\�#pW|��h<����A*�����͖!Qg[Y���;W+�{{�����T*_X�7��Ȱ%���g�N����\�]�5٤���l�֢�����-�A��%�ښ+<���ň�X�=7�72 �y�1��ā�~��B>�>��"ͪ	���GS3ʝ�{�h@FN�2y|/��։�.�o)M�";�|a�P����-{��DS�sB��Ug<��0d�l��^U5�^�L��J���ҵ]�S��(����{Z	6c� ��o��u��?�t�k��`94_�0��l㒫�"�;M�F�3d�s�Ǩ<tc�hR�y�%��H 祇x���d>usu�	@�źS/��ߨq������I8���6r�2%���J<Φh��M��Y�tOP+�?'�Bp�����a��
@��I�ЅO���U�ׇӂc?����%��
/�R���<�\�QVd���Ծ7)1�sj�1\��\-���� D`$a�`9ߕ1`���W��T����a���'E>�AE�\$�ܼ��9&r�_�QV��U���3��K��i��t�E�����$���Is���I=�Z�gz����2�_d���F^�e�-Z|?6-xPo[�r�B���^Cc��Q�/��ܴ)����� �x�	P=>���ț`Z���c<M�Cm��_�|��?�'w��9�{Q $�kS������$u�{.�-؛�}a<֭�F��ү��|�8�b���܃'��F�O�9@�{���B���=rU5-�o*���*��|�O<�?Li��66}=d���  ���}������ͷ�$���_�g*��81TE�>賸M�(n2�~��s�Iu��/����4%s
(!�㺭�l��lFM2O�C�ׇ�@>u�|����R������{p��鉌k`?S���`���o������ �ũ����3��U�%ս��n^�v]	ˢ�},W���,zO�ݘ��.L��X{�@\^�o����\s�L��4���R�Xt�ܙ�Kjoj};y�R�z@q���5����
f��9Bk��ʙ�Xn!��ߤ�|$�?z����i��BfBA˸�o#E��ޢ.�L��XVkDڵD4vD��\��$�Y��a�Z�/��ބ�t�b�]XJS�N�i鑡�'{a�s��1�S�2x��Zd랆�6��_��Ag�wҔA��v�����̱Ӿ�-��*MKJ�5OX�4��(����_��G����x���N���O������$�A�A�7�ݶY���	���bN�*��_�?yެV�d����x"-H#��p���OU�F��;@���X�!�*D�*���3��_n���(Pcr^�����|Pz:��"�v% "�8�c�ǆ!W�3���D��do�(Mj��^Hv�m�Q��,����z��^؞Z�o��>%����t�Қg��D�W�.A�*�n]�������;������˃�z(_4Rl�2�;8O>DeY�iR�[�l>8j��c�!op��+�Ga*�2sD+�u�zr~�d7!}x�&cukF�ǣ4�,�H���E�ʉ�)I�OmD�K�to�*(:�e$A�M�B4[0��r�%v���a^4��A�	,)���t�� ^�r������2�b=���f�\}�{�Ϻ(6�w3��m����\O��唦���VZ�,1�?�_p3>�t�8����<��1���+0ր++������<����8����T���6��ca��B_�s�./bv�P2�<�Q�G9���#z�_��Z�FeU~�c���x��'Z���D�Юי�0����I->�]*_X��а����g�#ZRb��TIbd�q�+���f��0f�ʸ�9���c1�Q��������z�j�s� ��oXh�V�Y�vʗ���]p��~�Z��aif��w��Y5��z/��I<CpE�3 mlՑ}����j���]+9g��=n��}drB%e��;P>��q�ؕ��F�!�a�����}�fG�4"�/�0�wé�8!~�����~�U�Ҽq��Iq\���XsX�QK
ʳ��)�ǝe�p�����W����)�"$ӧ��[��B$�t((Bs�{|�Kѵ�F��qM��E�� �R�5�ur6<"���{҇�3*�.H��r�IZ������<2H���<JeLLIy��2t'_1iE�[r�ߎ��z<�`�	�W�\W�2���V*~A⦍|l$$�����-��2�n>�w�xvK^�-nn�ʣ��
���i���R�\�)��#��0��#�n�-r�AX�4�@e�m��(?�$c�HWK�_%��dVb�?�ȫ�2ZUܡsCT�f.�hbh���Q��,9+U����]-��3-�&aQ�'���f��P�/����A���$�)�y	�,K��'0�Z;ʨe���fG1��hy.3s�Wc�'��������t2b���� �fB�?ʄ'�j���@Dd
8U��ex��<�N@�W���;uY�J~�^��F-ױ2�;QUt&U�^;�D`����Tl��Q]�X��>�%r���_�p��.e�l2N�Ŀһ�-��Qv���펁�v�l�ݺ��ss�l�&2d"�Ǜ\�3���~rj��p���.���kK�����?CmȂ�Qʠ�f&���k�ĥse���J��ȏ����*?�V�Ǻ�0nX�K挒�-�	E����l�����N��e*��)��Zx����TQNG
��'k��,Y�(�|Q[Eض�T�͚�=Ԫ}����"��.A�p.�;,�����^����d�ҢpŅfop���u�0_�ItH���� �D�R�w�$�U�_M	��h5�ͧm��1�x*��^t>��\9���c)�U�\w��e��uf�*�t��m��j���ț�mt�P6d�D��?\X\|��ƽ��J��[ˑ�TL,bI�T�9>���68���_*�pUsS����{$#�+n%���XY�=���8;�P{V&앎�&�j�L*)�U@<~+��!����Ƶ��v��F��{.ܛI�T��4����S��h�}XgC����ɞD����Ħ������<b�gF�f*����n��4��J�M�K�� Ľ��jq@|����2��-���&?�� r�9�J���$���q������{=bukј�?\d3��0U���O1�#�b �F�NK/�6��L�5��2	�$+�oŜ d���U�I@q.3�0"��j28��u���q9uIA��9^׻���c M����2�
�M���#\>��S�M�Q:�3*j}�y��ITF��:Հ1Ҝ�]^�a�u�7V~��%��l�`��)��B%
��<a1��K+��v��~m��>��g\��$���+�߬�OĖM��L�M9Cw�����Yj���l��{���ߴ�C��5���@�3%q��C3�l���e
�>0�����͍1��#�3a��+��[�MF��Q,{�!D��7�*'��l�	�j�7��v�&��J�,7X���e�RNJ捇�e�6=����cr0���s����>3��D@�n�8�^>��'G��i��6����'Pp��	9A�l��n�e�0ʰU_��������Et���ֶ�~�C��_�3H�6�Zs�����u�2�2TW�[��C�́ ��|s�0��YT����t^�'I3�]�z}����7Y���76��OO��Xإ�q�'x(��+D@{k1�1�酂@6\4�s��7�I>|D�gzg��w�RH�F�jl��O�X!��2h�6�Q��+-��ݩ&N/.Dỽ+�����uK�b4sT8��{��:&	$��T��-���.�r���g<�:�=tG��MZ�A�n��"f�]P�b�O�i<�j��g�I�N<��R�����G�D5Q��,�j�����OKW�[	XZ��e�*A�"��g��:Kp��!������zz95�Lz�,$Fl�X��cS|�P���V�Po��\�V�TP�`ojՃ}��?؍��犔���<��s!�q��V�K��\�v�a������σ�S�q�C��jx��r��憚�" �;��UiX�1��ƥ!�d��@�K�C��	߽Q�v�{��*�j:�1���&��ֽH�ګv�-x}犞.3\�� ��(��w�`v({���\�C��N�Ԧo��1L�i�ĳ�!�Y��[��6
���\��bux&v�Β�{/�H���#x� ��n
;x;��,ģ��s~^"4�V��I
�Fۀ�1�]�9�Bbl�U��������$C2OD��f����Z�g���sO.�Fx����=	��F�_p��F�Т�Ն!�)�8��8�:}�0�&[��_EH���V��,u:cޕ�^aB0�,O��KE����L��T��{��ڹ�)��Ax	b�U!�_3�l�9�7-����D1�
�?;S�ӮU�$]+���S��W<��"��L%���s��(�W�șQ�Z�\e����'[��So�^�ZKn9��**���>6�`��
g���A��|+ B3��®���� ����:�M�JZ�A���Q�^��1fh�\z��3 �yQE0�=|��3>�4�ag/*�-�k)kP���b�GA�t׿���%��!�b�ژXzx|դ��������#2)ҁ�4�L�ˎE�9'FK�-5oqM�{3A��$�<$�o�=�w��0��_0�>���c��:S���3�'���q�[�T+l��U��{"�Li����m-��&|3�h���r�d/��z����Fv�[TJy���� <VOnv8>���Fz���kى)wM�7j���JҨʽ��&��
+�נݥ>��@9�q�`�ߛ��
jX�<ڝAE.뻐	�Z��]؜?�����5Y��YK�&3��h��A�C1��&w�Wj��ώ�	V(�G/~Pqf��b��(�W�x�!"QqP�XjE��[�u��!��5r�u`��_��]�0�>*���@*������󯏛��_ePr0���C���Ѵ2μ0�qI�bdQ�ր����1�H
���C�r���j;B6Y�����9��������p�]|��;�ggҭ$�*9w a�?4�A��5�M!�yMI�e%��<9n�y Z�̵VH	����is��6p�nY�-�H�V��I������0Y�O��[9�W����2���SF �k��yx���R�j�V�� ����Xa!^s?�ǩ}�����sH��3M`rܩ��Ȯ��׉H\\#\M���i�0�{����͎�?�R �>	��L]����o�7.�Os8wp�UQ��/X4X<Tbsn��9���G���K��'JQ���Z3�_���&c]
�Iח��>�%��]rE�L�3�/�o��<�R�7���EVn�o�o�َ��T�"4�4�y��Z�檧a�߆�M���-����YN�����>ٻ�MA
)�ڏ���D%�E���'��T���D�-����!F��+�`m���<J��PZ�6Kn��L�}�lf8MÔ��ljv�C�:�!�i	OM��k,���؇b*.��{B��Նbd�	� ��B1a�:�Ꭱ'��v�k ԩmmF:L�n���Ok���%���5���-qmW�f�.y<�?��R��[�*\�3�s�U��Z��O(���Q����ۦ�u�q?l���y2#q�Ԛ>��m}Mt0�J'�u-i��$���v;#��?��n�[�Z���>��٫�;G�fCTB�0�%�
���۾Q��c�M��a��1���U�A��3l9���{/�ו�L�g�'�&�_��M�"��e�|u�X����@����OW`)��!�
h�~���>6����C=�+���M�zy=��u }��O(����a�Ճ���G���-��ޯ3Tď�n7Ǽ݆lf��Uڴ�Zs8
��]��$��=]�V�F�4I����4�W;���.P�[3�?�����*[�WW�cA����[2_��$��ǧF�j{��|��j
?d�گ#>���I�)�	� Y��h{�x;�дwDN��,Bȴ�7�>�^�`5�f��݉'�ނ��.�%��x�\
()�=@В58�3�ov��^��o\M��
�]��a��҇q���#�iw���#Ӹ��e_�� �@���{$��U[�GP�{�����?����}9=H��'����	8�FJ�n��B`�"�2�B�?���x-��j �y+,}���ڔ�3�2q;r3��L���p(��2|�R�`��9PF!F���o���=��BM�L�'�������p߈��"��H��?�!}�9=�H���n$rY?�%߀�j��$���S�0��'�,t�U��ܔ�������fٴ*l�˾5�a�Lq�iA�nO}��W���(��y�O�	�Y����(�f8���Z*���k�(�}�O��e���NT]-"���J�ܻ�������f�� �Y���K�����J���3}��Bf�����p_P�T7|���=�-o}psB#	K�؍]D-�aIb��2��ɨE�&K5��\��z�z#,��l�p4�Ĺ��hR��\�F^�I�3%g���+��A9
�������yܮ��8X/��y��k���)�/[!~'������6�l}q���,P`S��ጥ�QIj�k����ǧ��=\)��F�����7�4�������^����K�DDT4�k���v�VS�[xa�I�wU^��X0���%)��v�T�	�-C�9}����"4�l')f���yZIm���!��8��š�;ĹA	NI�˪t�h~�{Ջ�Vq!h��v�0��V��Gp��b?u�Y�ci�F|\[�%7%�r�t��{�Ϫ���2����t��JD�׿�O��/k1�|8^�����X"���c�7������)��>ڮڋBN�T����G�v��"Bʠ1��h���KqG�	|�;Vy%��wy(-p�q��UU���b'Qj�vp��W�����+Β��+�Q�W�y����PK����FrHQ��'��q���B
0��E�ġe1��
������ܫ�I��ΐy�1��j�_7�~vL�ʵ�̭������#�|klht��� ��VB�3IZV ��V�;��ez�^*T? �����~��4d���L~�+��
��(:X#�^�F�=m'��ĸ'}@�+�֩�P3�E=� J+��Z"k*X�6)��]1�tLi�V��~����&���_o�6���
�p����S4��zQr)���j=��Q�T�$$X5 >'�s51s��%,��-�@:�(����:�!4�s?��2� 1��)���?:q)Z���P��u�����"z�
3�����Y
�B��e�Č9���^Ʀ��k��� 	!�rC��"����B�t{�L�cզ��LPm���8V��ӾCq��-�}�����I������IYh��(XA�	����t2��h�Mh�/UjJ��y���S�_����~ 8������C)�k ��i�_/
 �EV����-�TCp�؍*r}K��E���eO0F�ܕ��u�ϐY���g���.W��j��W�7}Q�$i$��#;AQ�[�t��B�)�^b?�|�i�/m����o�2V����qz�ݧ����@������T��ݗ�ʺ�0��;g=.�r�EB�X�'�_�ըzT
3 ��T|���d���Y ��k�#Wt^i�}�6o.Y,�o*ϴ%@�?h�l�E�P���lC+�d����mh��RLK8����x��>L��;���؄����j!�/�,+�����w�O.>�䣬4
AN�+\��Rm��7��7B��ʯ7�G�[�*pG�o�4�<�2 ��ܟ���)bj�;-�-�� 	p)&.h��(V�iE�I�}޳xh�Ϯ����ꌌ5�	���U��-�����%ti:��p2���%�-�K/b�(DH^�2m(vĐyjC�WD�!�9�a�cU]m:k�`��2;S5��ZG��A�X��:�ښz?��{�:�XM�����Z`���@�TJ��}5���aa�}<��l�z~�Zx�L�gԅ/k�9z#
�LUۯj�NϽf�@��J	��y��|5!�ෞoZ�x/�?�`Y�5T�;�؜�*dF`~=�/F��!0��;kW~�;d��h�������T�"�f�ču��[�-��Ʈ~�l�/�G
�\n�����9Y�@�2�"�U)mM}#�ZW�; D�$[�I�#D�ۈ��Z�;!\/����a\�*�K�=Vڀ�?��C���E[��E*�K��[_��_"�F����*�p�$U� ��E�����-�N\��b]����8�Sb����M`�~�r୏u5���?$��{� �����pU"r!��㯋BF{"cӀ*��Z�+$�Q�'� d-��<
.)��s�ʮ!�s�-�=j�M�*�O� �ۑ��,�W�&�&�u��X�ܔP��	��G���a���|������d֍�F�8s��B�\'OI���v'��xўs��u�!�Uw���_���>�?�"�t%���1��C:��(�)0jE���B1l������ͤ({�X���T�rG�8��]������Q49��I����(]`��uF�����EA�1��.��+^���\�a�U��8iFDY�&q�<sy�` ]���uEXF����'�N�ý�7��B)fY�N���F�Tp:K���>q3��+n���cg�[�~�q���v�����dGkXx�дǟ��˰y��zՍ��{:0z\u5�/���c������>�䲖�;���-Ѳn���Vbвjk�v�B�'�p�ޯ�%���Қ���]f.vw�N�icwCj�V��f��{�6�=�%�or��ͽ�f`�g�N���P���>�	�� U���g��@���P����ȷ��I���/�$���>��'q	��;|��J�bMϛ�$Y���F����Hl�:��E#^X�gM��r6�XF`�Q��,I�j3҉���z>�'^�F�/����U���-���0x���T+���D�9q�����x罏U��	��W���%6�kkCy�H_r^�Z�L��u��8�q
;�⒑G���=S8Q�K�ӇD�_��
`$�)K%�N&�d*h��Յ��@��� <6kǎ��.��]D#�	�0�e�xݙ�%�9�;�2�J���M&C�9�Ds���fIk���Dz7��mL�ǡ�29�O�0v=h�� e��O^���D'��t/��Q�+i[,�p9��,� ��9�i�J5$Sj�{�Q�H�62�N�3s�ȿ�K���1�߰��Ͷq����%ދd�%��6�$��EV���T�YP6��	٫�^)��?�jlU�,ZF~�חq��/::�\�^_�fS�+�5TI98��d�J����Ɏ�S�b/	I#����p����D]I���Aھ~՚�M�)]��&?#�b���e
���,g� �n��:��ܳ�%�Y@���5���;�BN���W��,@����
ƽ9ȳ9c��6ƥf9J�d�]r��Q��U�^�d����v�:����IGк�Rh�[���RE�j6Z�0ܵ7�Ό��)�����Z��6i�H�͸�0�SJi#׭y���.|�3Ɲ����B�<d;L��ҊqBm�`1Q���Ҽ�po��{=+8긧�=o)Hm�\���L
�=ѪT�7������7��!���Q���mV�V�biJҤ#��9P����3y��ثr&8��M"I����P��k|�(;pIk��� <Zg;Qד��b�%�d���]u���0<��Pb~I��똥1�R\����J����ʐv����d*y1q��-����(�� �>R�N�wa��G� �?������ݎ8[7�8�z|8���yNQ�|4&F����b�	����%�d{%'Å���ٺ�`H�t}3Er�����t���yډQ�.�,�0�1l+���j%�8(�g�rU��n��8���@�,4����c]�6�ڪ0P�����~����<�B��'�%���s��ᨃa���o��0��=㩍ݰ�N�)<�v��y����d�Ȋ�ᮐ��@��`u��Z����0=�
��+3*�!��iG�%m[N��ۍ�e;?��f��r��wK?+^��)Qk��n(�;�R[SuM'~�ǲ����ۛ/�P�b3��l���5��2�G��uSd��_Ѿ����
.��C�����#:[��[Z��o Ԍ������>��nc;Eb��L�٠L68Vn1 �(�aꍻ���������G�����R�D��y�gY=�W��w���R��`o�0fEb(�T#$x��������	j������^�U_���w���lk���5�s�
�Uy�%7�p��k��ő��tPU�ҊD����W2G;�E��ܞ�-�kaQH����^��B7S]�&�s�N?*u��ݾ��x���W�o�o�O�Y���t�Kт��e����>��"!;>d�mk���	>������n����n�lV�@錧�#��%n]��О�j���I���Fq}����x��W�v�S�h�A��m��ǿ��Еij�k�u�O_�4���N�Y 9��go�.t�W��N��n����-B���A`�1�,�F��/���k��.���%!�t&�p��|�6�����yr��CsQ�Pz�+f�Re�y�,��An����4(e��#M�Wÿ�8���)�m�H�p�e��q�8��ŉ��*���A�� A 7H#��!�{�HX�e>l��$�)�!�uEf��yy��*��)�����Ĭ��uڕ�!(cG��z�0� U������w.�(�:_�{�)�v��2-/�`�J\bGC��':vڕ�N�>KH?j��ۇ�ጭ��x{�3�� \�.�:B��
%�$]cT���$�̃O�1�k�8�8�Tg�T~7E�[�
8�iX[��
Q7�jA�c��A]��/�'�+׻���J�wf#ᓮ[V�Q�~�Kj� Oη��<�^�<��\O4z�a��1I�Ks��B#8��2B�
��/��3vt�C�����|*�Q[�7)�$�v6I�Q)��0�b-p]cF�B���>G
0_L%�\,����hh\��<�3 ^�R�k�"��^�����XGg�'Юj��4QH�O�a�%kH6t�	�����
ߟ���6 f!�^��p��k��2�E�'$K�J��xc+<<�!h����R~���ￗ��	<���S1 �ꢝ��C�� �$x+�޽2��!\�L�>a��7e6�����ӏq���8*�(`M����ץv����X�i�|1y���n+����Q�1x����w�C����V�gB�S�B@�ǥm$�����r0pW\ln>	�W�Ph�:d �ѝ@�R���k��Z}�L�7z9�?v���:?zO`W�IcJ��]�j�Xo=�?ӝ��<Q41�͢G��i���$��^.�0��O�-T�[����+9쨍wb0� D���{/N��y�cG*�g��c��u�����#-u���d`=Sc�u�T3K�C��_�)�r�O�l��'��y�N����  f)6���r���V�6p� ��V�y�+��^x�X��^��;��]9@��C�qg&f�d�.x8��?����� �BZ�]d0cV�I����D�MpB�4N�dB9��� sb+�[��m^���Rຐ�l�)����F\�E�j�w�#Ao��B�W���O2q�?����d�(�4m��V���S~���Cr�/~��?�z�)�ݪ�č_W_��:� 1O)@�Z����%�R3U����q���\C&�s���=�]l����fY�`H����g�퓢@,倁r-X�d�i��c=xY|YڅW9%���<��&���k2h��|M-��9�lgU��%UgKap;C�O����M*�o�I� 'RAs������M�����Gѣ��v�d�Z��M����d�AJ�7�%� a�*�a�e�7�@����O3#���+p�^o4�p���Q�3�ܛ�`��,E!,aR�6���ںOr��	c�)l��Ēc҉��w7:�����I~�ti�'��ġ��l��|�'?��8R����2=�,�7���>���|�!=��!����%&I�5�yu(�W���߆N�/��~����Դp�B\j�"@�J�­E&t�B�{@q~�����X���;'`q����2FA��u^DuD¸A�%g�$L�RH���Kj���ͭqn��gD��H�y*B���@o��d1<��j���h���2�.}�#}�~�=q`��oBD�(E0&�jJ�{f3>����#�tz�o�����l.�s̉�Xd	��Ѝ˞�O܀n����?�ӥP����׸�O����޷Nm�:%�͚d��cp2���ɫ)��"���B�y���ύ~\�d/�YZ�"�B��k'�<꘻���YL�5��������'��B�T�� +�CMa��kB�:���P{�0%ϻ���frKi��~A+�*�	�z��ǌ���o〝.'���u��>�Uh�g�}�<o,*���qT�>����f�b�N���^��~���#��tHwQ>m������ڸ?v�:8=	)\e���g��h��0 �c<Ov�(�	�һ��A������u����_�4f� ������Pӑ��l޽���^�aں�^-%�.,oʦ��1HzHA�@ ����()����@P�N+R���pH����ͭ$9L�o��kW�k�,8L����N����d�qX�/���-E��Lɿm�#Z������S�*d�g.D �D�>�#��b�s�x�з+O�孰�77ǐ�LP./�'^���۔aC���@���s�z�K��u��l*�%�VُB�}q�1PI{}�^|��I�T�=��t�޷�m��[Oចq��\�_���BԝW �Ț�"�:O*ȹx
20��$2�΀��B-���sbE�]�h��?�}UYT��J]'������IF��6����&Ì�-J�&�%z�R!z1�����1���Y�~��.���mf�m�VHR ��9�x?�aR�#	JQ�]M�k";F�����~���vM��m��v��f?6�3��ٲe�!���A�)����1�!��n]��=�o}���|��5 r���X�x%����%wB]#"�#v�,k!�)�ط_�E��[X��fc ���{�NTX;�!� ������;��%���?� ���$*�?��� �"��N�=1szO*�c�3��>��ۉ����&���t�� zsC�=hRU�4@A��r�㯋�"cܶ���=ycȤ��� |MS�׵�j�L��"�QS�ܱ�Yĝ�� ?�+.B��R�S?���"���S}V�h@���R�yq��ëF��U`���{��Q^bJ�m͛e%��o�����Q����^�T��Kv/���3��G���l��)����#h,��A�� �&!�w&�^#�|Q��B�G��������ǌ >b�	J �1��?!k�nӹsC gh)�����G�!�Gl���%]P��T����)����O`q�ù�d�yޘΤ %�;��p�jC{�Y'��}'q�������w�oG^j��vg]P�l��.J�f�{e�j��=Lz{6a�5�ۧn(��d_���A`R��aE�5�.pw������@���$o-�HͲxB�9_By������	���ڢ[�VnE�ijgK�D3�9�YT�G� ���zD�$���icx�+J�
6�p�~;��,�ܴ�s��1��t�p���P�&�$��F�-:|]��	�Z�r��
�|���.�1��H�ܜ6��JlgɁ2pb�P����ǈ�ڗ�i���
�����XX���d���&*�O�"ih���ɋ����d�}��]~�J�ܫG�.�.�;?W��rkV�ҩ�L��0؞�
�?��}���k BR(,0�!�����5�n �<R|���/���z_�]F?��[�D|��@
���a�<e��r���w�'xg|��a��E@IŃ����A�Xoj^��v�r��gA��{�����9k_k�;��s��RY�F�[6��
�Ӱ�X#ۺ����vK]Ky��̤�Uag����eW�*'f&{"l�\�t�y��ۍ��w@T��F�;�	z�y�+�u�{���ypB�� �p�Q��q���`�-"�/Uk ��(� �!o�K�?Zo��m��(��.2��~�ր�F�n�U�8vPy���1C&�E�9G#ꀝbz��|�gH�+���H������%�Z�����37u۠K�|@��-Paq�z	Gr$w���FJ&.ro��rlc��_�w#t��X�����4$a�N�j���AI@�mɟ�6�_J�*��E�Gy�e�;.�3�k<k�}^K0m�_��Vk��o@)�y�)K��J3��)�K;���k)B�Q�������Y0�]���o�)T5h�l�4�X^��ZǱX��I_��ζ� ct��K غ�uOF�^?IIJ�Ы}���7��'�)���R� �gw��pD|P�G���'N=������F4S��]�0�J�/o��V*�lp�V`���\3�6��}����L"LyD��
$��G�PGr�R�K�Pz�٫��A�R*��9$�O�2v(��J|��젓�A�tV_���S%�8 ��а��9�MHr���0�n-�kJ��q8NSxA�R��؞�֨ ��Rۊ�R���i�n/Qnŧ&��Up��dJ���e���>��'�Ή�6v���x�n��^�[jpBg�B�B#���׿��YC��4{�(��s���t1�ge��Ӓ��1�\�UaJ�|�>#��H� ����>@c/�l�3�s�mB����ٖ��0��V
����g%;C�n$;D9�MW�j$L��K@?�E�uܣ���*��Z�bԣ�b�_2��d�Ύ _�Ʃ|n��M�x�[��5Ma��G����Q�&�ү�بk�j.���.	E�2�>���T� I_e�N#V9k S̮p��c*^���*	q(�+*��D3M��� �#�e�%���ރ��]ȿ��Q�΁x��K����a�Y׌��	�rK�Il_����	]*@)4s�±�hA����W!�f����,�-�1ǷX�u�T#��<�&&��X�G�ץъ�⊠�4-�#V��Ϛ����2
*�T�U��5���G���D'��B5nr1��W�'�I���9ęX#������]w&w�����%�XA����,t�w��U���Jxs�k���-UKq�R�ܿ@� �|�:����]���19��T�Z�5��X��G��+��:����m���@y#��qj��D�M��k�����S4ZP(�ߢ4rM��QΙ��&VA�o� X��m'�Z&+���"D1b��i���;���6i��� �wK��STD�ea'O�s��Rx]�$�+IX�+���
ؙi.�=1t�<}\�u�i�(���+
q/	�>�9V�"�f6q,y�a����CS�I?7��WQK-go>��xK5p���҉����b^�xP�V��@��ɥ����neZ��~�3֖���q@(�j��ΉW	Ph�lB��P�,$�g&Yģu(����1�v1BexywL)1���)�����3��߽6f���d��`�����h���`��&Fr6��� ��Q(;2!ُ!��i5u���!�3��+ζf�c~(h�r�Ƕ�tp*N6\��`ӎ�huqN����{����r�U�O񴀽�)�U�� Bd ���rU��$7���� V���8=�4���<�t�oh#�#�^;fqM+Dg
P��%/�j����kaxy�_l�K+�|�忛7����G2Kk�us��,�tj8&8��*�R1ҙZ�+ƕ��5	���R����ouq0�����T*��φg���s'�C�宥��rUd�O�ҁ�K��D&*�Tۘ�ך=���9����H��iFe�>5�+��L�_��T�/O���	���*�+%��C�W�	���	�L�jLz���aT�|���Jh*n}k�%mEɁq����fK��N/��:�3P��p�f�ͩ �5��#AITp�e�e� w2,&�Sh_T��)T�������t�@J������\07r��$�'���������=1[φD}^�m�غ,��	��^��U��W��:?̫�YJ2X��Q�ZYE�o>������2Z�}�{lgLp��M@�Ade��h��n�]{w*!T5߭T%]R�Fƽ0�/��wߥ5>�?��|�r�$T�b��Y^r�9L9��/��c��e* *��Y�<��7���	_Z�3��iOk����vU�L���v�e�:x*3r�Vz�=��ǹJnA+|��l#�-f��׻c6���j!m�ʆA�>Wy�����J�HT�#l=�4�!�;a��6��}y\�ۍ@�D%��Y�~��MG5��	����.c�t���YO�S�\�!��_��y�a`����<+���j�l�<��	����B�%�j��3@JM�)i�p���3v�fc�Y�����XX�,i�B���}6	X�����%�G�(B`H�,m�8�T�gf��Z@�
�_�{oő�Y�L\�Bċ]��`�V����H��|8�3r�����^�i��	C|��䶜����3��#,h"�hMTZמE#Ƌ)N��k�Q��X���w��W�-2�ڠ' ��Ub��rl/=9!jd.H�{�&��{��L���8��x������WU� wMg�����V�$`���pb���Ƴ�Y�َX2�a��y�2�+i$:�پ�~�΃�6�L��5u2�1:�	��v\ NKg�@�|3����cn�O�Z��74��a�{�buW����m+V��� �w6��yf�W!���d����S�VU�@Y�+4�o��&0G9��0��4��=���L���L9���z�D��
!: ��48b�C��^�+&*�S�`�U�F&D;5,2�h|�d��s�+���1��=hc��j��l�t
Ε�.9�t�i�\O<a�W���b�!L-��[5I�w�\.�x����~lU���o�F#�z����*Һ�jD]b$��������n��N�[�;�j���i&Y�ʖ��n72�%���8��ÃrCϠ]�1�#ø����R{���|Y���c��S'uI���p��y|}G(�H8��Q[f���K����ͥr�iq#�jB�_�rU5,a��	���!�����W���R�������_��&u]7�vַj:�:�ȶƪ��\����QI\�2�);L��ŵ�Ҡ��_��-r���ApMG~^Ex��ص�=�Ԁ�����6�fTb�V��XFb���<3s�F��U�(���PJ�Ӿ�~��HoNX�ѧ=_J��\����F�E�A�tVO��i\&�kT��Oϑԧ��Ɔ�X���Wc	�@�dx��뵕o
��LK�ccA5#{�(j9�i� �%D3ۄuHܤ���ؽ>��	Fu�Y��֩����n;Ƚj��3�8BBz��j���\�=�me&���'����`�F���Mn�b�T?�Q�K�C�(8�^��rx� 5�����v��NVh�z��r��}gb�B�A<�ӛ:�ku�����pB��\�ɍeLa�
r�3����d M�H����qOΫ��!ks=.^��c�� ��f6"G����Ns�o*��%��(HN���?
n�@��v2CΣ��i���0z�zT;�2x<K&�/�(�����Q��`�/��8FB���u����?�8�Ks�l��I6�.�d�B�)dn:2��5��,��JAb�]�v�2��+_}�zR9���2.���{J�lb��{���R�����q��P����&@.�՛y�ԆIl.Oc}�%I���
g��R~��A?� ]�%�ĩN XRioKLo���� ?��	#�*�Q��"�k�Q^�j�����g�+���7qH��t7m��������[�Ѕ脋BW���������K4���¼lI2���:�W����n#� ��Ÿ�A�c%�h���4AM�l��+m��50^�-Ay�f�[���G}�~���7���ݺ�-�\*m6ű�h��h��
Ù��yb$�~Q������Ŧ|,t L����7�x�E`��J���Ȋ�X� �/k��,@A�h�m����c��PC<�V��X��P\1��/#~�d�>����P-� ��h� ��E[��H�����Kg����Q����`ӓ��NyAe�8��@�^Pe��0��* �RN���\PZ��a�$U�cJe�}�]te/U�B��d�՜��SԲ|��;�_{�3uп�i�T��̦H��:�i���d�6O�d6���m����>v�3�f��d�J~�s�3�!���æ�S��adP���c[�A.�J�� �E�Ҍ��N�\�6�5iᖋ���8�nV�#�?3y�j)��e�꫸��o*�no��ްm|����?��n��ھ��{�ž=�?O� �J����8*҆�Cu�e^�������&�ˡf��RD���� 6�p�ao3��h��h��!b�WA#�L`٥�	 _(�AfҰ���`alۊ�J�
|�7���Fbs�k%��!j6z�5(�x���7t�K��a�~�|���R34�O��T�Dx(/�W�U�#�L�]����W�[
��!����up��&�V���o���T����A޽���̐�_����˨-%IuZ�s�2M����])���}�@}j�2DC��z�h��Tbj��ڑd�;�f����}�S�,f�2��&$b�k��6/�C� �kZڀ�"c��%]D�6�%qQ�%��L�[�0�Pm�5�Ӓ�D���Y�1�=�1�c�H�a������@�d��s�Yp]`JI7��
�Xt�U:�Ļa~�^�`���Ƒ��9E2NS���Q%�b(� ���Hk��S� �q<��8�Nt���|�W�q��3z�0�K�P�e�v����j�������!� MgG��s�Bʛ�O��.OQ�5#l�S���-i[2fЯ~��81�µKo�M�y�L-�lo�ȥH3v�ڙQ�e�1J�%`� �����'���m�.��`&mTI�Ĵ�	��.2�ڎ'���G�ǭ#b4��0���E�qw�XcA4��F�o�+a2��;���_��ƒ	M�`��Z�gP���)qH�W��l���k̢�T�jéo�I���3� / Rr�h|-����~XG�>Ɩ��(M��a滑hJBM�C��~b��rg����,7���q!�ntf\%vn��P���k�!�V~����xtD2�[����V�ڮ �`y�m��%�]�Ӵzj'���q16��FPw�ۜ���T�|L�� ybO�|N�vJ+@�~yypzٞ(��f�\Cm�/�R1�����TŲ�B"6#��{�v�|f���a�#:��O^I�f�8��$#�����ְ��>�?�FJF���(��O�w30�ږ7�gp���Y��6%�wF�̊��g\��d���y��LW1�ȣ����FP�����<�$�{��ۅO�_|	/qS�eiBה,d5|`���E#3��BS�������蛸|-ᵤ��E$� ۥ%$�i�9�̲�?��oU@�ۂ8^��`U�t��f�n}�������V���݁Nk��V��0���S$0H��,-\�Y�"ə�
��f�fR���_�s�� 1�
^I]�ܘ�p��߃��^���8��W�i}zVc�W>=�"�Li�D����e�4��3P7�t9��;>���:��/^��سU[�C.��u���SH�cI���X��1��:�����Ƭ;/��m�_]�ɱ[M���1���z�H�V���ͰR�sO�nƫ��3M�Z{�qf4^5fGG�n�����*&M�e���s��Ƶ�<��m�rL$�g:�]g�j1�2����j�� ������T�٥k�g]g
e�.u���QȔK?�W��	5"zwdT���Ǔ����i�����:*9�M�ř��I�L����Fyd�9�T�$�$�����BF�X�������Nh�Rߟ����{�X�-`|���-i��A�A�̷v�B+�e�Β"b�-Y�\Rۥa(���\����_��݃���;�{y�Lnd����H� Vk�Y�=�ߵ�����I'Q�N9��%D����K��[ �(U�2�'v�s�RZ4�^�ZЮm�Tl�X�o��o83�3��&�����4�U�f�m5����V�P��7B��Fs�:'�
�8�I
y�;��_Ѵ�Kp$4p�����0Q��Y�VɎ�^��缂P�=T��M������Y�E�M�Q����'|]�����P"�řܡ��t_j�[�ќ���L6]����l�{!�6@��$��o3 ����F@�X~����2�5��L����g��Il0 gDm$\��>�U.��
�u��^F5W��D~�B0��af�/�wP��k*Skt`K+���_?g��]�9��֟�-��ޫ��DgR�09�x�d0�U��X�r��a5��?�Ҵ��Z�Mʦ�hX��?�x��)��tB�F��=�4
�7�&����v�5��r�59�|c�m�ȃ��fd�n. 7�[��:�`tB�'�!@WƳ��b��ё����(��
��Wđ��}��`�'}\KfA/;�x�/t���9�k�9�(�0߲�P����4B��<Blv�k���w��������ʜ��DV%q��@W��@�䈑��]������+�X�AK�V%�i{ڻ/2�)�O�K��+�KG���!m��U.�g�np�ODj��<��Vv����N0�f`��t���q{~X��;���@Th�7ţ5�����Rk�]r��2�����$8�jv
������|9���L��%��4�P��1=>|D3����cQ�	�*7I*D�'+|<�xFO�|�4d[*����YM�1X?�|^�������u�?�j�}��5�G��P� �O�M��td�/"{�9Zgی��'�M�Oq�K�|�d$����$^��*Ȧ���QB���v4��6���ʫ�0>#�w>�![O�Px�!���C��!{�$�A��1|���Ư=g��+nW�'(�5J5r�!q�^>2$̛��=�1o�5p���O_��c�㫬U��%�`^��Hv�*v�}�.�F�%?+Pⷃ�Ta�N's��{cmT��
}A���_��ɧ�L��~_������'cn�J���5$0�ߟ�RK��|�/��}�����=2IO�n��� F�T��m���P�`q:0����bD�9V���O#��k,p�Zˡ�\�l�M ���XNY��MZ�b�^����Q��f2;����_ӎ[f�ӫнN���tI��,�2	��{?^uD���3X��r�ʩ6_V<A��L��R�y|�1P߬����V(�(/���ru����O���g�<�r )�[C��L(֍����k�M�F#fk	;�����'�JH����d���zp������ʪ�Z��Q�.�G�E檄��to�O
��sq��� �y4��.�y&��?������cv�cM�}���9b�	�Vh�¤��N��H�y`]����NQ���"�$am�A�����O�m�Ԉ`ܒ�ZS�HP)����(�`Ǜ��/�S�J��M�{����ǈ��#�~._{�W�D��矃�7�;� ��^,*��7�CC�Q�J�9� ��U+�J-���۹�����x����D��k�s�����h�5�[z'Ħ$l7�s��>M��t'ul?e�����h��Y�b���U���q��Qso��#���1�xS��dL�GGW����6y�R)D����ʣ�Ŝ����d�Wo-*&m��Z���d,5Ϛ*m=�����`<��1�l8�X_�1r��<��]������o��e�c^�$�����	�D�� ���m	�8��GlVD��҂��Ʊ�j�èNl��Oe~$�����Ǹ��Vf�}��O�!<���:���#��x��l����| �\�)��k�5�2���N�}�Deaw�e�lh��I/wϤVB߭D2H���t�y���&F����*��.����:s��a�r)#};�z.���.��آ*6@o�	�V
J1Ā!�N6VV\-m�`��*.�5�R{�I=�.0�e]q9T'�|灨�h|�҄*���OК��T�%���2CP����0R���Z���'��^ �e���>����8�庭�I���!2 ۑ�I�A�hF'D��n�N��ogy-�K��[z"7����o<(C�+�![Q�B�����*,��%��ps��G�O��k�2��l�K��ִ�[hsk����m���2�#�"�K�"ǡ��E~gC�[��n����2�I`�*���,�O���.H�&=b����Տ���|��7��;]�q~�M�ڵ�Ew[y�eI{�����;��Aܯ�;�9{�fw���e�8P$W�e��aT�F�/|:��;N
u��&ŽC���A���W�<�@E>���oq�!񸵋"3����WPb1T������Q��O�ax���>����y`�l�~�6���?Ω��R�0�󚘿��nO�Pd��[������yr0m 8�}.�):a�!+��m�oكP0��"���]�lӺ::q�pe=~���>E@y�q�v��D�&r�>Q�b�/�J�>@Je�����Β�{҅�>V[H]����v����+(�u�!֟����H�;I@�k|�:�=���j���k�u��"��� �8H*�L�v}�;H���U`���)��P�s��Ε:�Ў�b����R�D~��,:�ŧn1s��#T��؏�Gp�O9��ځ��'�����=���C��d-"$P4���L�H}���s_pV	`��!�U��	A�i��3��~����ޠ�a��Vg�O���֦�ii�$d�u�����È=��q�'�
��9n�)e���(!_���>�����6Npծ��I��'�������5�7��$�T�̸Z����\6�]�l�elAx�}��5P�*J*��3]|���o���P!����P�������f�;�G�;�N񒝨Ρ�����D��]�U#_U1�QZ���iU����,Y�9�
/Y����A��S��v��z�DYT3�Mq�xgU�h�b"_pt�	݈	��`!w�9��� ���H��]&s������G��/1�U��	U˰�$y��*�
Q�W�"a��KM��6����f|ζ|�7t�r�S��4�M��1.���XZ3d��寙�0�Gl����W�>��eT��wM�T[+��ꂄ�+O�]-0;�j� U0,�nޟC�ߥ��_��#$��W,�V6_f�|K<�@8��A���j�J���P%+E ���Ff�V�߳"�޲Z��3���%��0��u�hL�2�5���fy��4�E�j�L��Qۄ�[�Ѣ�=5}'�O�)_��Zߵc䩝(g���k%�o��>
t��G��^��vkdJL�0wZD�'��u4�E��ב$K���;xL�A��m���g|C���vN�IB��Z��"��O	`�"���
W{����d�P�_���Ǿ�$�%���'T<��xP�P�}RqF�E��}�2����T19���ٻ��{�p!Ï���hר�D4�Ջ��kW��_�Ҹs����[���A��;��\*�Vu+y�K�W��6N%����p8�.���g|�pq��'��� �!h0�zW�o�-��j��w���ו����ld�!���߰��=Ù2�}���w����#��N����g3���7 �9���U#<��6c�<D�[�/���nC�'�i���Ib5�zn�)��B7�1?6�I�Bh{�EOFe�'��|g��i)�S���tj{0F�]=@�V�mu�Dh\o����O���n��J�P��#��ʅ*QC��I8�s��?���_�s2`��VM���v�0���7��v�|��|���T�/��t	f����-� �s��}E.ĸ6nc��n@�II�|;P�i��^��λ=r��o{rZ�*���=�t��;%̱����UW��J���[����A�P�O�7���l ��5S�v�g�&�Zj��M[��.�����Q�fp?�����E��{�Wi�QI���8-�6�X�}y�d�>��=�a�c l�.A�E��9zN���uF�Ν� ���9��Ɩ3�r4c���@k>�^�V��1�{ߛ�$�D��6��������"�mU�T\!n�m�xu"RTd��}[��b}�����(��G�'F�P�/�U(dȽ�����Z|m!��0=H�;��	��%@�ԥ���]B���r�� ����l�\�H�3��~ɛ�}h��;r� q4�Z��Y$���N^�d�,P��O>��>=����ۀ.�j�-�R/n��B-5@�`��u	TL�p�,� ���/:WIS_W�#�OL�ݻ���ӎ>��$�iK�C_�����Y1�Ze�"����jj).�����B�PW|��7O�͝���͠�uiv�:�����(�|q`h:�;OزV�Y�w�}��G�ۍ���E�����O�ٌ���Aq#��D��2�#�@s����Axc,WMꤞ/26�H����s�=�����䥷|����<3G��?��� J�S0eȤC�����y`����䎤0��po�KY Di����s)	�j_����=mDӱ!��u�dH�M���3e��ތ�k��~����˯�_ų1$1��|��������l�d�>����F�|��A�?;�mN�'�*��Mg��s�������G�
_tsHp-��?^ކ��ԶY�\ ��K��{�!�����\2��]b�z0:�6��k���|wU��uU~��>�S�{��<�����4_h,Ez*���>ҕ]��mքQ����j,#/��8�F7g���_\�L�
�G��:{��3QOl�0-�� lT�f�yb����3Y'��{*�	�F[>�;���������@��j�PK�M��,���� �!i�?��0LBZEE������P���:�ﺚT�]��V����&;98��q����|�N֦_�6���OzV�,�i�U�:��fz2�VkEJ��Nc+H&1�Rxb*ƿfو��.,C���� �ݼ���?
]�_W����yw���y����������ꤼ1�U�͕}0Z���U���w���S���z26�X}������)%�+uZ?>�]� ��^�a�β�I�6�R2�'�~�%%�����`�1�/a5s�����<�����b�L�5T%4�[\эoh�I�i�$��1&g��ᶐ\���3���U�>����z�p=i1P]�z�M�(-�x5����U���l�IR��Wƹ׃�-;/s����#��I�/0����+Z>�a l���2G��a#V��ZQ�	�^,��nH��Dgz`�s��,�1=W<���P�O,��T���?��)���k��3 Wjq�0�60�U�^꺟��_| ���/�J}�1$��o���b�骭��_��,�N�<�NL��t^��@��V�������R��Ԇohg�h�T��h5b��rj_�/!v�[�s�m��W{��84�Q��Pwh����
�P�)�=���L����9�&���sd�n;ǑU	X��DP��V�-�RG� �*��2-������`2I�吏QzR��p����ˬZ�.�~G��Kq�c�^��f[���9V���bLMGG,��yr7MgO@��g�s��궋�-�eX���yp��oz���o��@���?r�F��F����-�0O/�Z��3�8���G9�F�J�M�&�[^\s����P _a+q���P���C��b�4[�$(�Hp�:,�7�߮U���P�d���8�'4��;{O��q���CJ�e/�@A:�b��xL�����z�6��4���r�wT��� -��5�����P]w�h�7jl�=y/���@��z��N |9fE$�QUC-
XG�7���;
�55�8��β�By9��	�*ꛩ����2t�b<j/�C����M��о!H5��"� ��p�F��ŏ�R�%�%'�	�@jڤ���%PU�x^`�s�]pzG)-t�$6�e��Z3 ��JTő~�����_���Τ�C���H�3�S�����^�nDI�m=}��9E���?Q���I,�-����L2<<'�� 3����]{(ݘv�U��V�с�a��9�X*ܓ1��nP��A#���<�1.���,�A�I]��=���?����`����m�t6G;�n����5���}Q[�O��ѯ�S5GD#�n+���z7UJ������I�"��Z���r����G1��Dz���,�<�_���1 A��-Y�B�v7|Q��i�c�G���)�|�ęh��9��6'3�
��;pN�R�0\�r���p��^�Q�T�R� 6����C~�*6�3��Փ.�p��r���t9!U(4����}�R>���.��)qNȖ&�М��`i�kp�#'.��.UD�WF��{�.6=*�w����
�|�><��s�*HYFd�rC���2��n�B�1������z�������������O?�Bxj�$2����8XY��`�{�F�����%�DF=P>��O@�C��"`԰C᡿+�[��)b�<ݦ�a�6�Cވ�k� ���E%�(<%�R)��6����[���u���b�
�����w�e�>M�Y�>Q�͆��;"6�c�yh�3ؼ�
�0�:������e�=�A���Vqo��F��A��q�bQJt�%�V����[����}�����)��X޾��	���r`y��z�pvZ'T�h�)ه���M�h>Ɲ�XC�"�fG(y	�9?��"�3��p?,����hGۣ�v�<�`�3�3ƹ���Xp1��8&RqY)���׉*ϐ��~Ҵ��o����sFB���^�{�f!�a�r��$B ��#"d@3����ɧɹ�D*1������RiC[�"i�LR���OĬI�_���/�����]�����B���̲���x�fT�C���"�ZQk�Do����2�Ӕ>F�U�+�W~���Lj�r�.G���1���&�Ɗ,�]��������AH�&� �'6,�=jWI{�i��
r ���Mugu`��e #���7���l�ř�=��]m��O�֨�YK��`x��W����*bD.RL��W�V����L��f;�
�ً�A�ݓ�n3<p�k�	�zs��xg4��ͷ�H_�7`"��2Y7x�Y������+]��G�|��b������`�;z����+�Rcy��ysTb����(�o����/#��i�,�v)�A bB��n@�e�h��Q]�_�����؀I)Q��V�4�U��V�-?O<� �V���?�q����M1�j�e,�����(���inը'��6I���t�5�J�Y�#�7�~}r���lT�١�
�M�?��E�u����CLO�ҁ���.�Wu"���Z$��'O��/���u%�Js�Q�|`s���nl�K����h�?�i�Tx��e/>p��4V�Hn�NQ��O3�I�� ��@PӢ�����>��ǅ����	��R5˫�o��a�}�v����K�c=׮I�uֵ��@�b{���bl�'���Ik��8~n.̩� ��R��g))��ZyJ�W8��a�Mv߾{���oEk�;����>e硴��5�D$�0g|ʒ;��&���|����2�ǭ��h�yǀt$�2��7�5'��Q�����N9�lٯ浸eV�Ct
�R���yL�l2z�jۘ����߱ߘ�|1 e	�)@Yl�ŗ���x(l�d�H���� [�]�����Q��sP���MJ�/�hT$��5H���..��C �~�t�z��|i0Ͳ�	�pX)�Qhj�_����|����65�F+���o&���<��\�b�t ��v=�T1(
��h�������
�<V�Cjp��NY,������H�:B�)��H�R��o�ү��[�cD?�; ����-U���+h� �'���$��	=~�˱��Q����bP�h!z
��?n��V�;9�����Wn�6[�]
��Z�^��� �x,I<�O?�Tf���@������0hp�֊��99�3��6��VKK�Պ`S��餿W�%+��z0Q�X��gk�\s���H�ͧϡ����%���UȆU�K��!n;�o�_�P���P������l����
M��V!�Y��Wb\���LK��Y��ľh-�Y=�6Ji���<򇏠�$x�2�	��sQ���#0c��W�rF�
 Xyy��p�J���������ҟ�&̛��ˬ$��<]7̖�wf �b>SG0�jH"8gm 6��f��d�d���#^��^���RRI��3�h ���ǤQ!�H�9?ۘ�Jd�#�nPBPC<˲m
�ݫ�D61Ǥ_��!.Nk#%���I��S����`K(��&��
pc�o���W���to�A:��f�!�у�� 0a�Z�j��g���g�m��f*UpL;�ڌf�X[״���+�|:�l�v.�K�l�L�4Z �c��.�D -b��m��g3����-����X4�8Ns3{���;�n����৻T穻x�%o�ҽ��KC��4�=L�0�F���������,Z|�J�/��3�%���Cek��]��D��3hiNGDO=d����6�Ǵ�^�Rv��_>ZK�4�E��6�݈#����SA�NNG&�%��"����^�ΚZ��q	�W����-鮞3ӎJ����3�5$p}{��g�Q�����f!U��Cv�����χ^S�Fy�;/?!+2�S=tr����ە�&]�����;q�ld�Gő���c��#']��C���/��
&x���[R
J����<���D���hOPipP�om4�0��5������S�@}�A9FML
*?m��r�Z�Jn�^c~u��؄�H�ѫ<|�V�*H�&�`�TliW2t��S	����x��=c
��³�q�7���E/�Ļu����,�Z� ��A��Q�������>�o��_�0��*�:�Lwh
v���}�E4x��lT��8�\� �Z؇��`�[F.D��|��-�ſ�?�(BK^d�WZ�m.�b�P+�_?:�c���4�eo/�gx�L#A����D��$���Jj�ߞ��UB�1�$��4��x��˧ޓ`��*�/�����3g F��A)���xs�`��ͽ�@Vi�8"f�6�0��wE0:B��o����]���Ho�
~ħ��i�_U��6�8��?mcnK�h���!c|� ���E�*w�1�pl�1�ѿ��fk�!HU\�	t��$^Y?���2r�7��Ƨ��z�*��LzQu{��J� �w=/` l�Mx�^^n��'/�T)���@o�Зv]#;��|���X�v��F"C����\� p�$yѲ���9fjK�M�5��(dq�^��<M��&Q���r�YiY~�䊄�o�"k�+y8���@�?,Ģ���P������8ԆN����Xv��?�I�p4']bYg��n=/U�،%qV���ˮ�W �O�%R�vPH�%VT��yH��ם�270�5r�v]�N��2CA�)Tjԛ|�>!^w$'Ҭ4;-�n�r|5� ��>�k���:����Vyn�̈e?�Cs�$��+���-� x8�#J�!P��ԉ8��;	�=�m�V���E_�P������t��v<G�L���߅;� �4�$W��2[�i�T�qyt ��!p�p\MБ��B�����(+#�p��$��u��_D���٨W[i�lҐ��FW���3,�k�&����d7���_"�|��ڙ��R�h/V]�g!�0�����E���0��K�ݒ}���]�:������#z��s�Ņf����(C����ހyl���;3P#:r��]6�蔻J1��MY��,%Ϡ�v5�3m	�%'�����-9��`���h��PG=Z�����q_&!��N�.B�@��L�P����F�x��y\�x��V�aawRK���n���Y�������P~ȅ��^�6q������k�.�Z	բW�,�k0���`|Bk�ǧ<��JO/S����z`H�,��p�+��o�<Vוh;2��A���3g��������PY 	sg2�+�`��@�/�o��x^:6W�z�6};sZݣ��ߑ�VdT�F�����n��	�U��C�1E���o�s�P亀&�79t�����ǃ"�K[#VG�n4�Z��_�y��/�{q�??
�5������������J���{�獴�\Em7Ƕ@P	?/���a+���bD��􈨷�ŭ;��D�eҜN�6��dY1��hQn-X��fƽ��v���(�9"�)�@iG��������T­�ک���r��K�JOQ9���)�<x�X���N�bY�͎�|S~���iN����!nj�]�\-���k���Q�V� umM�Cs�&��V�C�����@t��H��]R�����D�T!سbvx��������ǻD���l~�ʹ�}��*���?	��Q�&�#4>[�,�;�786BW�|a��ޥ��dߌ;Rݱql�Ã�9��V�4�����O�(Y7f�*^�9W&�'�;��0��m:�Ws��'���s�������)ܢ�<0�wC���mbD�����z����/t�k��LV;�띏��G���#���_3t�aE��ȳ2sU��,��G.��F����T|HJ����/M�����V��JmI�jH�_��7&P*~�6�4����z�����������+�;Ō��
\�L!NEx���X=ڮԉ�s�pw>j�l��;��x:��"E�r�ag%M����]`~��# :��7��Yy�����娠e��]��ף�ڸ���yDp�<t���{5�ޓ��۹�)�&Fm38Y{��
�������U�X�)Uvq9��L��.(�Dy��k�(];'9�:L|�I��[���U^�@�:���'�j�󀩄pv6��}�a�u��䵺6KpO�1B����?QT=�ި��͑�B�.��
F�\��G3�Lt��j���ldY%�/K����gi�J�N��ߧ%�*�3����#���������₧�������*0d�ѝ��_Ϋ�������R�<�W� ��$ԓ5�E�)vqk�g���)��0��v[�!Q�(��L�E�4�� �sn��@i~!D۩-^�C/sq�e*�~2��9���A�4Ҳ�+�mt�W�Y/F�u�W��A
i_	��3v����؆��;���7�2rm}$^<?�QN|a�������(\V�J��r��Z\�K�a�Դ0�ꟕ4c�7����f�+�a�z��P�k������gn�"�a��EY��\�"s���iLV�c��r���m����������5�hP�`a']E؀ g]ó���9/<�#�����z�u�4�d3�} ��:�$)���``�=��!;LS&�Ե���p�����0 D
��z��.�
��]F�%c�JG�Mݼ!�hv��Gw��%�E�g 1,����8�S��G��XM߰�S��s��|CQ���H��G��9�=UOh�4S7Zue�C�z�:5�2����1�"�N@��q�0�]�t�',����.K��� @��2�Ώ�iz�#5���M�cD�fq#�^]]N��a�X�1�޲��λ��9J�B�K��!->��c򿂽5��N�p��Gf���ʵ�3�`􂈚�w�7ߪ@nռ��ı@bs^��XDg�v��f �Od�#Udđ��x���0��U$����(vC�`��Y,�\�kKPAސI��W����Kr5�C\'��v���W�%�fN4��:�8�O���&Oqv��B�5���БZH A>B���X�ֈ����$.�pa:��MQ�KXś!��eM�)[���+3�!�z�:�Ev=�_�^�Ai�*�@l���y�@ƨ�8���z�y�� �h��D�oi����Q�s��QJ;�D��>1s
WB��&[�Xf���	m{[ƥy���Z�"�S���zM�yJ=C�آ��{������%��j5������d��]�Ю�U��Z�$b�
�����k��@�5��� �`5(A��c��z䍻��j4Y�����㈴b����0��^�4e�[(��4I 4��j���0⁉�S{b�����4���6{
KGx�'�5�2��OԠ2�K���^#D��ǹU�v 8ͦ�d�;%�HbG������!���<�	.XL闡�̭���wm-{�U�LN�`�h;��Qx��^�����9ȅg��N�P�����!)���&-ߤ,俉��ݥ(Uʏ+F7�a����Dp�����P�Hv|ӭ�h��w���-�����R�_�C���Ií(��2%��[���H�M������F��_����%�2L�f�b#���A�����x������s����S�'�%V�N�J}�iG)#�I�5�@|�<��0;BBd9�/���ӷ[&���\��/BO�; �c^=��^����ެy�X��"䮴e���z��N<)%e轃}��紭|P �A8�u� ���0V�N��w�_�|;� {�����sj��ψ%t�{ }o��G0�HB5u���{D�f����s�#{s5��a�|�cbR>�YF
`˜u��2 8�,�zg��/5��/�g�����8=>ɗ���~����~/��x�x���_̜� �^�b��Y�A���p��5�Я�b�P�w�[k����z�tu%a���X��� !��Df'Q�'���:%���Q��aW@S^��������.�^�j�"�#���D���"w�Jʻ�k��B6�e��[�6H�tD���I;���8x��!��(��&Ka�s*a��|٭%^Y�Gێ�����P#���8+��:��=������*�h��Krڸ����9��r��7����UO�]-��'I$c2�QⰘ�=o��1��E6g�C�j��Ҷ�!�|l����;'��	+�z_C���:1������<�3�4�Kf�N{�^'_������NR�L��f��!��^�<����!�mn��&%bf�6�0�����H�`�t9�!���Lڽ��_����_�*�U*UF�v�y�Fܚ�J'_��?��(6��a[�����w�p� 	osA�YSK	���ċ�Ϙ��^^��wiq%L�[1@�5yX�ς�b��-�_U��<
���^����㞤M�aHad|�h�Ó+ ����X1Dx�~K���:s�T���w@aF�q@>6-��(��'���I�E�4;���z���(8,s�@фj�k�Y�-Q�GE��W6�>Hڜ��mQ��)�c�#B|G�MMb��"rs���w.�4�Mp��E'�UhdƳW�Cp�J�EV�)��/.���'�:�/�q�/9 xO���ӄ&���W�� ��e'��L�C�^���ɶ��<z�vM
f�,��� C�S��1P`����<�GC�a5?�BU,D&@@Sq��w!�>��/�yy-�dd�����	.������Ժ`_L[-ũE^W�b��R;�z����=�[� ��L7H��\�t�h_��w�kB	�&2���l`&a®�^�e�kI��v�����'6��'����6����&�L��������|����a���_���?�����&�VU)ݎ�kV'Y��ҳ��pg$"���;w��J�'��zuo^��3���`Ba�oP��We�np�s�4��^��L%&�G�!�h��yF������7�����6c�p�Q�m��y�E���, �Q�vmq&���6����b3p�=�B���}l������d+�Iug2�~�
�����%sM� {4:��ޚ*�A����4���.9c�*/����4L�w��a>�Z�cd�S�p�o�Q�C�nf���mv�]5��Xݩ���"2������O��%�K�K�O�K��1:�nHh2�K�iJ�/I%_ޫ��W*�<�
�F�u#�ɯ��Z �� .*����5t��=�z4o����ʾo��D�p����F��Zd�9���8�oЃ��s�g�.v���rėɓe��Ϝ����ߺ��JO8I�/ )vM�0!^+���|u��&�6h�{./�sL�7��7P�g�bV~���z���W<Q|�}:�O��ȹ�&�g���������4"ҷ�a)(y��#l&�j��!�Oq���YI��W��Sk�#>��P�NƐs��B�t2�M��梕
 �.�E�h'&Q��5�`Z�;�'�FJ�.�R!��n�fo��D���/t\�˵O^z� ��+�9`^^�UyCB"z�f.�l�����V�B����
k�{�\�c�.į�?q���i��
�Y�,��_�e:b|J��i��I�n���	�A��|� �&GG������! ϰ	��S4�S�����jv�����,u�L|.�"�X%�Ԅm`�;Ro��a��x���Ȑ�c*6�W��kR�<y� ��_�v�w�0 �w���r��'cMoU#��P��"��P�<��r}�{k�#�p�kQᓹީ�}�����9E��z��TPeGY����t��-I9!(�����&��Љ�:���4?�DhnJ��Z(}C|�˾��E��0���6N\ā
i`����K�K�j�n�����_�>q�L�Lp��2�.o�bN[����N��X�d�����#Nc/���K�oBy�-����Đpѩ��R��
�sgIx
A�TNkw���	;���xd��=!\�k����=�Eb�H����h>�.�拆���?US(����e�Z�w��iC���g:z�#�����>�4��	��A���������d���>���B��4[�D�
���?�n�iH8둻;Ie�1f�s���o;X7D���P��!���<+'ޯCH�\c߶��V$`���j9�31��㞝:�}�Y��PuAe!�D���T�9�ڲ��x�9�vW�ŉQ��-+vQ..zcjq�Б���Q  �w���(-׃:�^�󬑏�q��nx���v�2���k����r O��h*2����aS�K��q�vr1~��O;��@�I���qw�8�>*y�7+L�E�#�K\v�(rL^�h���Ne=��E�\�O����)%A��ɿ��TA;^����m��8�vt��줴��"j(�K�����JV�zfa���Rk[�I����m�9܆=�gZxH��N�� =�ɘ��h��0�
�qb���ט^�K�t\�԰ ����Ê��Ú� ���Pr^i���0��r)�23�B �֔Xi7�KTh��$�:�84	Wq<|��)�e6�G�˫ �L��B�d?>F��jk��ê��ަ�7��p걻�h&�`G~��X�.����dS½��<;G��s��f�X�� �j�z�N������	�_'ɚp?]��Z�,����[��L0@��[��z ��l��� X¶d}J�&1ѯ���k7{��I�Q_38����:1p5L�	�:|�ܱ��<���L�^�9���q
þ�����x�r��r��{+��2��[Gn���gɏ~h��>��jdX�޺նS�*KGH�푁���Ģ�RW�JY/�>-� a�� M�ӎ�Y�"�K�##4~R}vͺQ�I��vD�F}%@w�_�I+x�?�VX���n>#,QQ�	/T�4�~���.T����-��?�O��7��W&{BU���4�86�͛�ȟ���2^&�Q3��A4$��-���fJ�NB��\{�5������O��_�p���L3r;�MtӔQ-}�G-�nV{���̫�v���j-2y�^�(�}�E�yo�����U�������I8B�*��>f����T��@����Z/���M��,����߈��8�����P5���l�l�WR��h�y���T�/�����u�5�n�Q�ꉳ�y���@A�Ud;�� �����p��}L���R��Y{ $��6�p{�=X66���=����Ѽ���C����XC�p��?��c�kV�]�i�2�x�Q�~e$3o����N�ʘ�'�.^�F�>0 ?wE�QT�&n������\���"Q�O$�����/�Oq��䒸��/�� Q�p�'���8��<�p����gO�!p��������e�������͵cC/����<�$4gAN��������LJ�%H�L�8�xJzpf�4D�����/�����[�'�.����k�⨬��GU��6���η�l�Bd�C�3P+R���o�u�k蜃�-�#��\\�Ƥ2K6���Y�䖌P�ܬ����CB��A-��_��T2^仙���� [��
M����.�y�`i� �G?`򟟠�s؟�P�0AUA�� ���X&�(YC��(�� �籑d,�#@����I��"���{�>�ϛK��0KZ�N^D<8��?�3�^~�k�R��K�I�(jmsF������ٶ`�VZ����҂*�Ϯ�aww䅸��\����im �{�fZf�w:�N�i��[X�{4ewLK�o+��nٮľ���E�3�]��.M\�b�?d) �$c��vTV�&jG�|��O��|z���p]�1�M(�����?��o��]g}�a�2Ee�>���>Wؤ�Pה����d&"A�Ql�� sT.���S~$�yfc��eH8��2{ti{��0n�!��P˥lhR-l�}e�ˈ��#�"������]o��"�]�{�2�S�IBr��.�Qw=��[
���]5�]pP�&{#i��M���w���^n��u���6����>L�Ŏ��U�j���͒G���٢�����\�RX�.5\ A�4q�4jnӪ�['`
N�w[�`N�[[M�9��Qp�����3��	�C�����q��ư�kD���8
�W�`/��z�%R�P2�>:�+Ğ�_v	�T��O�ז��h%�YF�8��,oޟ�)��:��|ܱ�W�Z�N���`�y{#eBP��ɑz>l���.
t��9#���ڡ�ɂ(# M�S�
�R�_ �6܁�A���m�7��s��+��(mA���y�[���V6��|9_�iw�p �x^J�1HN����Hzf4H��H�������AҖ�]�`��R=���;P%gh�Nm#��,���CD<s+��h	��>�<W?
1h��^��� ���.%D2��Ɇ�9���Sޞ��[���4��W�Zq��<��4�ˊ��L�^a6����Ϝ ,�k-�V1�3l����0��^���GZ���Ӈ��C�&������/%�[�h�G{M�69N��<�)��e��n�-��Ig^|����C%����}����dT����c�׸�N�N
��/�PQa��ɿi��:���Q��yD��>.g�Q�@ԹV�Ⱥ�A��#�8��o�O���m*�ݫZm���C��氺��|@����|��z��S��0Y��A~mt�mh��n�S��_w�4��`�F���j���,�>�4U2
ڼ�b���0�o��m���q5F�%^���s�Q�!�_N���+�)�U�7k��W�/�1u7���u�k��%�#�E'��.N
7ڣ��<k>ٷs޹���)F�����DxGH�ُ.�x:`1pU��� 22�(���B��j��G���;�aWe2���k������-��T؅����.�[�{��c�<b�u�ZP�Bz��U��`O���!bCF0f�B�����L������"��<z������/>E�e�� ��q�E���~�/�6��(��{uc�ZoZ�Z�Ծ4��-���`�����E�^������T�@�$�hĶg�Nvy��q���*��b%X�oǃda��8J�lz�T����n�x�~����e��P�00w"�$���TN���gq_k�Mo���rR:�G} ��<b������.u�8:<nqa���r�Y⫒��oO�fvyN�&կd�sS���atO�E�9��I�m�h!�f���s�_r�A��J���&'�D��m����W�m��Z?�\J6� ���P�G���6��\���^���rD�8� +���p���[;a�ބ�36�k���j��k�����5ܵKn���~�@�h��6�S��t�q 8Yk]{���>���kS�g����ȷ��cG#bo��i��[��yy�}|H8������Ȅ}�K�Gdbx�k��;`��R�<Kh����!�|�,����em��Cw���˙!ik�ȵ�,�o���e�lc~^)*vrև���;�¡%��"���S]оh*f�y�Ō.�@�	�
���cF���Q���a�!��?�>e���/?l�.p�>���8_�A���0��c��[6'o2AO�����@�olP�>��3|�hD2=��e�}��#^��_WH�U�&�}�6�L��I��жo���w�������-�ҭ9-W��ԝ@X�𛶅����B�it,m��s��L�H-2�5��J�a��j?�����M�$w�Tt�fw�r�[v �@�*t�J?�&e�v�G�"�WZX��m���4?3��O��3��T_�")QxB�T���p�^
�_��:΀s�S��r���&p	���S*,���4wu�Aq/���Dw,�/��SƮ��*����=�pl��.�$����N�&�Ej��X�Y<+�$<�w�7'T�:�7��h�u;�>��P��0�0�"��8FtԈQ��C_���e��t{'��j��H�[���L�kp��d)��[��J�".|d+�����X>@�s���;(�
EM�Yf=mD��̺T�	�4$L�l�e�A|�����7�r
d�F =���v܄u���)O��-��;��NY�K2hp�_y��v$�w�*����wD���4�AJ�DB7����2:�������9?�+��G((�Z���>[uh���h��Q^)�L���q8����be��EL�@o�6��{J8�L"jk
#n�+����YϾɘ��<&�$ 3�����r$L}@�SEb���
%bb�A�<���3�$Q/bzO>�x%�iWZ3��4��Y�S5����Y�!d$�Y	�?Li�aB�jƎW�NS%�* nP�G
>�|�\{%��,�0�?R�@��2��Q����Y�@L$�Q����~_gcZop�❁��_����ّ�[^^d fG�rB��e"þ[�w�<8	ew1�@E�>}I�asMx��E9��fW�8�����q���5�o���Be9��p�?�"9==�=N��c�1،M	�ڳB�[Ɯf#rֵo����q�yCr*���G'��ș�����KR��A��t���'��+�iG��Az%tv;9�����A�|y���F�$�@ (<��vy"�
��E��~����m���0�����@8�����p�u�wOhe�"���_�{��u
,�.,��	ɥ:��7J��d>N���ި�KK�M���cIylkMy�D����Y��1m,<ݺ�D�~G�٢T�˸��!v��&�>���7�P��'����njn_����y��y��X$���
�6�����W�ٟ�B{��L󭥐Yqlɓp.�(ώz"����_,�p�肄�ݜ!�K9A�� N���6��C�D�:H ��Ǥ;�;�0):ZW���K������	L:O�I��/<�}pP@!}�3� V*7�&�0H��%Em�)��4���\WP�yg�Y1@�a[TEW@�m"�(�x:Qr�Y�����_Pj y�����w�����<�U
h��fߧv��WJ������Xsk�UI��aI�6�+;�'������{p��)�XXJ#����d�m��W fa�Vb�F�Z+}DB �O���,�����T1�,=�D���S!����;��|B��ͱ��б������׎ق�L?H̆쥁���W:�H�n��6Zܠ,i3�.hT#��>[*�@��f�l�c,1.��Ⱖ��P�XI�5P��n�MԘg�{�k��,,m�Δ��A��4
~��O����C����n�db�D��HV��'`�&ȣ&[H� �&�M<s���@���{_'����+W�j~��`�w��6���VNUC������~�v"�Ρ~���^#�?bP*UC�}H��k��G�BM<��ȅ��z�T�`�#��N��h4�yw��V�|�x�c�4�C��~�$��xd�������e�*�x<�=n�Y�H���f�I��hy�f��Faۻ"�|��v~�h%oz��9��B����̄���hB�����_\�3ٯ�'̫�D�@2+X�J�եV��0��ŲW�o1���d�l�͡[p��ȹ�K'���|:�<�]�A�3k����,hF�'�->�Y�߿V�����g�M�)�%uVzUU�Y���}�����z��N�!3�Z�.M
� :B+�E	���$b�0&�����P�i�fH�o+9�;��UbjU�q%�AX�Ϊ$}9@slN��%{/����������.�,�����4��o�P�7}껯cwl,���$N�?���V�l���x�� ��M��>�*A`Z=k�TBp�9D4���@e^�%�
��n�r��`מBΘB���w��bڹCe�guv0�Rޱ����KN���3BQ�״9h5!�|wG���^��=z"�Myv.0vǸ�iT��K���<��9Pn������F���k�콁�+��U*B�=u~�>��L��^��@���տ���@�T�����R�^Е{��Yq[s��h���j$��tO�Ȁ��H?�����m���pul�,�
B�X_W�ON�ˈ�5�8����Fj
��-��.$�N��>��x[l��Z�_@� � G��s�@�g���dy�)���H:zR$��H`-�U�Z�m�K?������uk�,7 �;0U��I$<H*A��	F��~���4��_�<;'`"��	GS�rvT��T�6���x�}@Cp�K,�vԜ1�Vo�5-� ���j�آ���y��'ex/36�6��b��������H�f���5ϲ���� "m��6j�.����y�����o�Q�(��~��Pt�u&���Q	|��
��B�X���"���t�Ff�@`���x��!H=�BR��� �pL@�t^�Ur�D[��w���w�+�m>]�tٯ
���;Q&ꨟ�G��v�X�G�r�޾�h6�끵Y��ds]lVB�΋J�~?��_Bh�S����٠���Vzr��/.����KC�"��2߇{PHI_���.>u����6��&-6��>`{���ɳ�.s������h����_�RA�O�TƜtf�m���*�*?7�py�E5�Q#�����I3���5����,=>$�#�I�I��9�f;�����WuNS���'��s�%�'����8#]2|vB�N��u��Y�J>��67�"����#1�<�C��/�
��y�G���$	6C*��´c��cu[țfx�Z2"�o�2ϧ�+�����4�w�_�e��N��]�%͔�t �IF��G��EO��lJw�~���aB�r��8+���r�Fh�E�|��:B���L5¾�[�V44�����F��dNi����Ş2�Б��{��"R��9�L�l�k4=�M��R���II��;�'zQ���=g�ZX~�w���hA  ��a2G:��G�� �E��El�+81����rr ��p��fJDե���4}���ˇ���s��EwB�a�Y4B�5?QO!����:h����i��K��U��e������M�$!\g�����l�����$v��kd�P±&���]]>�VU�=n��Cc��T��;i� i{y=L�k&�6���>_�.Y�q�$�F�u�t��˽HJ���s��P�UQ?��Y�l�9(�s $�瑕P�%���RUS�����$z\�[e���y�d�^|o[b�����7�E�i����[��?S�
E_�erYB�V"#��l���~e�?�[c�^VM?���+2
�X7�s��Gc�ws�x(������h�󃌳y3T	R�C �V[B`vOZk��w3)���ڴ5$J�h0��K1╿B�X��Ft#n�d"y�j2�8d�*�cN�Au��s��E饃��dˎ�/�s@h�� N#�I���Z�+'A?���
G�<_��}z����k�4����> B�22x��
*�v�ʙ׏�N��݊��s�{Pnk�ͼ�|PD��
��~pŮ���Ǣ��EL�Gsҕ�i+��ҹ����`���:��v��\��D�K�-���眬}M4��1�'�#�K�ꣃ��~�����m;>~&cu��a,;x�H��+��@.	l<j0*Ƙ+��&w���)Y���K�&���=���O
����R1���5R��|	��:�=,"��;�[����iՌ\�fOp���;�c��=�����A-�^�A|��cTUɁ�Z�?/S�m/�9Ɏ��!{��TJ���;��M5�d�<�B>y1ҟ�A�	�����@�¸ɼ�i>+/�J�U��Y�����1q@`�Sq�
�?���((�,�S˩-P*��b%�.>�۹'�O��X���Mb��<B���4�I��l�P�ACuAkyF�{|�MR���?�ĩj+�h�ډ��W9vS�m�+p$����o~c��I��|o�����wmD.9�o�e�aH�y_o��~��-�5�0q�C$�`�3+�R�"U�Y�5ue[
���v�������q�����p�f\|�e8t�%8�m�2fȒI�Z2 ��/+�x<�F�}
9#+��%�_ r`�9Fd���o,������8g�g�O����\���x���R�V���������U�SX~���ŨS������-�����l��� ��D��G��t���"QX]��W���i>�ll�-ϲ�/�Ξ�N�@��̼��R�P �mJ���� [���)Z�p<�8���<��K�m�m�L��@��=I��Gw�P���B����P�b���j1`��}L���&k��H�����.����H��9+�/�u�>$xz���qpS�}(��h��G���j(D}*�D�%�v	}���R�b��/��r�v��{�`�}���]���;.�Jp]L��*6d��.�l��%��ɲ��m[�&��~�((�&�7{b��ߗ2��	�Ѯ��#^�n� l�9���^A��N���8Ty��=b�3i�Yu�<}ݖ�g�T��r���BYZ��P]���cc��4�����W$Z�)�v� �)�H'��" ���3	IX�YhT�v��%\ąsK�%���=|�@aA�ر�o�i]��ח_�f�P�{�����7��SBx����dQ�0�Kɵ^���� }vQ��˙ ���gHK_n_�^�UF������k��n���D�%ͽ�(��
a�"%��P��N��s�Q2;�O����A���[�A3�(�K��x[���w'���_5d(��Rh�!�L�Q֮�Jo-��X�#e�"�������(�h=΢���9�������E�ԝ�Z�<t���3=���G���Q�H��ܑ�79�p��W�NCD��
S�e��>��E9M)���?����y6/e�'�-���͖׋2.�I�qB��
Z֙u��|�|���=�J��;(_��l���J�[gΖ0~!E������w�z��B�@��ej����icN� 䊱�M��8Y���Ü����is�xi<M����+	-�V���3ȳ��0��|�� Q]��1�Q7{e{�_�����~Ղ��9�aV�ۂ�n�5�A����,�N��F;Je��(�j�	3�G�-�0�S�U�M	ms�������$Q&�E���N���B
��5��"�A@pɏo��C�W��6u�f��Rh�ZW�o^�8.�i �
����5X4 V%@rA6��/��E!W�W�_�n��1-̽��לCaH޾��D�%�y���
9�[�8���'��v@�y.R�94��]%�$e�1$�|u[c�܅/��k���S��\ɼ�e��ډڿ��u8�Zc� D2��"&��;@� �eq��b�<Fd����'\�6��zv��L���٤�oդ'u�H`�'��U7��}X�t��俯5,}�\Z�׈�*�ZA��~<�`I6�Y.U^�����,�Ι�K,uA�*N�(�����^��>,di-'J,�1`�8y�r�-X�s���. a���w��&��OvPaӦH�d�Y�(m�W>�Ł�kUR
vIV�A��ǿ�j�(����Zm<z��s�*B����.�u^�^H�����0��f�GnT!�?�����5������d,�{�� }�XS�(���d�u�-�hA�,���*�C$r���0�jL�x��b��O�{�R�<��2�?f��wu�ਜ਼���e9���)��l�e> |i�03K2l�$�m�F(HW�[��A��g[(
;!�LP?w�H���Y�^!H�&*+�"F�C����`It=��H��B`"}R�mW����ğ�+�1��˭\I���#�0"�ѥtA�^!w���j֮�Ɇ�Pv������hh|�����l��"�u51�.AB(H��g=��&Z��l��P��HH�O��4���7Z�����Nq�:M��#��݈���FIkҵ��Hk� �"����/�V1q�"���7����W�m�G��a���(�YDo�5������[��'R��4U��g�u��fx@zsf������.�(��R#jǣN�8cЁub�Ib�����c\�&W?|����$�ِ�L�tVF>�K�u�>,k5J;2oBi/�ݵ![J�6��8[���VP��}���!Z��D�-T	A�k�$��KMo���or��Ü!�]y�h�%�e�a��~�2}�4f�������嫙5rj����}�bM*�C�#.��^�]�a�b��
Կ�J��@W:ܗ�)Ų���|)�B�I��瓹u�
AQK�ru�-v�%o�~馪p�,�5P���8	P�$��^"�B�ag�q;��6<��fӳFs��/�� �� C��b�Q�Q�l���S�9��������Q@)P��VI��ϻ�#;1:BB��y�{����YGp�%�?�i�Y���� �������MUȦO!�&�M9te*о���,�kG��љEA���V=/��~��s��8�@�\ݥВ�z��+�Xk�g��bo,�<P����Zi���s��$�a�d�,d��t�)�@0�(5}ݻw&���(S]�$�d|i��@���Bi+	�Go���s��7� ���+��`n �4��fly��k>:�Ì�%{��D���)-^�aݩ�/awӏ���D�7O�Z����p������	F��Yk�qQz�D�e1�J��n%�P��MDՋ���s���� ���^p1��ŗ������@�OD��E	��W�qt��c�=�F�6گ�h�]Z���+ꅹb�Y~ڭ�"�`��<�b�y	�b&	=�<�vg�`��I�%yY����|/D�9V�Z��s���(',g@ �/��GW����SL����� �pp�xI��V����zFS��j�_ŷe0���r���`Ɣ� b �����{�*�)�R��؇ MFS��f�����U{�����j��ЇS�����0c	w�'� �TV��eR�ؗ��r}��telŦZȠ��Ɏ���f)�����c�Ol��!���RѪJ"%Q[�M�~k�uD$!qY� q%~�*��wچ6��~Z����E�[J\��p�6' �_`�X�8\1u?��y.���v����W�y俽�S��J?�?n�A�D{Ai��"�`��z ��޳�J���h䤷� �Z*T�צH$o��)У�ڈ
��p�︽܇dL�|y~���Y+����+�e!T�g�9O�E'A��[�����˴�К�H�F���Nu�7mW���[U����w��$�Z}���Sp�}�Ab�X%G�v!�Ӽ�Ke ������U��Z�>��PC�S�)%@ϐ̡�mAO���Az�:�!��/���{�q�Ԯ�s�v��HI'�?�n3-�}�ށ���;W3-i/��@򪱲F�E��Z�����֊ؗ|�w �6��z�B�jrI�U/��Tn?Ƿ��Y8�d�%��E���	$�ÿ]�������ZY���js�>m�e]�'���Q�88�tn�J�,W4��h�AB��E}b����p�����N%VO^8-;c��2��G��V�u_����fbߡm���;&��A�}��]RG�SK�$kaE޼��,vX�M/�fh0M��`�5�l��oHg�
q_:�J���	���:����8X4�-���l��)��R�d�]t���Ǟ�(�W����xYhq� X���>�%f���S::���NC��=,�Z��� 4�r`�I8z4u�.vN9�Y����f��Θ�L�������>3��-�7���Y�X��Tw��褲��' V_��n4��D�����.��n��4�ⶀ<�Z�Ç��,���r.�U0��RՕ5�x5�17��۹^GWM]��=�S� ����� ۰�x@`^f�����M�/�5aJ�w>6�8*`�*~��+B�2c�/,*rii� /�ph�Aj��r99׽y�"ߓ��4���;n��G�J����_�jIbVC�b�Q8'��Hpr,�+�%Cw��`��ُN#��$ֹ|6�.D@�.�9����Jҧ����"�<4�������7�3�]�����V�F�&���SN2���XP�`������@�p���h��e�O.��
h
39f$���`��v$z�A^.��%�jc1���5�;-� �Z�\�1vI���!ϸ炬��1�RJ(�aY ����IX�5�A/�ф����=J�h%����K��1�A�|y�f'H��a��!��DK�*��z���b}R�W�t̔%��n��M+jI��Y��߈���L(5ATq��������(��ena�Ā_,�\;���Ct)|��6�ţ�[�b�酲�\.�b�M���g�9�r���S9U�`|b�p'���9❋H�`j�8�#�Q� ���.�3P�RX����LB��A�&Ur�-^.�mث�è�sO^��û�}��w8]je��B^:�OdB�r��,?|ߙ������3u~b��1}��[ �9\���r{��/[$T }�5�(  ��C���)=|i.|�]�����0�M�v,ӵ�ɄG�J�<�v�Y��0�e\B�O�8�z�oTU8�[nw��B�^h=�r�F@��u�������,��ŭ��L�x���Ǧ��a�L6�h�8��k,�dh���5yE�uC��!x8�F���V"/c�����׎8��o�Ӿf��g�f��w?cϮϥ�� < ~���۫��M��gp9�]�^|f�e&f2�>O��*ߚYN���o֮�Αo5���fN�l� �\忸��[�[M��%i\ɶ���_���n�߭t��g@�������%��>\q�����/� �#Q:ަo�ȁ]� �dI�ܮ>���)�F�+�O~�6ǏP<l-8c�qr�r��.��,S�V��=�WX��(� ݿ�=�E#`&���0SY����=�<1U�wb?��o�ZO���>��4\����˾$�q�w�az1N���T�@W�,ehԿAJ��X0qn��o�~<Vr����^"[��%��i��bfy'�Ƴ���ⷐ�r
OD��Ҧ��jvJDH^�M� / �]�e]�Lڥ�g����Hw���<A!a�lw����k��е��ѧJ.Jc۰�"��|�%���nTdց���?�7��i����#�_��jp	'��]�Z"�m�������{�";�[��d�j9��xa��p@!��)j׃)���)q�@Y��Z�W��pk��M~�X��+�?��J����eD�zˇ��ZB���5��U�=��G��������Q'��񢃇�z,A#�5��#'��������XaU�a2����9�N]�Mo���*���E3짇�� ;�u�����}���3ϞQn�RHO��z'�j�ݵO���c��!�c��a+�w��w.��.�$.R�1�Y�B�@�w��{h9����AgY�䠘{�.Qu��1v����L��W>�Z�ƨD��;֞�鑑YB��"�J�"�s�o`,���3sQ-��_m�^<S
S��#V��6�s�t�*���_��DA��j�i�Ѫ�����uG�K�u��Ը�R�=T��L�����ڠ���=�'�_�컺��y���s؟+����R:�Q8�:�q�D�g}E�a��$[^gI S�3=M��{�9��j,;����?R��cCK�A���vl�r�~A;l�W���3��`rxƺ.	3l�q�D�H��Pz�t��eR�ʵ��I	1���d�}��	��r��ݟ ���O[��*��Z�jnH�l�f'�.�+�9	��_K=�ͩ]@����/������{�Tb�/���@�������P�	����V�R��E��h+�l���Y݉𙁚�a���?J�7��1=n+���n�CNwl��A,Q>֬B8W��Ir���Bd�:��0����@2���}`�$���W��OB.����Ԯ�E Y��/Z:eJGS���ZzrB���"�� �C�U	��"��)�#���h������y ga�wm
U���δ�WbH���T���N���8$�O�ci1�iEw�۬O��,�����ʑrCY�|�vCv Uk��2�'Ǻd�=_Dh�_�VL�u�_	R�����3ax���?����3k�	b�R�@$ ����?S���ǶSPĚ"o��aV��:���W��̼�a�w� ���-����������t��� ?�`�R�,Y��[�\�!h
ױ��l:�\�V����c?���H�2kf��J���=-N���>Ǩ�?��]���dR@��i�e�B_abD�MM��D4�;O���2,�U�rjD��N���y*(����[썽�sW�[D�0��
���/9�����g��&<��9��R�m��R�|՗�Č��^���{ɷp_3�/x�����9��e�_�^�k:�k�\�	mQA@��)�����~�G�- �H�=��sF4_�{�߮��c�#@��x����~�x_�hP"�z��+c����^d��%ֳ�ol��A���A8G�����I�%���!I	A��e��4����`٠��K�U 2��>����_n�*���x�!����$�#���S���n�NVʘ�Z�ϧ_�W�͕��%n V�hK��q��DT�/�Af��	`i��� XV�-����n���.�l�������^�V�n���\����B�VJ��6D�gB�%:SH{fHD_乥�^���8�2O�%[B�/�3�B^���~��xC�HgO�x�y�N��h��'�ȌsÝ,�6x�Q7(�'CXH�A��ִ>��ό(F��%��'D0����˴�r]��#��~9�+��s-���D�����(蛼�@(��*PW�65R���>	�4���Um�ah�PP�HHk���'w�a����S^܋��ҟN�d�Ny��r���w��A 1�4�Lߡ���D��^ܓ�������yP4����tg�)T?9�5�l�;�2�(���9T��i!��L���N��2�����9��<5VQ^>���e_��S\��*m���)���&�B� ���|�"%$Z� {�wbd�v��~]@3�x����K$�j<�z-��$����#*��1p��S� ��98}!�x�&a��x��1!^��&dvcx�}��]!,-y�����'VjJ ^�ʓ�q�px��L�%.�K�>��=��������J�jb��DW +�U�e���H�z*SnB���u|�َ�+v�U����#s8�N8fn���cQ-�,@�z���)|M��kUJ�7�@���K�h�hrBO�2�o�=3�<n�Й�ܞ�F+����'pr��xg����W�i���U��G/R4��T0{�3k�U����� ���'9e�P2۷^l[9��x�+��F�?��E�����ɍ#�����R���Z�n�����~Z�x��t♿�#�L�E�cr�^�荰zi��T,��J��_3�j�X�]�w�����1�2���Z�xǒ��������fuN��������R���H �U�ܤ������x�y&4*������4�cvlfq����i|�}=�9�"��X���$�,����?�]��Xw�}��0& �U�$���ʇ�:���t�@��#��Z�*��1���l +\�CڞĞ���Í�,��%�fW��kޞ	+>��W�T뚖)�a�T�s�A��@���x��;4{\��Q��(S�w��I�*�#wg���}�q��d`�#�
-�jz��
�Ч����H�����TB����^�����En;��̘��'y��;�^H���bv5&�ZD�~ӂ�����N\��Ă�ObY��LK����Fe3ܕ��c�[�#��ECj���"L�zD@�'2l���	 �J���c�L�sD���=�z2��R�kyg5ÌC�+a�~wʄw��%?Y}AD�u��[�|jm�)9
�1_D�:ߦ�+��8d�*xR�m��\�z�ݡe9VO������G�����4�>�9����W*w? {�0rk��D�F@N*q�N9���`�寚�ʼ	��#D%���Wh�̼M�7�#�<fqO��g�-�
*������57����]����'IU�t-��4��:�̌�в�@k �M sSA��Yo�A�y�WDހo�|�뫞���(4Z��dx�ĺ�])FR��M���4���2-:|����(*�b���e	]���nBw�����r2��7d��L�4҃����(��ف�[�|w6�Wbns��2��i g@��a��s����~��3�M{�
�<�h/��n�RC�� #̓m�"��-`W�`t��;1U$V35�F7m�^��5����^>�)fG��qa}����ٚ��A8�&>���1��{h�D��&��?���s�y�����&�4D@������&���̬n�� ���9�,�G�@���iP�%V]���5���Co���c-dH՛��M�]p�ee����O+}��cmw����	�$�w�|z�3-�b��F��V���cx���[�v�e�G��,π
r����Ne�8�vU�>��Q4���ӭ��`g>�B���H^��!#M0fS+�g�7+}yy�\��q���u�43�^��C�c͐���D<E���3�jb�X�7iY� ]��u44׮��>�&���N ����~Y>���W�d֢2	XD.Q�x�_���=O���P���>� e�f�T5S?�w�G03Z��6\A759+�}���K�>����v  �/{ܲ>�Q�ㆎM�]�~�l��([7< t�#�<p�2k�zx�e���"�g�����YYDjkƪ�^�@��k����K����7b'��5�y�2��/5>M#,�`F��C�ʕ��c���ه 3F	����"Zgm����z���S�*S[���h9*L�K�r��VJ[:�x��/�ׅ���{��S�U�l�T����L��R���P͹��rd�C�y�v��>��{��8V�e@�3�s#y�ft���*�zN-���N�c�Vn�	� ���)����_��z^H" ��C� �T���3����<��5f���H_*֊���9�Ap�V;(���l��ǳ"
����+-���_����Yy�,��ꭃ�V�>���aQ���i3����c	tf+�%˸��A_��	{b6�P7QU�[tg�`�+$_��Uu����?��-{Ćw$�Ⳃ�Z�
��j嗯G�>�F��n��̥��=���O6 �bC��GjӰp=Pl��x�xp-Ȱ��qJt'������
����Ю�v<�A�Լ�M�m"�N.�]�	��:|���&��+D�)[xl,�_|Pg�~��������R@7n�\wX��� �Z�X�
C�9���?傰�ϑ���*��H;�G��R}�pZ}���/�s���Hڠ5���B7�H?��M*:T����	��8q$jzǌ� ����֡�߁�[J����{�GC��PM��\����뛙�'4a��&D0���Q%�Ԯ��b�{��>�%�^�B0��j�,y	�wb?D�X�>@�R��}���4��(F�)uc�����0~�j���
y4(��d}x�,V��w�-�P��%e7��t+�����|^���]؛H�<��B �xmj��z���)��?9ґ�il)��v�|}�Ʃ`.c���#�2�1��E�~��7�d�g �T�G� �sB_H�~�U�.��k��t��-�-��<[>����s�R��dX�M� ׆hRg>&�������"C���e��⊘�|����m�Ȳ�xk��xf*,�QT���N?Ɂto� �A����y��f��Jc52���TJ�cO�1�r�*9����gLm�3�#��c8Z+�c�.�΀�GR!6��y:宺�9�<���R#�rM�bqգ���M�ʉ�ӡ��h�� 0�6�@��B��)�`�uR�[��" <����:�����1#Mh.i�|m�8�4C���������k)h5(w0Jt�g���&����0l�d$�5�r*:�O�G�$zsO�����&��+����eBc�J���v	=�ˢ���٨r�1B;!�����/�w:��	�qJ�$I�IJ=�f��X�W}����^h��^j�F�&_�A��Y[Hz���49s؅l�]�� .o�#<��n�|g���D�/H�F�H�U�C�̀m9#(��P���o�}����dyM�|~��_��~�ۆ�:-�����w�[X%)|ic�!0A�
�A�k(:�G��Ww��TH'~�n��P��.n&�^[$9=V��(���@vJV�v��w��d;Y����/��2�(W�����x<�ŷ�ٵrb��*�3��e#_��{1*�ꈭ���|t۾�
�$��E�;Pנ&��.r���aDe�h�[�nM�DO� f~�k�����y�|�֘�̂<1����r�Q!��֞�4mS:@?��0V9����o�-��]侵���t�&����n�K�](I������,�����m�o�wZ53��� 3��32�>0�d�z.��u-�V�G%F�P+�h��9��h�����+�[6f������!��p�:�x��y�s����>�JO5�a�Y�srƉ�/j`������%/m&^��	R����(��f�����	�Q-SZ��gT:p\c���(z��Bآ���\ ���3�#16w��Δ���+
��'��r6q��Ĭ� ��� +)IY#���Q�/	%Y���	8z߶)���Q��:�w}˸�%�nA�Ip�����y9�;*L��x��0�}�t?����l�L/��k���j�Ŏ5�oQ�=�#)�O݋]Oր��i�p��8�����ƫ>��:K�7�v	:��n?Վ����k�=ڝ�j��]��P� s6�G��r��{p]�`�\$�k��7���-o�S���Ĭ_�dd{�$	��El�݇�OT��%�,Қ�c�5F��J�ޖ*���~{Sf�5�W�Lw���w��:���dݚ�I�6E�Fp�����*���R�ͻ��n�Y�Յ�GŽ�a��v!��;�C ����/A������Q�i�� �v�+�c�g��c�N�-K,<��Y\c�Á�� ��B�b�P���̺�wgd��Ķ���iP��Ⱦ��|���Tpo>���:��	�rp�d�EU�*�đ��O�BA,�y���B�E�R
rz5��&�8;Y��6_:�L��cE�=-�QC���JI�7><���R.�Hu2^FK����jy/t����s�l[�sA[P��X.~<.��g��W�ˁU��s�f�7�7���x�����
�}k\�6��ˆ��tAz�">��bv�{�d�11���	n5�ڼ�xJ��H�����ɰ8�Iv�L��"�ϱ��@�z����F�kit\�=�D����Dv�'Ojz$�Bgrq J�����=l�?�Ln%	~���4��KN�=Uߵ�X�,W�Q��?��x��+��_q�&T��~k�dT�
2ιVF��v}k�����}C�^>�/�ǘ���� �ͳ~�Rsǩi���(~f�]I#閼�(�؉;S,���6�{����0���ouz������Q"�6�"�ش�҆��x�Ӵ�_��%���j�VN�f��"ĉ|�Kp�oFo:O�ks��$0��0��7+x��o�F�?x�6�7�-��!���0�&�Yػ�o+��ۥ>S�����-�? ���F,X-���w�a���h�ӄ�F���U4W���8�ω�?코�AA�\|�R��mN��[�7'h���PGP*U�i�v�t��1M�n��c� �7�U��Hd
S���o��U������R�j!������EmU|e��� �~S����#�N����@y'��ۤ�8	GEδ�啶L�ѣ?��`���B�����Z)'!���e
�5�_޵�;
�+���h��˖��3���S	��h!��t�۴;�V��-f18��G�����p�5j9:ie�J�LniC'��}���Q[~���[��b@��R�46�� �M�J}���h��Ҋa���^M%L��d3��sT�7r����h�*��z=�Y9)�ڍ�"��7�P�LoX@ޱ;�r��(c\��gj0a�+�F�-�'������s�j��ap�o9]�t�g9S�gm:�����ed���hN���q[����[��*�Õ�j��E�
Y�8lrpz�{��/6%"�=G�����S��	nG��]��٥�����ĸ��`��a�TV�??y���r�r$z�Ǣ�i�OKQL�e�p�w�N")�/i���~}�d�੮QkaP<{�[k+�-A��<P�&V��f%&�7�KcalTr��A���HQ�X����q���e�(�P��h�?0m����r�5F�yY: ~`� H r��Sw���X��iO�f�T����%5���M���9�ߕ���g؅��@ں���%�����ac�T��aW5�Ҭ����z��͚Ȅ��K�1��m�6��q�(���Z�9�)bd\�]T�H$=0���P1I��-~``b>։
�ͲD����8�J�ӓh�Y�葶7��ߍ��+�2�󠧮���b/,v�si�Bs�G�Y!�h���"(���Q�8Q��\����Ei�����t���_� `�~'(��Q��y��@�ր>w�� ��N�-���l<�����98�[�HpQ�xf���.��.���f���a!w��l�o3*=R4ʭS~�u���4Ch�
3�����=Y�������O*�)r)4\\A�	��[XձV�U��YV�e�O��PӒ��S��<�R��;�Uu�k�i���O��l�����YN{���F�st�����|��Kj!ھ���9�ym��Q�|'fF�!�w��`\���R��z����2��t�-���^��,��t���W{�K��_��4�H'��u��uՊ)^�\�.���l4�1��+;��h�a������D��+��	�߂�g���L���`H��=��zo�g˻�۶Ҫ�S�Ժ EV�ك���BJ�s,���W-�6T�J��6����;�lUZ��HY���u��Ԗ�Eay��8^uW��/�*�~1�hY�9�`2�o��ZWԱ����˸�, -��#N\����)b[� t��!���1�F:D�c�v�k���KD '	��!z���������zg���P8 ��3�n+;x�$���nP-�{�} E1�� �bg�x��=D��W0%�R���{�߸�.Q�.~-YFެ���k�������O���rҞ��I�?�G��r��:�,O�e.8�677�^�T�����2ʂf�yV�bh��I�R�Ug--�3R��3��4��r���4Y�vɂ���'z/I%��������>���f<�#���$7�z��q�O��1?�.�0�wfz!��l�7�I�	���D�4jt�����4��X+���o]�JU�@�tw�����g؇v�7��Bw/&Β�)�c����M��<�W�*O��-KZ���6��e�GX������(�FtEJ�g12@>#�����+�d��$�#�܋�I8�;�hR��,�o��)Y��b#@H3�K9�Ǽ��oi�w!)��~>����Ѿװc���ב2�؃���Ȅ��n�}- ����?[�j���Nj��\K��@:����?��F���������nx�|���CTb��<H[�Xp<��r��4����K�͞I��r�� �&*��Y{�%:��8�U��(%�%K�W[�ߐ_��ҩP�l��H�w�_Q �'���ی��2�A�k�z8=����U"���5���m�"�O��.84�Q�$xo���9�Pm�V�!=O�lq ��6�@��gܭC=��)/.��R���Ȟ9<t����+�o#�Z�L p��a�n�R�(tZ���$��൶�S��S�����M柽�jN⨂��%��@�(�m��r<�x�������s�<�������
64��3�r�����]^]�(P�z�y����z7�^�0�� ̞϶88�<�����kvy�� 4��X�H�|Ia�6��xSF�L�G��o�R��b�譖��٥��(�\hŌp�M.���<��fc��U�yy:���;B�b�6r���C�AUT�;�K!���	�2#�	[��5��D~��6�jw7�U��-Q�Z�e�]O�����[xA"{W�P=7nO��z���X�*L���b��ׅp�b��_+�=n��a{`��U��@���RqF�/��s�`�ѧ4;��=]�_^��y2Y�K����0��#�˛���X���e//�~ق��诊���_�kGJ���ġ��P���Z�>��~�O�XΥJ/%eq���kx5���.p��@��o2F�UP���/��Pq�L��Ra��f��<��\�Zfٕ����2V��� �v����ܤHH�i���$�aΧ�y��f2��H�̟qN�d��Q O��"6R6$�
�c���fp?d똫��^��v�"I�j��K���A���`�dy>�M� 6\u�=M[�A��H��k�J�^��N���ΈG�Ʊk^�M�#�dF� W��Gx��5ب����]��z���u_Йy[^��MO���8h�QLt�dL�|�|�ʲ��W}v���8d�ծ��	g5�L�K���r�Kh��/fڬ��g�gy8�[�,0ՍWV������3k`��!AO򩒄U�\<l�ߓ\g�n�`gt�Y��)�6ɞ^[��R	i(v ����[	�{�yx���	w��E��Y�Ća�{��*ޯd��Fw]��g��� ���7X2�NH^��Lev�-o��+�{'��d5J趭 �W���5fߩ�;�c Q���D�LfV�=�K� ���Ӕ6"z�
�	����D�V�íaf��dh��L��[\���A��[[�oLJu��_U��F-&i؁|G�G?Oq7T�B���56��? ܇��w��o����� *��x��֛_��Z����%=���9�J}y/��oNT{����*�J��Ն��iŪ/1�h��tf����e)T{��\�T҇53��Xb�w �v�>���ca�$�T�*�����2 �����8����?������Lt�hh��
B���7�f�^t�V�� ��U����X.\�C@Sw.�e��ۢ���A: F��C��tK��h;ו"��[O����3Пm���A��S\��:�����M���X�Gj>K��  a���uJQ+�Wٔ�?k]@��`�����òk�N?a��t�9l$5
��*,w�;`
;����{��x�%�Q_~[o�j��hC���'w�����*D�VH�K�C,XC�q>��s�g�U����}$~�^�α܄��ۏvY0�d���ws���T��֋�Z2VmvZ�`����1��J&K�nk���]](M���Z=�gXaܶ��󇳬���Јγ�p������);��]Wc$-9���5�D�
xsD���bzi����J?��-�_B}㣟��2�MY��ZѱR��:�� �1�}=�c;ɂ���L�lǶ*p��WGSm��M)>��Vb���6O� ��mJ�>�E}.<→`��.F�&%}T]6��h��GS��>�%���z�6��NC�KWĿ�缤�L*�l�b�-��V�Ap6M�죿&Y�T.s�+��
���<��ֈ��c�)zOX�Ӄ��wьS�$B�crÃt��l�O�<#��������0n�xh���Wv�`�0��D�
�0�5zh1�B�/	����+�Nռ��֭�+��b0�,d�Ěy��b�g�N�.k��n�T��E˓��ղ�[_���Χw�^x�7��;cpw��f�h@��m�Kz.�L���=|�Ņ�&���#��P��֥&JUin�?%R%-h�a�"@�Y |v57�̫+"[�'�N�	V��,���#��m�	���Ziv��WLj �oL�'��ͳ�r�G�C�j���n���r�a3�=�xM��o�@����^�M'��9z��?9��7�;�RFXx��,�J��τK��к,+e�x�d����z^���KZ����_�A���{�R���n��ǯ��d��;�e�C�dǪ��p18/�x�x_�U5�p ��_��O�Q}*��_�`(v-2o.ݝ����V��ݢ�����t�jewu� �$)�)H|a�Ў�3�w]�Ŕ��L���!�^�QMd�9N��6�+��]������~�lZ�&2[����<ۛ~(��.Z|<�����]ͫ�x3ȍ`�k��V\�_v.�v��zY����,�D|��ê�P�B�y��ې(S~���o�����]2��fR��!�گ��H��Q;��(T�����Sw��4R�Q��Ӣ`�����
� X���A�����:\�~q1n�;ע<�R��$w��i~;�Bi'���z����v3/���c�����(G7)\Xs�6���-o���[(�-<Q�����7Xͧ�"R򿒠��n׸��ʫwY�ȅaB�gnK���� ��L�����,羽����������[`'OC`m�Sl&M�.M��	֞�|wnz`GRE�ڶ��|��B|H���_��Ή�Z'�NJUb���ک�S��~�4�&�9����I`���|=5�w4��>S��� Ĭ`C�`GR��`��;{f�Lz]����Pj!W]��.Ě�aŅ�U/`��G"��o�x�ƥ��tga�+�f�7r��yJ^�O�,������f�4cl��@K%y��$�?̸���0��LLϺ��E�(��q�{�=�N���_��zb;���iD��
Us��B|蚴�g�A�ڿ�Y��v�X�X�zl��"�Lm�7]a([=��7��V!샊H~	[���˧AKю��� ԗr�Bd�S�U�'	�˫�5G��B��2�����o�OT�y����0�;���c%�T~nX�h�1�؎�I��yV� :)oL��L�� '�"<���VF�,��Tuި�Ö:%�1W���m��@w����\h���I�3V�J�z/`�g}?�}R&ĉz�u	@Ͽ�P��y�\��ۆ�v\t~\�L,��\�8�A>)���Lg�y���h�Ff^�X�x-.y�E�ڶ����?���'�:s �:�.8^}IAB!�R|��G;�}K�JXs�#͚'�K�h.s3c6��<�z䌖ʿ��#|*@u�P�Ś6M�[RQZ˕�{c��*��S��[�J.R��<���*?&�:�Z] 2قZk Q�nvC-�"���9��m���'&��f�Hhy(ǟ�����{�t�L�,��T�/����b��׎ �#�`��P\��SP<@$$Ȩ"bc<9Ʊ�3Q��.�+W�(t(+鄂.�o��վ��[�Y��i4��R_�-�_�4�b8�d�uQ�;-�C^l�5��n�3Pu����^HQ�>�]���R$�Wt��3+���܅�H-�NMm����#T��R�(�)�5�W �9����Ui;Ђ�H�H��[  ����w	U:���bP�q��VXD��������-�?GT�n�1X�c2�1bE��(?7.AjDaF�ձ��)77�h�^��N!�F JS�}�^��*l����+����a�\1�E��iV��9,R�(� �I
j`��(׉���5�0�%�o�==�B��*RL�o���j�:����4�"�UY{6�d/i�h��5���m��όA���}�tR��Q.~�m�B�] {����~ȏ���Μb���9��,c� �����,�G7������=d�Ek�Pz���g+�8�0��:�d��yh]��,�^�"��U|4/���>ص4������k.� ������7���-ҁ�]n���0Jqu&�KH�9���nP�Z������#4a/N�uG�pz�a5(�-UݗǄ�(�\��8Ô�@c�v�%�c��+��)�heZF �����qK��bd�N���r�;�n����n�+ot�>eq�������^G	�Ӫ]6�n�#���^C5Vq�W�b>.)l�g''=I׶�u��!���"I���d�{3�D��*�F�"uJ�W}3����`:i�p]D�Q��(u�M�ܵ��t 潸!~	`��u�r"���O��e-�T-Xh ���Ҍ�9gE�}�ڕ^�񲶍M�kj�V��|Ķ��]a�R���FK����A{zi	�`l�l��j ��I;J��f����%�Rr�B�{[�4=����]{�����~>�u�: �I��>�_䐴3z����Dś�yk�mu��Nzp�v�¯G����WZ���'���׽�>���ڰ#i��v�Í�u����_������.�����bNL@�)��p�f�<lW{pG;�G,�Cͥ�ى����;/�,L�������>s��He�$��=�c�}�;a�r�S�~<YK�T�HVOe���.���}�)(��>T7�#�=�,���T>��yN?L	Ps)�rf�SRw��F|MU��,��hS?8�.��S0�e�*`wh��f�T=�};g��J�)�/7� �k�ӝm���Yqc���?3�/	∝͹����O�V�!�U[�3B��u#��c��4@�}�G�@A��)�W	q=g�4F�&�r�R�Nw�TS��,��ɑ}��V	5�؉��{͂ȩ��y���w(�,i5?����tK�S��`��9����WU26��6�OmE�wMv낃d�k�Y~�އ����M�`%�������<����1 ����*��j�pp8�*0ӇQ�:S.�C��9�����4J'�Z�q�/���5D�(������]�|�ա������l���t��:Gro �+v��v��� ��N�9�gPi==h@��e�P����*�$��{+nX
��4U��}y(����\C�H�D�"T�����Y�2;8��\uz��J��:&B�x"�¨���6b��v[qX�6�L�z+��phHP������D��[��_I
ߙ?+��LD ��@���.}p:�~#�\G�MU�_3�z�ȱW.51r��4�EH���u�T�T�����:��^��R�ŽUw���. �|��{�����A\��������8sQ�Y���h�b�䃞T����0*d��6WL�q�/�j}PiM�=����D0I����˵j)&�$\J�9cf�yE�%������,�8C��A��^�OMV���ɔ����P,��Kx�G;*���g�'`��q	7 ƴ�8A0�4X#�Ūl��@c������~2�]
�9�Ά%HzN��a�*P�s׬F&��t1������u�z�ӱ�TAf��T��u��xbK�~���(R�q��jZ�E.��p�O܃9�My�3D�YQ�*��f�������EIbZ�Of��@�5yD��.�!�A��Y����a�������5EA>b�w�F���ϳ���5�-3�V�}��z:�ޕ� Ԫ�ܭ��B������]_\��0o
�i>�ү�L.?1���+��`�2Y�=������"wF�!U ��瑖�ڰ�8� F���oU\��1�
���0q2Wev�Z|B9����<{�v��7jڄ��>�ޚy@����ZP�s�R��͞��o�����!8�~�I��6�����������T��~`������0�ܓG�VGϚ-a���S����W�R2�u^�
 i�=ڝ�L�y�5\��*��OMC���M[f�����5�9�!�A<�5�ˌn���2��уȥ�r(����D��ra*��K�f��Bq%4�N�N��89N���<���c�����<t�+q�ö�ڽ��,�"3!��W�����ggb��8/�Ͻ-����(��/^�o�Sx��4
~��/�gm���
�RU�Y;�ȥ�`ESea�v�Q�N0{���>-�{hݒ3�A��G���$��p�6u���6m%L���h
�K��ҙ��y','�BϏJ�Oش ,�ts��R�W�Cr�Z����2Zv��~E�o����om�L����ꪈ֘TF�����L�<�!i�-�j���cV��}�� ���/�$m#�|뻯0��i��ow���Kf���oR�l�O�+��7)���b�F�D�L
�T�z*�~��1�z��Gm��MU}����`����������2k₏������x=�#�Z�*���N��$*��ܶ�_��W��4�1���q��K�f\o&����x�ɘ���F�Y؍���F2�Ypݏ� ��Cʊ�&���5=@��G��&�}��3����Y���.���jq��9¾} ݙt�}��h��A��Nf�"f`�tDl����T�&]O?R~c��4��!�[5Ωr�;T���3��	����S���(���X\  VI��e��h�0}�N��&��X!��l3�R����3��&��_k[�v�湷$���эݰ
)�Y)�lG�l�1�&��H+1�~�B�*%����Ԡ�d?�"V �����5�)�IW�xp�A7ñ�0NQv��<��X����Cl��2-�v]��������+��ǌ6��N�V�4�z�d�U9�Es1���>|SFE
�
�W����t�r�*�@��<�[4���3^I�t�~������A�f$�����Mh$���=jB��_ei�"������A�ncF�Ѳ����@|Y]�֊�v��E���0:��B��a�d�2�y�����̹U��7�h;�� sa#d��U�G�D�s��&ჟɘ�����S�� � h��.K_�Ծ�`Q?��X(��*p�IX�[a�����X�&�ܑ�F<�i87��c�=�?	T�F9�x���"��SIl��m�rj U.4��Z�3ÐJ���#A	�/��\�
��[b5錻�֥_6�B];���~ԏb�a7���b;�IC��\�����&��lc��Z���x�rT��I4�L���D襝�����g[� �=�t�o��eS�c�MYU���m�p��	p´B�e�r��^d�˪��1�t{,6$O����I��(�=Q5$�o�TV-�Rb�I��Cf�cri�u��+T0}�ѣ(�-S$�Cɸ����^7�Y:Xx��!D��E�@ږ�^r��P�xdĽg�5��.�9ik���L�І	*ݠH+�&)�?%Ք�]m�9w	ⷾĴe�:=���w��Z�����t�n񫙟�
���Z��V:��2�W���j�R�^CK�ɫ} ���swH�j�Ao�W����C����)
�Gsps�p��-%��ӁuV��g�+�{Y�a��/�*퐚���At���%y��@2.5�I2L}��m�����|�nT���<C��@��iXV���Z4�	���4h���
�=M��?(C��8x�ǆ��	��!c�"'��D�����'� �0�nVQ�$����Af��4�n��Tsn�8[\p�|&���Uj�)wd1��/�:�)&�İ�#�	��ʧ��e�[��c=&hT���9����ʦ_"|a$��l�	�72}�`�f���?���&�5m�q�!ւ�=0�^Wz ��^�Vw��MT�^k.�JC?]�2�Ҍ��Rh'�����������
������QՏ��M�r�U�ǿmG��՜Y��@��=�`��܊��N6nv������?B��kM�e�,*.�X��Y�&yi�'���.���!�������.�O�Aɺ�.�n� ����̷[sz*�p,������ug&JV����B�Xz�-7�|�7%�*ҶN��v��ir(����k)c�SP�duo�$
�����qw�E�P���-:`޸#��HIgqE.��S�<���e��F���n!�T6�� E�#�
�ۂV_k�8�����J�48[���k�jn؀q�fϊ����q�s�w��h��(�V����2���x��~�q
"�4��~�X�Vy�j�ĩ��!�]�����S���"�Rk�V���1���L��ӅT)&�I�R�'����?˻��'RH�0$�+�.��1�Ó�����8�K��$����'+�#o�w!ǳ(;�v��\���kn&d(Z_����=H i��H� Te�_�LBc�v8d�)�=u��fɬ�ލ�,�P\^�Gt7�����H1Y?�~�э�R�/pֳ땳�p b��.��Y�i�V�:#������������+Έ���b��"�~.D�8x��.��F�^w�\/�w�#�)��#�N�#�iK��e=/	�i�+����3��vp:)������2�����2�L��9p�zM���s;!H󆷸�eq��j����N�Y�(ܯ�9/����R~=��c��)���σ8	ؚ�1?�F3�����zX��d9p�ǚ��p)�-�M	
j������]*����G�Q�wXk� �l�~����P���`2[C@�o���j��"'�om��i[AX�m�<vS|յ�/�����h���u���_0�D����O��d-@F��xb�L>&�
*� �K��5詨�\�-��Ssw�&�q)C�z�LV������r0�)g���
#�E��E4�Di�	RF(�xw"Uv�h�q�OD�����"�"��|��Xo·Ƽ܄���p��QYD٧.J�:^j!>�5�g�k!���x7�jz���T�e�~��V��Yݙ׽���g� �[���Z80����T���φW���f�TL����v��In��=-w���D��cu�wk��B�����C��K3M��Z(��s���OK��|^�-��ʁ���S����֕��NFG���w\cϋ=�����nɇv��eS�C�ח�n����!C�����qP;�a�t�Em���sh�^�eimNq�؄m)���y�܊��5é2�`Z�K�1F:;i�{��R9�i�ʨq!�*��������4zϼ�Yoc~3C�n��#�_�Bt>V��n�}��ۥ�8i8;WHtNg
ϔ���F$k�[<����6`~�� �q�n}�n�/�/C��!)����@�>+*���ҜJ�v�p�DY��LIn�Z)`�]���q�iG!9mu��3�RY@�h�(/$c��y7���y��9BZBm ��Hr�bo��|p���w�NC�Spz]�#絆:^�9�1(A����9��)|��p��hr�ʁ�0��#�K��WM4��B�?��@��n���fv%�Rxn�c�V��!��J++c���R�aj6��Y�Ϊ͍��������-���D��rב��4/������{s'�������(����<!I5�σH�"r��z
Jee��@Ƥ[co��$��\�i#+���G�h8���C��aqb\!峤���z	v�̛��9�ܰ�p+j���C�$��f8*�u2Ҳ��$��E��Ae��ř�ok�>�١{{*�a�e�iU�/%���I�~�Y�j7b�ϡ�Fc$vNOS�u�s#����H0H�p����(˷�<P��tU�O�xB���=&��p�n�7��\���t铹Ν������?_S�  �4�Yѵus��w��ܔ��UR.�>�~2Y4����Qsx���ڕ`�`I���2+�%�G�XX���j�6��Cz��)�����'8ǯ���1�W�t�hG��m7<���97C/��ӆ��)�I{$�6��L�4ď�T�kaħ3�ͭ�*#}b��%�}T��w\�v�ς.��Q�P0�36�֑H��}bO���ʃ���ix<ϋ���T�Cm�AtU�+��d��%�#7�h7	����e�̻%�tJ��z�nٳ����Qmڍ�tD�?�����+�,4G���m���9?��/l�5���K�x�U[���E���z`b����n�ڬ���%�zN|������h�~�W���r7;�NQ�~ K�����d �*ӑ�c�T��R��L��SB�K`&�=���k��I!km?��Jri�s�t_t��œ��4.�DZO�:6�kf�ݮ"]H#	��Y���W\�sU�/>^½��Fd�O�v�	� 3�ml#��vm��0���Ǐ�V���v�z�L���Sˊ��U�9i�.����zhɻv����c�T�H���%=[�.@���$Dd�����rv)~���!�.�`�0������i.7-?������ey��DT�e5�m�<FXQ�&�=��"D�~�6�_����	܏�A:5!�|<�� ����
�y������D�"GLD��C��Pmԝ7��wNůmf�e��L.�� Y�#�Fgu���u��<�2A���%��G�r0��G��� {��nz9�B�겵�ّ gѧ�_�#3Y	L~�j��O�䖚�����D����:�
�Qp�g��.�[S�m�u��U�xL��s�	���y���F゜3���Ȏ�KBd���t�u��M�)��РI>ek��?�� ����R���QZ6���@�E)�)�˚�
�႟Z�:����1L"�������_�zh���w<�Ȼ
Yt�j<=���zq�QדZ�|����s�CV�xX��-�$x!���~'�%�ד�gQ[wH2�٠ȏM�?@���}Ӹǒ�QW0����;��`"��fr?�D��a�@3b@c�ۆ�$�A��$#;�/D�#H��\�8�u�G�I�)񃗱���◌>���=z=�q�k9R�F]�
,Wvo�4`7�G���p�����2]n��x>x�����>4��� �#6e����7��FI�2���������dJ�;܆�Y-4|~
a��N�<���0�F���ƭs�V��y�a��zF�ټ�t��A��?4l�z~݃�L
o�?��iۣ�d��}���ѣ_��z���n?�>n�����xW(����\���<F�b��cW�ڿz&Y���ӹL���!x�)�+��0���]j?�H:���6������lU�1ӥ?~����������XL��2�k��Y�X�-ܢ��~�v`}8G���ƹu��(󩛘s뱬~Q���~� ��T�:���2YO��Pu����w�u`�{zH�>w����c�/��ȏ��b@fX��`���$��ڒ�t�Kwo�7GS$G��N����$/�����:K�n:�s~ղa��u��{��0��b� ��5�ȩ���wx@ǁ9�+j��Z�,�X9O[8���!�l���N�dF([���%զ��#�W�f�L(�Zg|h�Bq����d���K�!�ۦ��n�#�P:�p~,脈�]��	$7Xɞ/�Y�IL�R�/�V�w����wf���_�`��uv�)�*x�I_@�h�?Gޯu	��V���S��P؛Ӄ��+2�(ԀI���r���>l�hJ�m<Ǵ��#z�e9v�?y'�)j���4֐�[��xn?����s�� �}�E�d촚���N=�׼"n�cI���	S�5
Y�dv<]���x�_��͙��Yr�'�E�_#R���rO|�h ���J'�Ϩ\qQe ?^�]0�J����2{6\Ó�zRZ�y���t��_����3o��Jo��?ר�~���}�������0�ƃ��1���?Z���,<�'4�l�P����ӵj��Qc���ɏ8�B���I&g�Ӟf>݅����ZU�{)�@�����r�i�0��A�ͥwQ�(=����u:.��^:S\T{M��q��Lŋ��z���9������bI��̤�X@{#�8�����,����D��MK�͔�6����j�_�B�,eګ�*���k�&�	 \����~}!��_�;�#Q.��bx_XUl1��
����ٓ�)���5��Iqa�4G�f���E�W�+Ev�������rFp��d��6���ʮGq)�d�;�@�P�y
��t�Æ���Qg��|s>�=PC(���Nn��5[�1�1�S������LT6v{�.~m�θJd7�yk�4��ék8�.-�Vx�t�����Ի��}w�H�dș_��V\Q�㲢�D/1���6��I	uY�qb�,���ҶU
�޷GZ��
`^a�a�g3#����at���>&u�g]҇�"�}MR҆��2LI�+r���1�dT��\���j�vl���	�4�Gu�ѓvMԘO�~wз�3�VJb�]�'u�bG��m�p��}�C� ����A���t;��f�����$p&��1ю�`[�η�b�<�\X��@�d��x߂�J��	�p����?tvO'�e߬��?�<��[����J�)Q���$T2�#���NK�N=t��Z��&s�3G]Š�k���Ub>���t���ϭ-&�
�[n^n�3�d܍�T��b;Ͱ#�E%����YKB�0A��o3EK���Z�%!�<����? V`ۚ�k�@���¡_�Ȓ�VV�3��8!Gi���yUC����4�����r��o6���XV�H��H$��Z�bW?�<��>4���|��'b�Tian=���kK��Ng�Ztr9hL�[�k�p	�����,�)9a�8�FӪu�&N������$���5k"��Av\�c�\�*C
��������vǬ`����Y<A�2��g ����/�+iS�@�{��0��[�:6�k����hJ��  /����6j&�b�ITy��c0��%����)؞��&49݃�J),�`ص���Wʜ��S�W���m#l_ �~.�8���k3��׍�֦��=�I��d��X�ק�;)����r�L`��Hvĳ{�X5!r2H�arX���]PW�xW��;��)��3���t�����:ʕ7�����@��LX%��i�����-��d���5��>P�R�\�:�q7E;w�"j�Ĩ�th�W)6��
�Y�aEVT+�Qv��;ۻ��j�W[�;��p�
�T^K.S��W����rh��Ԯ�,�&���3����@��F�s}j��\��e�Q>*8I�i�_�Ƅb��|9Y��3*����Sl���/G��������6�4?FD�����{D�|�O�x@��D�2��(��<�l?�S�FB66�+cM�I',yo+�|
 8�7�&ǃ$��_L_�!�,���adV�
K*�=��)�E�^X��5e��p���f��zz�,mt$Ơ������I�c��&R�@�ƹ���I�)�蜅�"�]B`-�Vo�FQ
U*Al�5�^"�	�K�h�Z% b��Jh6��_�Q�K�U�(�*ae�C�&�W`�=��@y���-4��)P����s�A8|���Z�տ��
G���ݽ!��&�(������k���h%�˾8[ �|#L=�w	����{�,�AZ�HuV�||���I{���$E�s*�ԸeK=8��c�%z�<9t+�oz���iO^IO�����a��w�_ �'�d��_�q'��=*����5�c�N}d_�O�G��m-V�_�yD�yT�����Ϯ_�VL�/�\x�s�Y��5UΪ�8���~3r��h���魈�n����A��Qr�����:����X8`��i���� l���Ȕ4W��V,]�' �����P���@�ynZ�*4�����3/e�;*�6-8�Tv�x\o[�����ϸ�?�;�Qz��l_�^WR�E�w�%ݡb3���+���]��!�r8�����A�9,�jg=�3�*�ӥ�E��� W	K��V1o�]ZG�j�����FNK6Jy���#� ���D�b�>��%BXk��:!*N@���Q!�(]+THE����}�vl��Uf�gut��0Ɠ�Mn�[8��۰���k����|1�Vz�W�i|�ؑ�T�
��U��-�H!����o��	u l��5�x���!���۬�0sQm/�ܞ�u3iv*T �"P�B8N�Ei_��n
HYBn`�4y��i�w����o=���{����][.^jei�7��Fw��7W;f�UQ`�94�gB��9��
�����&0j��۶��_�6��>2'�B�C�˿��2��;u��t�H�vE7l�c��c���Q��@S��Y?�.O{��A�S����O�ѴQ�o̲�v����i���O���H�ә��D���^��N]�	ϡk�ܒ�헾�����?�g���ʦ��"V���r��9��@@�L����N�=���WX�ۺ~�0�.�2�?�e{m39��~�v�UT��Z62[ !�e��W�Z��4a���O�j���oЧ��s#��t&�{�m�Xxf� ��:�J���#p�d�'�{ �]����w|Μ�ك�]��Z7�h��(;��E��ݬ��o��z�$�q����&���m	3T��Ĝ����l�z
�*�� Y|��
+�j���[�4�l!Ig!���	w��l��FZG:�]#�k}t�@������=�� uu|�?d�gx: ��n��@fT'�ϫĨ��)���e�y�KRmrzi�B ����kzc�Md�.�&M�}.a)փxP��=q,4Bw�Q�呠�e���s���l���B��^�H�;�@�]
��H�hP٨M^��e�vP-bQ������ �$�)�"���&)�̾<?�Q������+��+h�Lե@�tn�*Gu���qs@ٴ�&2�~�b�%e
���,#g/8���7^7zݟ�ˑo�)���zޅ��T�+�~D�c{�b>��0_Sh13��C�7�O���W;m��Z���+�7��g��V!��l��O ���;Ç���gR#�L���d6��\=�^�k��K$�Z{[~�b]ԛ0��':	��$Z�.�5�ё}Lq:-;���k(۸�U:��������f��Q�b��� P����	�����ań��n�3MF�",�\!3N�!��W�np��nX��y�)�����~��e|�Q�1_�Ԗ!.��q���Ք+_Q4h,",�w*X\E����$}׺[�}90���#�l�T���G��cG�J��~�n^a���<Z�f��7=�ў'�j�����琽O�����岫�`�ʞ0��TZiɍ��
�����t�P�~�@�7�i�(;������0B�MF�p¡e�9�Sr&�Y����Ɗ��=`�g��}����N����*�(��!��ʇ��S�2�\���"0\.O�4��Vh�t7*��V u,.��ǘ��VV���JU�*�C��Y"�Z��o���>Z&P�� 4j�Y#÷�Z/')D�JӽOD{씸G���!�
�8�iԩ�
a"F��yg���/Ԝ����� ���-��l��h����R��*T�&R�f*����x
��.�}U�ש7}!!�7����*t��u�?}�=�~Ky�2 �o��~�m�m POv���f�tLq̇]j����|T-;;�_�o߶�R�sB�L�2O������U\׆֖f`�[�=��!D!"�:Z�$�aȐ���hH�f��s�����K�� �q�a���1�a��}@�D��P�=A��[F��ǲ�hQ��\�Ϣx5�����$����1fL��͟�\j��\|-�M��<��5�-����C)"dK ��S���]3Dc��o �y�V�;'���<�a��jyhm�H�߅�q��1�s�.N�i�z�9=�W�ٍ�ஐ�d�<lb�U?R�k+���nk�=P�E���\�B����4٤_m�'_�����39��N{��� ��5�Ŕr9�(Gu^V��B��^�4��x�Hԁs�,&?g�Ԓ,�<�&�F�\����<�HlS�� �ve,�*��:�s�_m�j(����ӻ\�&Dr��-с@b`�,_�����v쐸�|�k!X�u�9de.&�x� 3|	�P��"4_Wɥ�Yd�l7�iӨ{�]UZi9����~ܗ</Jli��r�[�xz�K
����mB�6�"�[�'9݇���n�a������q�=H�'=�:�ުvp�Y���c����'ƨ�^�(as����H�_���^�r����,�@q�2S�E�R4N�5B�)o���Ja�܋�|x���/����0�=a����ֿEE-H������t�����dR�����Q���lܨ�J�����v'��z]O*՞cR8�;x�˄��lF<�ں���]�o	D���N���m<�J�*��v�c�΂�&�\k(%=�QzҬ"�IF/ͯE�z)��	dc��WE���~;v����'���?,�!2e��w<H�4��$@R��c��3�������J�2��XQ���un�B�:iD��:����s�n�k�)��[��G��g���V����ڳp7��L�]� _J��N^lfV.t�Q�������ܜ+���38hM>�����O ^� O���qX[�,��Nh��-D,8����섒��)/q���A퓣���7��''5�J\�ר�i�e1�Ǳ��R��Bx�	��yX�!��Q�t9߫�U�����%W'�v'd��m�t݉θ�	^���X��>�p��"~���D)r��zL@��Ճ�>��˔t����&U������yJV��
��.s�7�"Eav��:�������-�4�r����_H��F�M[Έ���#�*��]жo�58�֍>&QDt���"=MA�ef�ޜ����3Ѧ.�S!;oB��/-�L��_$];΂Y
�ԑ�'^m�nˎnȎ�A��b�e�d�D�Ύj;@)kl�/"�@�,��p�����f>g(9�-W��q��B,���^�璯?Ȯ���jr�/u��O�V)(X;�Z6;[<8����L�J�z|8 ���C����3�^���2�s�r���J��qt��Gd�3�#�"�Y���=W<,�5���M;#l-0���������0.g	udU�:��׋W�ih^�1YM��8lH�����J,���-i�I^�+M��|%�V�9�Ƌ�"q�����[��G�C��<5� ��W�XX�R-c'aF�ڿ�*5]X���gڬ���W�{�ǺI�� ��`р�wd�����O�Q�._A�9fM-Zr�}���Y6e��v��Q�jx6	��9�0�?�$+�.F����oȹU<Hö0������"��,��xBil~�G�| ��*�I!����Q����.�~�EeqE��;AkGTeQM����gK����c�)J��I�ڛq��K���z��ڛ@<h>��Urk�;*�AK�?B�D=��nFRvd�+t��Xh&����ɍ ��)(Z�0�����2����SPS��:<�/����=k��1��n���#�^q��B@YK�5f��f�A�|3�+1T�т��kl<���l�Ͷ4����������Z_U�Q%5����לA+<8�����ݢ��ˤ� {��ݞOY������tA��@_8UaOp�N�Fר^�mIj�&0������"#=�V��Dޒ��R,�O�U~��3�����r��� ɕ1ᴚF�_����ꄹ;��n��7,x*�}<��&�46����ۜ�����>��y�Cg;�F^]0B��(�؍���9&�:Vع��h8[�īh+��N`�g�@�@���4��wp���BQ���g 	��bA��e�N�8�w�%UP|�D��~�B�kIP۾��A�Orh�W��L ��-:a��>��M%�Z��6Js��~�)�w)�����W��5ʕ��0~s��G�a�Tq��$�H$i����K��㎂��E9^��t]�ab:�F�KS�
�'1�]b'<G�Ò��r�'�M���x�n2�U=*�H���l�.�P��G僴�My�~E).��U�[L��{�bK�T��������Jܧ�Ҁ�@�3�����(�#p�dj��M���4�#9|6���f��	L�ԙ~�X��&�f�����X���~I���h@h�U��*��#�US�g'H=UV�0ӯ�&�Os���i�L��/$����J�n{�>��^�f�FKfE�a���]�"YO[-#��a�����R�کxϢ�����N�w����Κ���f0uC�'�Y�F��Tl�+�y�H$2+Kx�b�$�'e(��=�u{)D#E�0��_.}��M�e�h�ꙁ��qF����Sq!���~�v�e��y�5ԣ�S	���]%���U	b�4���K�<%e~g�B�Ax��Y��Ud�����)!�v�z.(���+/�(���z#vgE`�J"0��o�)���ZF�`J�\�s����b�RЃ�P�d�hO�\�4G�����N��Y��)m���ªOH-L���,�q����7����W�>���Y��p:��Fs����H�Νd����,^n��C��iKw��=o'Y��j����z�1G#�f���|8�p�p��ޢ*,��#���)����"�d�7v�~�G��ԫ���]�&�7��"#4n�߈9�Ur�����%�F��2/2n����-ګ"Y�~}fb��my���]P�<U�!11>C�C�آ��2��ci�I��_ބS����U��Ce�x�0Z"F�*@������elMe�0b�]�g}=�6z}?�]�߮�S���~J�^t�����}J�܀)�D�?8�]�vyz���9����:�Fo]?p�Q+z^]�O��LF�+��C7R�p<x��Hi�3�F�TC5���E��,�_��T���Sg<��H�GF���X�$iővM����L5��;��]�V�x�Ӂ9O��u��	7%S���k��f�[bPt㘈��jq�C�ݱhܣi���a��<2�X���l &}���{�5O�WNsl&�;`�zbAu2���ö�õ��L��ԕ�B�^�V����F��ܦ=e'C������ Wx�h�w��U��b�9K�v�"LI���Wn�@���8<;z�4U~<��T[d2i��;��bV�r�T��G��;b��\���r�����<����d�T�h�?��{�M �L���M�{��E,$�߈��;��_��69�F��s'�����Y���7�^	3��w�,���g�L��J��g�ViO�a��r���������� 0P���������]�K�
5�z̀8>I�Ig{��[����x��y�8+&�e������Cr��Yi~H�1������/O���~I��G��e���Q��-T���f#0a�;�K�,��f�*��?�3�������A_��[1���0�n�Pی)jg#؜pI��ٶ<�G'���~W7 '�D��򣪸;��ǦX�CF���<̚��Bv�B�К���D?4\���)@�x�����o���X;��(�������59ܢ������Nz���'�.���O�P}���;��I:�����o���9?�����j�y}�!1X�y0h�7b���B�7t�)�����
0�����9�wZ�<�����{�Ú���O�0��`���:'�OyCM�J5ʥ���F��/��P(��x���h�sEu�3Y�q�,��Z�E�eL��xx��ȶ��`�bV���Z��!?I�ς+n轉���t(����{̻^_�������\�h%�2I��;p���7��Z~�8��6���u%�S3�t�2˦E\{�VO��&'pR�dx8܎Ш�[��'�jwb��Hי�u�џ���p�A2�D9�gMn�>��Ȣ�ʾ�H׫H�K�^j��8A���,.��� �VJ�Gv:q���n�P?
��|!�?^�~�0�~���Z]0Û{t2�!�I��@��E#7X��V�u �E��)Xٲ�Ũ��±�y���7T+��I3�6��cU�36��P@E(���
Ot��"z��r`hk�6��h�(I�8��d��,������yG�*�"�]�	3D����&��l�5�s��y)�T�ڦ,�;��I)����/�� �{�l7��y?�5������j;|����<�}�r.��#н�I�L���	iTt��%����V�E�ƪ�U*�]$Ow�(�������d@!�U�)�gB��ˬ dm���ʥڭ����[MMK���0GPC |Sjk�孿	�����x<#sp��c��5�^�|��j����nz�j��9�2ɶ�Hغ�hbo'0jB)5_%kK�c��؝����D�Xk�v�׹d��O�ȷ�����ߨ��k�ؗ�խY��̄-�(��*0y�W�O�����r
���<����,
�t�֬c�p�n��4�"�Q���j�x]|�a�a���y?M�&�g�mѫћ�n8��E�%�����d[
���W���0uR�e�Sa�b�6��}�H�$������ 'Y��Ȳ�C������i.;_�ǊB�<c&L��^��&~�aSjT������P�wG"�0�ގ&🥜x+vƌV��p�re�����0|!	~C��]~ �ɕ\Z���)��!��^�oq�;A��iƟyb���iH����=�AU�45:br
ga���?�puX���}��3����ou�z�O��d��dm%�;L����ӯ0`�F$�P�����+�5�:1'�9�����#W�\���-�W�Wb_ |�!��tȗ�fQ�3��l*鍄�N��4�v�B��Z,U�{���.�P��,сk�PU�@�U�ʎZ�F�F~�Qۅ�x�/ '��T�f�� ��Z!(��I/�������\k0D��&{v�9Q����`x����=��U`uu�����u�[枰x���n���
�F�6�ʐ=}ۼ��H�!��w���˫�!���?�̆�t�f|C ������9�S��3=���k�Fj�.wgnf��R��T㱐�<���E&ÿ�)����k�7H�� 93%����\��}��,�3�q��o`J�_S������)��5�n��5o��;G��-�֊�O�M��Y���<si� ��)���<ޝ+�h�`�W�L��<�蒘j�2�֮'���k�.8�ۜ	�
�f�~�G��B�V�U����t�]��?ـ_�	��bk&I+���ݡ�MJ\
�_��g�R~�aFw��I��m�J�=7�!�dM���� ����t0aÙ9��{$yF��V�0�LY�`b��32�Rр��c�:!�A��:�|�б�J�.���_ܶgo�"\	�=79�l�x���)0B��dN��X��lf���5�H�F��ۤ(��ݟc����Ȏ�p�u/��˾l6V�J{����H�C[Խ"?L� �sR�g(�;Oz�$��7,Z=�=[�ٮ|	�}�ݷ��kC�������Zn[]:�eH��ʱ�!�ڌyS��D�i~��	;3�X�h��)�E�RJ�Uξ�6ǔ��j���Z���'����:]7��?{s��l~��F<��Qw�`Rӡx���\�Vjv��p�*��@��3�5����: ��'���M���]RI*Ƴ���~q��#P�]��TڿI�4�7�Ǝ-|{�+��&�*��@����~��
3�Oɖ���������� �	~ ��}9�GX�ch�u���P�#��G)%tPƩ|S�}`�~�N[���������,�-|pST���b�buX�s����J �����Z��]�1}�����&�DFGB�գ� ��1��$��]� �5Ft�"���̘���ש"I��t����"�޵#��f�Xfxm�mw��'@z�|�<1�c���(Q���(겤��!�eU�Q緤�=c��$O��Gm��Qǥ�ZO�� �	���MCf������bW�����j\�a�N[+�2%�R�@ݏ7�wAYSk���H0���.�I۸Ղ�Ze�ԧR0|7z�P�A��m���� ��}�!bi2�ϟt�LL�
k)�M�н�/%,�L�cPHL�okx��؇`uOB�ȵ:R|���6���Jp�����hh܁�����<?6l8o28G�R�;�G=��1o=� 10�6�d����t�`�߶7��Db���u7�mdR޲�}�`&����8%BG#���;}�<.X�{��b_)]�]��
�t��Ј	��y;O��B28�w�����5�ȍv&�<X��r�x�H�����s�΁fZ�+NM!����nM�fb�� <yq����4�R�±*	8�����ޛ�r�M4d�+��	4bK5�o��`+�K����7����G����Җ�ݮ���z��ƫ���D1�G�� gA�q(�1g��!��@��+��>�T>Շ�I��������*�mu n����|_�T%&#P��ե��ә��3����'�������l{�Dμ/䊗A�vj�<>7�}����_�{6�a�t�n�sF�OTE3R�o
h� �&��E%����W�e�.�>�#����~/�VO���|{ڢm�q�w�R���d��@h����;y�
+mT�U���G��y O�~cO��](�������m�F,p��z|����+qE�H�s�0��C������+f�>�/��ǩ�c�����q:��{=0��k���+X�@����/�C,�T�bg�����H�t~+�ȗ�ah~��mgvBv���k�;��!�䡻��ԡ�m��хf�����R�
h�Ʌl�����������`4�Bh7���/[J��E���W��%<]��Zx	�4h��9��}'�.M?m���Y�`����w�f3�A(��N&91=RD�mQ�)\vHݤA��*��N��t.�4'�/����SkO�G�v!
2�e`/<d��u�ԛ����"�Џ�7xyo���i���w����Bs�Z�D11�1��#xfVa�7.��n�-�7V3\=F"�>e���zt��F:7���g�^:�� ܏k���Qﳐuh��ۉ�	�I׎�v�} ;��f䖡�<�/3�E �\�G�d_�~��o�a>}P�0�آl���(xE�1h�ʣT�"�#��A	O�ǱT��U|��><�o��C�>K�{��c�$��
��� �n����	�� �[ɭH��5&.�8��9�#k�ɪ˳���F�M�#�⦈d�ݠ2�Y�����?J1w�k��Q�:087@�!'�U�'���oJ��B���	/fppyEtf�_(�sG�I��"dϞ/>t�BF������܏v�nbo9�u���Z&x�����;�<ɾD0%�7��i�]PY�4�9����LG� �[}@uSk�*��ܜvi?52�ҍލ���"��&5�E`�_�8{0��}�>@���U�d#0�k��~3���������jgu�'��ܹ\þ�TJx� tsT�מ�ל5ݺ\, ���-LPS@v��f�UYݎ�iCX8��g5m�q��
.]��j�L��]`��օax�L�)��H��  ���ϯ��Yb�0���h�/�)�t�k�*���>uj�{~���brߎ��a�&��B��Ռ\)�
��<�/��M�ح�И�~���r?�c��M����=+e��jd3�Z ��i���T��M��P�¦�d���� (k�"9�c��7.gSu��j�3�j/�I�����,ĉ*��%iU�	`6��������"��Μ{fn�Ss�ĂMK��9��W�$�eH3e �~P"��v��R�)nB���٢	�o�̀.�/��ya����:G����=�]��3����=~H!+`��!��,���!`���,7O�1Z�:�A��3�&\=:-���|�jHb����@�L%��$Y	5bq'��6����tňq8_]��z��6��[�fS}�w�C�ݛ�9l�������T�W�/`2��W���ã�s�h	��c��<��ә4<y�&�4���6X�s 	K���m00��-l}�u��9�Zx��'@���*��ߌ�<�w\"�����`:�u+9�nC±[�����b����W�x)OE��2F8FÑU�XC�ӨMM�>��.�ch$D̖tQ��77�����d�L����iP��6!~�4�SHу���RHHf�_�� e���/1���)z���aD���~Z�&��$�'WT�������&O��gb������W�D/�gы�V�ķ&���-_A�4�K�r����k$���0����q�8�b�3�4�=M"��cx����������'\ ��*B�g3�(��z��3�|�0{�3�#;���r�L��A�|��`2֍ry#��y��sc��<�؉3s�x՞�W�!_c�r�=�Y�_��n���A��)����G�^F�uۙ��j��q	}@�.Y���S���H���y�x��]��(��t���b$?��࡙�o�	��;�k������F���-ˁMh騞D���C�w�|�q�`xJ��-[,_�ڦ�ErY5#�Ͱ�B9��i?�'������;lڕ�Өu����t�<���	*�ˤ�^�6a���fk�K�ظ	:�\����A����?�d0	3d��-ʭ� �����՟R�bYr�wF��+I`���=�_u���H��?��(�-�)l���Vn�;^Ŭ�x�}+.{��i�ݐ=HGHr�5�&�Tr�)e�2�>��{r� 	�����o���R,*������"����O?��|]�3f*S�[��p�+��Y�1��)�pC��=�xy �ql��|�Ga���q�i��ϱ,������Ҟ�ҡ��N���b���+t��d���<_0a�cܳ*H,f�>��=�܅뮢C1b/��Xe8	�;t�����"�m��i�͊���)FP'l�+ƢLMlj#��X<a��>o$�����<m�`�T�.�5��IC�/3]�
N%�����@�i���%�V��S2�y{I�b[�ҥ����!DJ�	w+~5�&��M�Ё����iwy �ޜȬ��\�Ӗf�b׺�w<=�$�#�Nr���;���K/0ޝ6���Rй�1�n��/�{ِ�٨�S�p���H?+hfy��u�-��4�;^��c"��(K"[~��s����6��#O����`>����4
���]<���OYZ#[n+8Z�vǵ�-�%����U�7w� �$<J�0��iK��5�[�d�ZzrH��p������H��x�J۸��� ���up�r�`�:�����~��Z���ol5�čVB<uv����=܁�U�z��$�S���d_��H��NP����P<3B�fi��c�@K3��
��}x��b<N�����r���s?�F��6F�0�
:����楙C�������������l��V���`W�K�i�|,��,�8��x߫y�k�4lIv�@Z�%GpH��5|�4�i�NH��d�B��!���;��BG�?��,X�oӉxs��4k6N6�h=���Eu]��T@�T�Uck�jr�D����&̈1�cd����J�"V?&9��t��U�k�t�d��*�=l�{.���]z��ʽF��϶m|�V������G�;�ܳF^�I\66F�*�O6T jp�H�U>��c�C��l�4v0H��h����̛���(6=c����ih��rK�����5Q,	+�u�P� �ܗ�:A���j����;��Iu`K$��o�P���?�tZ�ק��1�Wt��E���*�Yh��[��`���2�x:n��E^����7�h�ܟ#Y��[?*6��K�� �p)�^z.��.żh��gH�~��$Ls=������{���i�E��E��kG�(�$֩�`�Ĳ�B1�6�_�˳�Ϡ�j͗EI˴�,���������� �|�+�TJ!g��̊����F��6�\1VW� ��]w]j��#D���L���gz����,�aQ���j2�(B�FM�4]�H����k!	D8[���E.S`gv8�:"������g�"��|�d⏭��ڪ!{�#�V��<��8�"T��<ւ�0g>�tm��=�� �wr��J�]Q���5U}��M,��k��[�4����Fʩ5��
��e�*o?�j�!Ҳ�9��/PG��y|��;~�E�r�-h��ӏ�H2�㠌�ۇ�2 �?I���)��h�Π�2�{@�\w���xTr�߿II�g}ZN��{��v���V�K��Qa�߭F�������i�٩�`�w��˒������'1����l<cH�d�v�7�EK��u��� /�j.���Ǝ%�j�nEU$}�#��:���k��8�D,��$7p�۾��b�F�~FŻ�,�8��W����Jѕ���^������EL��[2�b�(`�)�W����'�{Li)�r��!�ߐ��HHH=����$r�;f�zu�eT��ٺ�Q}M�x����cF�'N���M�t���v�Ѷ�BN?���ɰb����Y������yҰq����{�]S����1�!'�{�h��N�8;�C=/�=ƦI,+{OUg�3�\76=,~hU��c��>���Rn)p����������7�s ��&��.@G_���m$Q�[���"a�N^Sݢ��_�p :220���ЖcT�f1����5���`��neb�mt�y)E�[�-N,Z��������W"��Q���VQh�$8�@���_�≺h�I70	��"A(	pگz+R�^�Y��RÀN�Z��A#T�hy����Vs�+��*�[-�N3��!8�����U����Y���6���t����q�C}�ꍋ��_����	�5�Ѯ�0'��r���p��e҉K���(_�$GyϺ=N�JF��|*��RU�|e%��
�����N�WB��4�������z�2�����kg�?DH4���8��}}w�	��h�u<A�1�1kW�`�ClFز�,7Oy	d����Q��j���^�7�֠�e)��� �iV�С��&���w��3�W���yq���!?�L�D���J����Te�g�+�Eg$o3T�f���g��kO�g>ِbnE�m�(��N-������@��|z 9��B��(Լ�zO�b�D�v�K��ݮu��t<��8��E�Cs�F�B����Jbb	~�[�d�ܳ�����{��(�"=-d ���`�L�s���0���k
I�q"��}�'?@@F�#68eW�����=h<d1ѽq��#i)�܅N��Z���c?B�pi�� K�3�P������3q�i��#��YZ�o�0ȆF5of��Zy<�!��X+H0�q�_� H�Un�=�w�4�i���{�Ww��o�/}!?�e�O���IW����ԅ�6F��I��3�:��ᩍ��鵃�1�/��=ᖼn ����?�R�o�B�D]�7\F�������-g�������C�]|%0!9>�����O��=B����Q!�oh���~%3¡Dx��y�Qn�b���7�F�x�Z��迚�>'���Q�Y*���[�� Qe��C��:G���5l.��y��z.��7�Y�<A$�t1.~
��. ����ѱn��`&�9��_����e�[�?(6@��˪����1n�M�M���Q�"qcz��.��f�'�>Y,��(Y�9�'g��q����`8SN��S�^)?Q�py:�]J��)�nͤ��<�\�_\5�eQ�"�R��;��~��EC�_.�-��a�K�6F��xUyP�-�ٯ���s
�LZ����EFC�Y�$����C�����j����M	���6H�*O��H�e 67�J.����6V�z�eD��$��0�����
),p���t�����2�	���@�~�^f�D��v�o}�_~|�ݿ�w7p��x��~�kZɠ9�l��������btBt�4ռa��t���	ؼ4�i���:�w��þ^�����&�@؝:�Ƞ^ҧ\A5��'�Ɔ�dk,����=U!�a8����Ő��˷-
�3�ڦa4�43*��Z����X�.f��� �0���4�V�ޥO�pª��H�(���[AkZrF-�dL�k��H���iגzL����0��u�z%���D8��@�}��ħ���Bk�]�,c�L��l�(L4�/�\���� �'��uOT8�L��>D�7Z�C� *L�!t��[w.P�v�T�BU��ާ���6��6�E�f����Z���]��.�6�ܸ��G���IsLr��Y�ơ�Z���BI�_�P�s,�$њ�u�IS\�p�oѱ&W�����h+�=��&:o���_J_p����<���UǃJ˄�&��G�g���{�ə%œX�hE���dT>E�;Y��������� �՟ʔ�(�[}\nE�k��3:�`o����a��(�e��3w�G���=,$�Rƍ��x�b�t��4"�l�*�=L�e�ӕ������tY��cF��Gu��D��)���e�1�����.ܤe��<��x�<���\W� ��u
��4l�p"�@6�#Ww:���U7�0/^pj6���}l�����|t�?2FBN�>t;�0����Y?�Pi}}�1'H�x9}���=��;���+��Ќ�]�pIy#�����������Z�ՀNBA*%� ]��V�Q��J�jp��ނI�	������H�P�,�(��_���\�QZU����Hñ�c$�m4�ksjYc��v��t���n��]%�R���
��򿊷��}��:�Zf^8϶Nz���%��kZS�����iGa��Ֆ��}�ڢf���C�e�D��E|UȆ.��Rl8\.ޑx��xrqX"����rɱXn
jEa��IX��K��8�;�r�X�?��s��G����#�42.l�����+-L%����Er[{ֶ�Q:<�G�q=/����O��׳��3Y�D۟�,��m�?]�bk��K������fϦ�T�J(bࢡ6 �	�ڃ𐠆J�ٿ��Bq��k�{<�'E
'��G��o_>�Zn�P����K�M��EO�J�e�F �!�fL��=���ާNy��?ܘl�(ñ�\�\%��d)r�Gx���9+ݍe֊��2v�yG3��n�:����9��a���śJy���[���&@�����
�d�e�C8%z� 	J*�^@�����O��bf�օ~p��D9i����.)R7>5i!��s(���{��p�c�]C�@���?@����]�5�5D�VS�W ������N�㬅��a���~a
�.9�զ����~�|�?�7Mr/���'%�<8:bո��a��V{���� �B��W�Q@�LD�,#%8��y?�r��kqlwӄ�zs�xũ?���g��7:��n�ࣃ�5���1!;�d'������ԧ���1C�d��)���5c��,q/�Gs6�/�e�3����t8���C$��Y{4&>[�7[P�j���k9+��Us����s.:(���ֿ��߃F�
֖6�G*�;=�+'1�y�'�2��h��b�(��5�_��'5�#��j�@¶��Nm���й^!��P�M|u����;ǩ.�M}���Y��MoiS���y���|lA�����>�j^q��(��hq!&G��K=�v�g�u֟�$�費���%��W�i�Ͳ.l�(�l�����'sj�����!S�����qˎu��B���B��}m"�,�pChC���AE�`<X�_B<�kq���#1��Q��n����F?\x v��C�UD���?��l�5�L�G��Ӛޙ+�i{���|L�f�����X����+���϶YZ_Iq���1���WU�Ҕ���`O��N� �a�I�t+l�H���wx|�jSo�fP[2X���-�C��bh�	T
�Q�}�����ɍ	�R��N��3NC�eę����.f�f����y=�"�~M���<�gF8�1w��6Ĕ�j7@���Z?Qi�#_��cM���2{smto��q�����khu�d{�N��A�x6^{�����U�Po�^�k}R�I�86jQ���v�hb�H���eZ)��D�^���Zw��q��P?�\C�u�r�6~E�v�|�S��Nc��Qxn���|5�*�}�t;bDw�%XG��z6C��ޕÚ�/zo�K�v�g��g��%> c�K&]+�� OC��a���/�t�s�����;@���8��(��(@.R�x;���ݙ��&M^��C�W1
�&}��1�Z�04�^#�K��ܶz�;D�)��=�ݵ�M�8�]���(���oL�s�-���q���jK���|��+"~)eKB���h٥��ُ��XZ��"��K�}ӯF�|��%� �滵3m
D��B�T�Q��"�N�'�T��p�O��UKh��]��f��ĩB�}�;0�"<A�p���k�\���qj�wl�8�Iq��?
P��915X5�cHT՘a��]�=7p&	ā�QPHHT�����l��\/ʹ�	)����J�X�a�����p���Ҡ����~�������E��f@Bp�u��\��e*1���iӈ�7�ta1/�R�ר�^�w:�L���i"O��s@�z_��!����n�걇&�/^����L��l(*̗�$ఫ��Y���F��?-鸑A��|iƧ��=	�͝�T�( ���4?��Ax����\�&o�P��5R9]�j�t�
�ׯ�ڝ�	�� �(y�=o��C�ŀ�M�{�F�l���fn��=t��T�Qg��f�c�D�Z�v�Z�x$�����?"�'�( 
�@���6l��(^貽{��|�S����H��Ȅb5J�Q&�dwwz���v�z�5�>��5�0ߡ�G���G�Ⱦm���L�<*Y�G��z�\8r�d���qW�M�t�t9o��'e-=��}�h���;���.��?��. L}��@8v�v�S�ӝ���-=1��vҝ�I��2��5�7w�+U��W��!�����+�'F����,?Jn:1ʷ"P	����]GF̅�}|���/��˙8C�
�����=X�r���E������d�A+�]�+� 5z�ħ�7��1,l������M�;�݈1%�_ڊ����}��q�٩��[@&g��?^pj�[k�x������_���1�|"JR�Qn0]�]5{FB4W�@<�]=���;i���h�A�,�76w7���<SƩ�����}��t�'�%P�ig���<����<g���8>S?{�O)�FQR]�%m��A��&:��|,�Sߣ7|gKB��, g�%	:�U�jǾ�b����s��a�5k%Q�˓{�9IvcY����HJ�^I�u���q*N
�D/�V�Ah��^��qX� L�]�}�,,jG��t��
>y�R�09q1�}�b џ�7�EY_R�}��Qb�]�Q����[�B!8;�ؗ@����V��.��jJ�A����Rbs�F�T}V�1D�|E���@��F�����qʨSk#S*�)b������-���q�֪�0�눛�8�bD�쮹aM7lt\G����4�����㨾��ˏ,��/bJ��J(\;nJY��w?��í����q�fo�+,/�����&���QF4�E���v�V��Y%]�a�HNη5 �줲�]�|�X�+hT�0V U�U$7j��ȩc��m��a
�sNt=�Xm9gV�!S�y�Gz�5�mL�Yj͢��t��l�j�awԙOτPJ�,��1%i��+nAQ=��Q�D>_��L��}vLl.Q�Z��2Q�%���i�U�\�
��A`"c�g0e�vR"bMV`z˲�b�
'a�yN��U�{	�G��'���d��oܾ�J�Q��([0x�̚��}���l$9���u���C�:���uq)�/۱��g6aU�H����z>����4cO(��&h�h�صr���q���y'ni0��I��WE��0~�fΘbe�E�s�+>�����e1�Z�����)�7+����1RX��#��`�U�ح\:'6}'��vx�u
��P2J�I��<O�a���с4�!hN�ڀ�9����K"��uφ��4@�ߜ��$iqƍ���띨ȯ��t\#�p��2�fԶ֖t��L#�&�P˸�e�
~ЁEv�������c�����	�rf�c�i{������$�>�/+tr��mj��*�����  ��'N-&�o�n�)�[����v�e��Js���L,%j��s�4GԹ~����Wd݉��!o�cP|<6-�)�g֖Sm��D ����(��=�lh��U�F���~��=�����Gj�Ȥ���Ŷ�a����Sc�5�,S(o��zUr����%��i�߾�_�o3��I`�<��dK�0��mJG}��r��*&�|4�W���e�#����O�.5Ӣ�E���]nD�
�U��)Ã�}��9�j�E����u�����׶mn�ٙ�%� *�W�\�����_�-�i�(��������tYh{��Ԩ�V�`��k9
u�'���8�. ���#��Ť}B�4���i���'%�xp��~)G%E�.4�D�Lm�2#j �p�h��ڃ{�j>�'p�6/u���8��ć�+ߐ�u1�������i�Й�����`?RV����,-�ޖF�2G�v�Y�����Q����/�%s��%��q@�R�֘J���!9�d�yԝ��WXxL��91�Qԋ����L
�{����h�EF�`{ծ�����Gr��[a0MA��<�D����f��
�C�ҥI���#\\	����A�EH�9��9���`���� Ғ]w���l��6��*�J0)Lʢ%�6���t7�ǜ_�N���h��3YWb�y=�<m��l����
�f:�_�&Q|�RjY0<�����2 �����,���<j�E?k�k�V�j>�\�s�H-n'g(��_s��2	e�?����.>��;�����L$��`������ku�+t�HE�JN��@ƭv]�|�I����X!8���ehH��Ay֬�is�?�s"��4�ճ{��_�IԌ�h3���6��O0/S�T��4`��j`� ������4��ق����o����v�V؍)��펌�H!g��CL,.�}ލ->�f��d5�n�����Ic0-�r�$�ٹ��^�� "��H9۾�v�1�z�cqҒ�nR�3&��f��a�Z|�}p��%���
)�}&����%���@ܿ��$K�~��:~�gԖFp��|��+�c�8,r4��]P�B�ư�7Pid/u�|:a�E�\� ��k��X�!����U�%�� �w]�����owu����[���b���	�60ѵ��$G����)\�]��g<�G�)�*���u_�
��-k8 ���S�� 	�i�a!y]�Y�J�h+�Y#p��e��"��Q.�V����'A_�fU���͔�㜃�Sz��/޿ٓŀ.�R�t��5<a�`�Y��`��#,_�b��Z9" ��F+����	������alcdɗ�� �cX�$���� ����m��t /<͛���N�{�� &!��qJ��0N��W�
��$C�G���i������X�K��h�T=a���<�z }��.5V�U'��{����k��;	���]�H�]���b
q�#YY�'b��tr4�t�c��p�'�]��ٞ����Jt�=2
�ucϲ������~s�Q/�>�]cR�&.wY���5wwr6V�����FTX�7���i[��xE������Y�2��������[Fz7�-9�4�1��ۀь��.���e��$��H��w�� ����PK1ì�=ts�DT8N��F� K�o�����^����/W4���9S��/����R�}�ua
&�>{'���Ib�*#��NF�j�K)���`x���|S+�g�����*�g����yp��L���e�u��r����� �/��t�4���[dUߙݨ�
���'Y�R���^D���P��QX雺�h$�ؓ7z��UC;��D�$7�����2W_ ��d��I5���`�R搅��\UW-Z���
MkaYWv�9Z"�A),�p��,}v�g;��P�"��ӏ1�d ����m��G�6:r����.pi�zI@���n��������_�>�$@�^����ԍ���\I9��0�ѡ��7������c�+�+�5H���/ob� y�8��lI����k}��Xy�%�����i����_�������[k�_��e"���~I��ݖ�tr���
��\���[�V���%A��NJK�&���C��:��.��y������\8?cAoJ��Id�9��fx����_`��+$�fK���u"n2�F��	F�%3���@��K��G����e;;ԲfDo/���/�ǫv��ǀiCƇh���z�x&�V��5��� �`�ENȋ��4�J;`���]i�
阎<nL
f9�N`B��sӏ�Wct��{���G�b����^�:]���hY ]�I�8#��6�)��`�%�&{��$��P8�_���Dc�����-�S��!a��k�=�7��8�2HV	�kq�^D�a�Gqճ�-i}MYS7�"�#9#Q��0�����`�. ��m�o�g'��xC@y��}ʨl�nxy5Xl�V:���>�91�'Hj��"+-�i�m|S�n	��P�I��XaL�s:s^�hQ톚�A	��%��u��xbEb��t�7�D���x�@�ٷS�?��oIykq��ﲭ�� I㭆 0%a+Q�-C�J�L�[�F}=��Ŵ=&��2�"Y��#R����ܦ;�F�y��.�-��9)S�?l���ȿ���-ml��~e��긊/,5�E���q+��Jd|>ᮄG������&3��y�����+���͠j�-6i����0�x��|-� �@�'�E�8ӣ��� x^&,�ܬ��4И���I���,իI�\]#��U��m]�iW�p�&D)x3hY�C��K��h@�nh�K-�Rd�%����_ 	Y��w��O��5y�U��{��������O��
�ڸџ�e�isZ�b�B���H����x.um�"~Y�6�O(��c6Jp��� �<�T�ْ�+Чz��0�0����$����;	��S"e��ݽ`n���q̮E4����%&�M|��}���ݕ�|һN�|(�H �nm�����LE��7�h�b��<g��Yض��f�B���������R3��?x��b�9�P?(�P��_��Dc:��vB���ٳ�\R��6.�?W��K��_)�-s^�I�!_��H��)"Ysu%'/Q�XNb.��ȉ���s�P��f��*����(y�5���Z���`����iL�_�C��FTL�k����;�X��O��d4��;�֚Rg7r���u������R��I3ܷ=���*g����OiVTw��#�دA���:b��+]_��;�HMqι���R��ee�ܦ�+��Bơ�rr�o���y�Q����iÈ����ƶ���*4L�9*Y����<�gl��t�]zT��0^p�d+��a�|ez������\�3Eq;�i��AЬ٫-��F	����^�s���??�\���*�^�3��;GaxR�~pW�u�]��������ԔYX_&ZzOR�����Q�Ub~��c�����H���X�v�*��	��*�����l��qG���c��:�z�g��Z���� dE`�!�
��%nc6_��gu���rG��LH��ٙ�=��rh9�F��MJ �ۤ��6[΁-�_�$6���~{ʹ )�#�v<V~@���k�%/�����I¾{]��պV�q�ѯP^�_�AI�ϵy�b}�d���A�3A�{�4����! N��� x7�C����t�wƋ�V �m��&���\����ɑ�����| ��(3,����n��l7O�е=�c�_p�DG�YsC��O��I⠂�$Nm_b��GG�}���'pݘ�3䄋����hɘ�ꘀ�ȉ��SS�ˆ���-�^��88F��Jv��RB��^�S��X,�����U��B���P��-R2v��O	�5;4��<�����z=;�%L�2�z�x9&qZ�]@��`f��e����Z#����Ay;3Hp�m���tm�uc��f���Nu1d5uR�pwzt(�۰[2O�g�"@+M�
��a�)o��I�'��d6�����ԒVg���YiU<�'�<67��M+Ƒ���~�?���w`K��}�R�z���(V�+�i��8�1nb0\;B���V�"Vu?H�V��6pPlH7�9��}�y�Z�9��_W��3|��p��n�$f>9���*6u�d������f�7r����!��k�u��@�ޡ9�P���&G-1��P/a���T�~��x��j� -ٙ��}��~�.�Ѱ��$�$vA�������&z\X��P�O[�-�� ]�.�]_I_��!��X��3��{��z��_��Xȍ\��bMB�������ׂK6$�T�C�4;��\�A�ze:�M*=nc>��S�~��_�y�ι�&^�t����L����}�i[���3����u%Sc���t�"��^l,�f��n��\N_�T��]v��qe��ӻ7F���*�Zy�b9G�^^mb���^>pVA��ü�o���qb(�+d_3��+ӫZ5�N�m�r=;{�c(�4�X��xl���&B���޵��)�fz�*i�g��@��C�� ��ڂ�C̷ c�F�J9q����8�qnp)�`}�ǣ���}q��0��M~C2�Z'��p�{�F$��:Vo�۟�Oq�2	�&XxM���.z��1�p��A҃�)@�-Bpn�1�LQ�Ź:����k��k��ĖleF0m���;�\Io��L������h�qr.eV�ꄖ�8��Lk�VK�c�v4��m�\<ا��Q��'�XݩWn��#`4�؛O���-���3eC�c�Jj�Ց���w�H�Қ�ligk�#�~�9�;�?�ҿu��M�ʍ?:�:��[�p���j=�/N�?�v�a/����ZV!�)��U��^�3���{F��ګ]P����s����Nw�kw�j˵��׭!��g�<�l �[Rz��3a��]Y��#ѕT+ـ2A�m؝&B�>�wM%5V��WJޙ�	�����Nc�~+�F/k�׳�!�`.�g�����=h�����#J]��K~7�Q\��H�af'd��ޮ���R4��I�( �}�Ӥ��X_"�z�'|���t����U��#v�ㇶ��J4l �j�\���z7�-�n.��+��Æu>��N�D��(/.9b�f������P�������T߯�5j��4�X\�I�}�rǈK�]a�Q�0ی�NO�L�HAF���8�Tn�*S*$o�@ׅ��9�K���T��� �n�vq�<�xF	Ǜc�� ��j��ֿ�/�uٶ�XA ������ ��|Dpx���A'��u�ذț�4P��\�4��qk��HpO4�5�Dض5oK`��a?��3$ㅋ%��Lz�:�bǗm!�Uu��T4]���V�G3��Y�O1&5ټ3��i�Q�Y�)V�b��S����j����MM/���Gfz ��l)�A����B4N�!+2��'!`vC�����hbp�^�>PB�'�kBj��;��f�R�����}I�2P>`
&?fEW�T����6r�D�kOaD��o�R��%o&ǴE)��My�q3�S3!�q��Qz/����G��p�]��
��xV�F#0 ��:a�[�>(�;<�Jk�B�^�˸>�(,��h�C@����
�J�?�JTyr�+Z}���(��kY>Q1��-�G�Enec
���l>��$C��6J-t��O$(}�1��#���Lǅv�����kűL��!�w��P���'�-�Du�ܛ��l�u�P��X,bAbz����9Y�h��uY@������ŕ�wk����Z'�][��̄��P�t�{c:�T�/^�DS��G���W����ݴ��2�4-�?��S��
&�Bl��A=6x��DB�i�8�#?����(�8̬h
�e��	��ґN���x-Rt ٵ��͜���}��C�����i�3F�x�DÇ62߿�=c�{MY���a�$����IA�lmmr�$索BD]ꖄ����ft9�-��,O�����")XdYY���C�mf��&R
�y~��7���A�%qg1bdX����y�>y�[�V&�cl�J�����A�-�c,���E?M�|���nD1������V�� �G�=���lt"><�mja���5'kO��"BϦ�d"�9�qc���Rv��p���yY��FZ
?X֔u�hx�8���4��-���Y4�Df��H偋�a�Q�k��5} �lj���?��.�h(5�G�Y���/ug����~.�fˁ,�[)&���2�p��4o	�Pb%]$�:���D�]5��#Y�"N��P�7`~���Hl���.G�7�2u�0��}��b�h�����0](�N�u�cUq/@���Z<1DX�J�O�	��h̝���N��f�5�+�5^.��&�͎Tm�>�&�w-&�`��@H?�h���E8��1/|w��;��t�"�m2K�U��g$���pm2�ϻ���5�����;?	E��Ɵ�'V2��?�ڠ�����Ρvz����|�Ջ�`�ҧ���4��˸�y6U�[�����L�:ȷM9���=j�6j�&f�^��5de�u[���Au�//�|ܳ��ы� Ϊ�1u��v#˞��Ξ� yd�p�E���1Tԭ$���vq3](qpb���6K}�u?�?�:��No�H�Zk��HLO`����>�j�w%z�b"6-��4�@��7qT��R����HP�C��F���#�ˍy�����7*��|���a���}
���a_V�C�r&ţT���߁��V��	�~ ��lW�CKq���eEY�^M��u���粂$�s�)I:)�6"Q��$��u	li��&(M�b�u�_@���v�O�ߜ�qf'����q<F�8��7뿉~]6�����6}�v�f6E}hw�F�8��#T��fY���93��� S�*��^�G;b�F���������[5��y:ňR�H�2з�����hǿ�+b�Kt�� ��
��ꥫ�������l�*����G�1u�����׵�۱�"�1�:Mڪ��$�|wl��6��ݻS�O���c��X|��E?{�MaY�yf��`n�x!��Lټgt���7��AZj��x�o�t�d���}UMo\~�3[����Xx��	���C5e�,�<`>'��d��7���V!��W����� Z����i}�Ʀ������o	R�W�8]Ȣۈ�zKٟ�����c�]3���Ԋ�j���g�٦f���P�f	�ۺ�N=PQr�)�G�׏B��Sl�-TY��c����O�����h���%g��o|ƿ�W��Te��][��#��(�$�[I	�a�`�|���_r��3�ks��9���/�r<P�ۆ���
H	eu�
�aT�//K83Bx��uef�f�ע=��dĨ��<���MB*"-L^?ՙLBM!�n�=�.0�p$]�=&��U�i(�<�UtH۱���~MAE�����+�IQ�� ���8gc�F2�]p�I��C[ ��!!xWY����
�3��-��#�)�8p���K��ZyM'�	�'"Xug��1����O�9�y������'b�Q<�(}�d*<��d��=��k� �0R�[�����KƓ�{%d0J^$gU:�����q�:\�}��f��>̹N���q=2���T�����)m�[MVc\���䵠.�eZ���ǂ���%�Y�jl����kM���X��W�'��|����"H��)D+<f��cT�C�@��v��4��;+��޴�9#
e��
g o���p]��¯R��N*�7�B�l�jvdA��I���a"��Æ�4
��C\��Z7��Ďn_��H;WN��d�_,]11��2Uk���IYv��߮��2-E�9-E�Բ���,�ֺ����}���(�Պd4L[�0����N{��wf���K �����O*h��:y�#�?|�i�Hގ�f~�-�S%I�ܬ%�B�\W�S��Q�x��!�EVeBmV��UιK��M�Dz�5@sk�v����~������k�kt�t OrSCe��rH��^�9"�Y���}(���pgA�!P���D	�C���hu�=u�y����R�ɲkvg����Q۱ߏ���j��d����U�K�:�]�4@ŧgX��m$x�%�)�����z}�fu��C�VS�r�wƬ����
л��ф����e0�G\)R�ǳ?I[�8T�Xt� ��-bi�U��D����WD`��k��}d�h��>_HP�v1>CW9_z��l��YF1�18U�]��	;����Я���IY\��̔�^b8ү�V�[�{|l��D���.��N㚌͘�Q[Y/�1��'<	i@<p�0�fZQ�}ষK
�U�u��������Vz���
u)��3FC���f�3J!]홦�#��I���`ƺ������K2m����+m�x�W>|X�y�7og60X_�!(�-��$���,2�7�ˑj��=V���ՊW,8ᖯ�"�����L��S�$���w5_�c���c��5�9N�,�+:�"��0z�֙�K�u�Ď���ĕ�#�X�[�;?��R�_P{�M�Hb�QFDP:���R����U�/�䳄a_�X��>��v=�!�Z
w�YA75��7�ƙ�> ����mf����,į�����g����՘�^P�_���FH����0"����ES�	P�&3	��ժ��:qΤ|��T��#nF����pQk���D�=n��{ ���y�Ԓ�����y-���c�ʘ�p �����[2w*p����]��� �jAk*||��x���٬�X5u�=�K�g"Բ�l��|
����F$.s{:�6Ĕx���������F1��� 2��t�Kz
�4�V��r�V�H���[	���{X7٩�W�G���\ɟ����K����}������<��֎�0$��%ѰT��NDI�Fp�������g{	D3<fY�n3�_t��z_W	]-�F�}��>m{ ]�Ӆ��]����xkI\E¥�I.��7��I�ո��Ԛ�=�m�.�揳ǘ�e���'�u��<]h�}�d]#��0a�w�s�23�S�a��r�D- �"4�?X�6>�� ��H��50��#�M� BG(5R��3:�XC>s�A���Li��K�Ezg5g�2/�D��Տo��kS��N[�*Y��|�_�l<n�&�l�A����M��IC:�{��]\��]�A��@uamX�~���4k/�J�{ώC@-��ȭ�%���g������Ȩ����W�3�-����:4^��`Y@nħ����X�i74O�C8�{7�7OK�ww�]{g|�ﭟHv�>(�6�mR�9���T╳8W'EF����%x����杈C'Va"q���"ˑy�O5Y:�&����wrr��s����jpbe� �WߋL�m���Z�V�Kӯ��ڵ#J���I&k�t�h�&<Ru�|�T��NmgF��)�'��n�`)��Kyò�d�mip��us��%���1�rI�q��T�]��P��J��h��U��s#y4�{(n>�ۖ�p+�i���i�W�v����Z��/+�q������+Z�Y}�]�A���g���ws������S:��$�-7p�Q�ڙ"[5 '"�$�8�֓����_k�� E6s�Y��(5>�s6��6�d�EW�&&y>G���s�j��U��g7�9y��6�ݡQ=B����3�//���:m>�Ng�;�ܳ��>,�3#6(Y"�Te���mG�e�#�Wc �w�L�wq2;�������3��o�6�Y�݃���t]���<�62ms�{�6�y�tF��qz�o�t���'����.��ʥ ����7�����w�Ӛδ���!�=�`�˖m�1�Sg'Eu����C�a�(�ͣ�g�M�`bƓ��,,̰k�Q��E�J�,��ӄ���!b`x��k�v\�c۠4b�B�|�GR���	��М|�@���eTo����{�W9.@�=�;0~uB�]�#�P�V�@���+�����+h�g�a�}���+��_��խ&Pw*��*�$�($�A�^�ˍ1��*�����<�,�P�#D.�x�N��V�u$H�������x\���AaZӨ�q�A.��K�a��5�215�l��u;�aS-�N���,!��Ϩhri9�
���̂O{V3����n�[&Z�?ż�&>�|���n��k|�T�����-T�b�дw	v�}}���?1ZC����@�K[��6��9�r���ʅ���x���r7���a�y��3;������
���&�&N\���ᑩ<N����h|'p:��m�ł�
b�<�E���~_ 3��W�p� �g�/e@�u��[�d�7'c����h��ԃ�j}�,l����y������O�E3O�$���sNSV�Z|A�!"���s�i�ݩV�ܫ\��p���s��QI\t=$�EH�6ک�idpK7y@CI�J���l�=ȸ��nw��v`#�j@��G���x`�<:F	Ae��
�'���(���q��,�\�/����$��UN��`����+�Ξ{��:����Sz���P�f���)q�W絳�U$�g�os:�2�l j2tQk�W�݂��#B��	T�{�+Z��'�	�R#�gB�|���׮��FOܔ9�R���?�
!�3��CXF�_�����A���l-�Rh�x�o�7Z��[�7f=�f�n�,5�Tv5� ��0V]�j�?��`�@8�?�.��f����(���t�@����W~W3�e	1��v��8>���J]TE+�_N?���r�(���omO�N�!�B���ځ��"�7��e�<�y��gC�fjw�du�M\Kb��+p:�vƣB�}�B����~�+_*ˇ�7%`^xJ�-�}lV��Ǯݒ `�*L�[T�f���� �a�5��`����V�[yId��ķ- ۑ��h$��*
����T� E��� RD�� �݉]�_�����yc�?��D���Xt�*��7`�`��4����T#aR�|�mx����Ϳ�W�X��P4`Μ�w�V�vAq��tk�!�Le�Q���Uns���	�DE`�����!*#=9���|�x4N���ҾU�����ah7v?X�	���?�:�zЯ�4���ShHtk4j��	��zdc���m�Wa{�=��1��;=�������P�0C�N�9k�tg�Ԇ��l^�	�n�YV�'��9M���*EX��A�B�l���?0��*6�:�����RO�և]��:�]�������j䩬�� ����9�����}���G���p��Fƌ�Ԓ����^.�� �2�g�
��R�4oK��?2�q� ����P*l8[h�u��G-�8�cp��*�z��NM�)�ó�젲2��`��O}����� ��a���T|���ܸ[e��p�0�ģ�AD�5�跛7�}���A+���a/�O�◠S#r��q�����7;�W�'R\���_��)_塦̄�i�z�(Rm�Ol	��;����w����~`�����/��P��"��K�)d�-�)o,㪊g���ȉ�T�6���(�Q�(���uN����)�\��=�d�O���v)%*E�W��1�@��s|%��8�x��!�|�2�0�#��;s�+�0j ��b��'�^�k%2��^�[3A�7a�/����/�q����
&������Y����n���l����7� `�7*�:"1%��ډҩJŀiVP4�4�5?a?�U����9/�s��s�t��������l� O�+�<V�he�0�������\�rX��\Ӈ����Bu���)h�p�,#鈅��BS���M��9��/����=������m��4����$XPQ�R�pz��f �Q����a���8O�c7�Gwf'�m�pQ���_��%���#DU;�^ʟr�8�:����	��H������z�_��6��}�x��H�1ށ�Ղ�E�$i�4��>�xK]��ǀa�s���os�B��k����3���y&���� L�C��-��
$ ����7�R�����2*�魢�b� |sy���E��@v/K��5j���f�4I���?K�,w�a�AH_��!Ktze>^B�(�����m���ݴ��\P�ׂZ8��W7��:�p�p����E�(��ُ�}fw�1�7Ŝ�w�t��;zPz���{��s��Ś�،�X�N�X�|��']�Qo�iB��H'�+A���Jg�p]��}d���l�'����=!V^o�:����n�j�(Dj��;����Od#�
��ǜ��]���,��iz�9�pj�����O5:N�wt7Ϝ�`������?5r�&�ˈ��?��38�8�N�$ӭ�-t����}�΁d ���H��/�@d�o��ʚ�>!p��ō;'eއL9}Ƅ0tؠW���K�M�� ��F׺�u�ĸ�O�.�����D5�N�I���ySӁzZ�f�������9�<+8"����X����Z��x|�Ul�þܝ�m2�������m1�B6O�E{��W�9�P����?;����_9��|�z<��T�������Q�������T��na� 3��-�E7)������SQ6�������^v1@֊�����0̿W�����gl�sIh�C4T|B�/S\&0�0�
�aU��ѣL]�����.CE4^BI�
��O|+gd/��	i����NB�1�I	�Td��9����q�82S�O�麙�~S����s��lB�Lh�k��u5AT�.����0�Q�Ƌ7�}��w}�cY���5��to�Y�Tb?��6>��A��6�o����f-;�����V ���4cR�8Ы`@�m�X�Cd�Op��2~�l��|�1BU����Mtpބ�p�q�Y���,�x�"e�VK�-1���@�n$_r�"�g9{��$l�Q3��@����~fi5�_�AV��y��7(�4q��Qu���,�da����ُ���BR�:1�%I��ݬ��)����*�8���Q�Z��U��8	e�ݩ&��ٔ���Z��b@��
�\�MH�r3�+1����m.кa��!We�hW�F:D�g_�e�8�(EpP��Ĥ����T��b����	佾A�I�q�8m�E���ǇNaL�I0�x�FJ�Urj�3q���v��:���ڭ�-��!z�3h7ިlMNek�^�����]_�~�!��<I(������]XKt]e8_� ����z���T�y�e�0znB��8AϮ�aC�ڏr�Y��<�K����%�:eu���Z��z�j�����F�0�H�1
鐯}��xm�aԄ�V�����>��1��Ǆ�΁�;��0��s����n^#sԗ���b�|LƗڛ����Pԅ��^�?��O)�W^���+�Lg��=��n��G7�g����g���~����A�aC�B/ؤ��K�ϙw2ۭ0�}k�F����7���^a��YA���h���.�c�w�z��=�X��9d�[&F>��7�.������"�K %5�!�r:&/�)��s��6�[�Ւ_���� �֏���[�}Ó�\ԅ��Z��5�)j:�*�������{��+� _.�x.;B��`��t�炂�,!�;2����i��z�A�0�X$F���V�\�s��w�z˙uFC��g�������3x��Kӳ��7"���K�d�0B��(�gfY?"�~���ie�0a���e��"�i�T�M
��'~��b /�Pо��I@���jw�W⧍�!��`�11k�)c?�ܘ�j������V�ތ�Vf:3��V��x����t�i��?�8^:�<��v>oڱNL݇�s	�C�����$��]�xJ�Cb���#�b��<�ޠ+�����ȭjλ"P�D����$J�>Дhs�Zв��w�׾��#�t8�Sf�����n���7��i>�w���Ϻ"��P\4�����F8?�Q���LZg����P_���{���&��Q��Z�F*�|�o��
ZZ??����E�1�u�Q���CIGz��������D��P&�"Nv��#&.|،�������ϐ͆��������Y�����l�f�蹲2���T�#����U���7.4P�釭�=ۈ�3g\��� ffpߖNÛ��N&�(.����2�T�:��|�ƙ���+��+���<t���w
Ĵ��9�Êe�I�k���~h�G���t���Co�B��Mu#NM-�3�p�N��� x�T��`W	�p0�`���N�}��t�<z3ݹ�o8�Q`�M)�gf�Q,V�l��G��t��v(�T :٤o����b����zݔ�M&a^��\eJX��n�U,�3$Jn�p;J����H��U���Qo >�d�^	�Z,Lqf��<?��º�@����%�{�>�r )�_ƾ,9��
Л����Qb�p��}�ķc��d`�1�w�ϣJ��7ց^0�ڙ�=���:M�V5$�K�@����>�C}��Yq�w���&R�&'�Ϗυ�~�2�K�M���
����Ҥ/}E9�Tau�1��L���p�6�q����5E� ����t19Ma�1�BE�@�$���}�3���Gdjݖ��'|s6ӕ�?�	����S}�V�������8Y� (����z�ag����.��C���>�=�~�~>���ذ����s�J�-7JW��:1�U]�z�W�a�=FJ����ɫ%p33=���r0��Bu�n��WP[��U7�`փ3�0M乃�������*�7�T��z}|�g9���j�+�"�\̼c�+��v6r8g��$��"���Z�bC.�>@����� �tZ�r���E�!Qb+�[ޝ`�X���
�g_\�f�wÂJ�J?ݕ�`��v,ŉ��s��F
8�n��؃�\�֟�<����C%�/�܆\h`<k����6�ez0��6�.�y�����j 9!�����.����!�͒%��{�n�}�D� e3�d��|��ڦ���:��&��	Ǯ�
��������-�r�S,W)�N5]y� 3-8A1��@-txX)k���!��d^�P\Ah}�_� ��[����:����w$����U��F���J��d�ᏨƾY/`�S!�?Bu���T:}K*Q��K�a�I�QbI6y��ۆ��_&22j��MC�%���֗�+SB�H
�ePg=��hC_��ب��0_��w�츀������c�-6p��ڪ��.������D���Rz��"���Gi�6���ޢ37������H�#z�_����Z@���gF2���cn�1�e��IEA�o��Tq8)q؉�P����r��e�eΠ䃗�,����إ&v��%�����J�K_h:G�\L#�P�e9�aG�6zv�w�}�v�ifjj�J�	Y(F�Sk=&���(dO4���Z ����J�X��uQ9��-�S����5&5���=�@(�M�0Pl��豌�4�LM �һ���}��i0�75/d��\�
�� ��}�(���vT��Z�Ve_�t��Χ���C��N�/H��%/?�g��H���;��@�\�x�L]�^(;��ps5��?"L� ��X�����}�oF\��5��O�^5O.�<K�{�Kv�T�l��HI�_�Tq���ϳ�`�[K3�Y qD����y3����r͸I�x���ډt'��{�H��YjPNgI��$��"Z�ë�$1֟�������PL�m��ׅ�߇��C<n��:����S�U�k蓐����/��-���}���k�Z��`�wU�(mTc���1�a+Z��4��}?A+�p�V��&Β�m*���,R�����t��`�����c�i��H%��/�%���ǀ�XC�)@<X�8��I��|�%F��dp�#	"�N�_�l ��$��-��I�#K�>��o㠚���Ad��Y�\�?{�ܖ�p���H���FV{�gTϟ>�� 8��F�wI�XW����\q�u��{0�O�.��B��U�?X��;`�eנ㡤�~�?��R�u�꽌ְ�P�b�I!���L;|��ӄEq�k6�I���Tj%;hZ�c9��+3	���!u���b��C&��j�ߡ�ua�i$�p	�q�S�酰�m ��[�����8�
��U���G2��{��:`�0Q�� d(n�����&6eOHb ��?k�OG�`�n���Cԏ�$b�C�ʅ��{}JX8�ӆsKmh d���JX��[b�܍���p��v3ȋV��,�	 �8�'�:�7�I���ʐ� ����PJ�6��
�o,#���:n#��)lQ���n��H����btI�Â���f��kg�M|x(�����ۦ����k�kU�����L<���m��e+G0q}H���}���N��)N`�9���v4�LR��!@U��&ۑzxcC��1���9a�hĝIv�I����JN�=��,�;�y�R^������n�M��7X���ݾ�i=�UҤ��1Ǐ��/�D�o�fb�t�ù7Ր��q[gIG�b�8�iͬ�Eӟ�Sn���u�U�ګ��gF��U1%\�����Q�|X�U:_�N��c��芋s�|}��Tbh%5�����f�ZF�l��,�LC�n�++�̦,���o� 4���,t��Ab�!�`�4s��u�\>]�ϣ��MV���{3ӂ�@�������U��9�s��Ϟ�6]�7��JŐ ���#Ȑ�}�d�%��h�N?=������1�q+�C�Wӄy�� �(�:q�O1�/F�V�����q\�{��X���͐Y���������f��8���q[�/�����F4���E��)�g�(G}�H��<J(�_������٘cWbqL�¨���@�v���ɨ�50Cΰ���,�����	C�<45B��0���܄�
_9t�x-�̆~M�ңE|w���$�g[;���H�j�w0�s���?J�#1gfu�5�8�R���cb�&��%q��}xD÷�83�d�kU6Z���-��d���,]7�r��a3�E	���?��J�~�#��$ؿ3������x5wӆYᵇX0�s'��
[�na��[��}�	�6�U`�|�����ن�Ǆ�9%��֗��sWz}�������7F�ݞ��v�ľ���1�Jw}��oq�@.*���U������u$f���tZ����<ǂ��̈���Gb�]/h!����\�&Q�����),^� ��+;�zR�=��5��O�?L�צɢJ�qb��7P�t��,]�<e,���x�Aâ��UKw%�.l[	�2��&��b���0\���G���at������2���Y���!�v�F�EHꜾ �ܲ>��k\2b�Cᦺ/+��>�.�G�~�!g�m��	��PǓ���!�p�R�j=�U�g�)����M`V�B���"�W��nH�6R�t�2��!<�!�ofpi�}5��6�sڟ�E+�BW�RP#_�w�mM8�+'3^���N���NM�y*�`!����KZ��*F�P�Dt@%�O�n1<��+e�m;�,��J��ذ[|��Е���]�9�>���K�H?��Q�9�-�:�f�&�Uk&����(��.�A�1!l��oj�a�T��!O6��O����Dz���rY!,=�դԌ�7����RB���}���2-�r�0,eM`���/��P�	K�O��W.]q8�t�U��B�AEST�v:|���'���M�k;�^oN�C ףɧ�&:MTH����飼h����y�2���<X0���hh
��2z�ZB��b'���V����D3���E����T_8�a�Ә�i�Eџ� ����c�U�.�g�Q��LC��;�d�x���dAR�>k�*H��ޓ��� ��n�?^��H�K%H(���X���.�K����!r��F�,g�C���"������޼n!a��4ȴv�C��뎦Em:v@����%�������{�i�V6<�T+X�����0'O|X��d8ȇ�^��"H�ɘ���ɞ���ZB��a�1�@6O�h#ڏ�a`�<��}����Z��0��)n�o��Z�Mw�?46�O�Z�4��Zh�kS�����֢%.�J��|��)z9��9P�p����7�a��K-��fX� W��2������16>��z�
��k�")����k�Ԗ����s�sB5w�7t��ܨB�W,�E�Q��ײ���۲�N���HsQQ��ae�ˋ/����ǀ���O5��Up��)�<L"�<3@��)��+��	�L���\Y
��Jy�\���l�ReiO!t�_�p���xDd�����5)�g|F�D��w��k\�)��kť�̍��6���,�%27��>^!,:�H����ڳ"��ϖ����#���$���J��]�x�=d�B/���f݂R<�=�:��<�ܺ���K��6�4�[��������G@���6��ux��O�]�E���Pح��&��P���!�7��V��WI~{!?�}�p���h=��b�8X�$�Y5��{�޾��ÇN97�$A�t���t�����>�b^{��r������I��3��Is���!��o�T�M�V;G�/K�t��!��T���-�p���ɰ��`���֕�2����Ə�"�1�'�%���8y���oP��?�#���݅�%)z1�[�PQ���&ܖo>;7�D;g󱊉��?Z�}'���j�}�~\��nE���Ev��@)[w�Y��w�h�8�ђ�\"e[I�M��lW��l����D�<�b3'�(�o..��:M��1�q���2�F��[2f� X��7.�����ū�����HP��Qh
g2�0k�j+TO&�V�(�SG5}�^�*`���y��#�S&̲�?&��S�/_ő�$��@$���-��,�B�k�D���j���cg�#�-�'lu��J���5�'�y]$��������-��|"ވ��/`��2��A!�> �T����{z�$�@���+�P��~j�w��Z��Q��]0� �X��y��К^�����C��H4�%|�fN���A��a�:S���|k���sB�j��p|�L���.�k�ϊ�����WYj�:�{΄*��x����~��iK9�y�VvJ��4cZ{�9��S wkF��]��h6��]�8�Z1gBl���x�D�Օ#@^j,�;K#X��7��q�h�E�HF�7���ij�Cc{[A")p��<���Z��c��̑"&R/�3��-Ǝ�����`'{j:@yL묡`��o�O˱S$����*'���g����[uTJ��T���mt�����V�T�dEVt��Oǚ�s�w�ڿX��Gi>I�<Zc���ɐ2S�e�;{4���
ϸ�C�^� ����|�|e��S+3���6�Vm^��o;�o�'�ɍ���_�jw'ܙB'{� �z��}�hd�R�G�>p�N�m�Ʈ�l�6���u�Rf����0A��?���D���Ѿ2�h�h�)2��c���^���*.�F�C(�_ԃz.��-�u�X?��������Ki��nO�g������Z4��������PR]��)���l\$JKt�c[}�<ކ����� |�7��/vA���d4�s��MY��e�*��ܲ;/��#��3��P<�D�T�e�j
�&�B^�T�/�;QUb��j�(%-aIS���Y��"
~�R�R^�s�7v�b�)U]�E�k���C��;�	�mW!�Ђm~����1�.�Y0�;v��'�&�?\����|52�(���&vA=k�D{��׉�!s�-T'����M�@�X)>a?���;����˫'n�pHOR���49|drǵ�aVq�X�D2��K\m�fՙ}-��u����EV�  ���>�Ժ�ʠ	#�X�*z��4��>���d�a��9~t �>�����m�\?�(tgsNۙƅKݢ09Tuq�R�$̀�)�th����PMp�s��aI�e�T��ÐNss?L�\���g�6{`A�(�]Ʌ����z��͊�>ʷS})�=�������R����YyH���#�eެ��S{{#^K�=�	i�/�A��wӮC"�����R8��aQ�j	i
��=]�7\����3$�"s���DFbL$ �t���c�eo��lF� ��Ti�4)�����b��P�Do$�`����벋�r� ڏ�.gH�`�m�g� �ȸ<��p]"d���(ͩ~�O�\��g���9��Xs���|;���X_ʄ�ƲK�ZD��,Ֆ�b�������iU�~!:m�:�`����RXay"D��W۟(���q*�f�	.��H��Z\@~YxR��`_Z���L�>p��[�c��3����S�fW�����v����@�@�"��\pۿ�O�����|�5@���j�?.�NI����Γ�O(AX{?~��4[�pR�R9>^�)�LN�~�0=���+��<J`۫��j��H�<�_WK���T�_�y���;�h��8�aL��6 9�`[)4D�r�����v̜����*�0�d�yP�gu��	h�3?��q[{�#����S�H�9KZ��������bs�\�h�J�E���i�2�@�;ۙ�.��{����nY�R���;�$P2щT#	��?�������w\k:HPj i�Z����d`��	6	�5���#D������mU(�K����㠭B�Q�U���Z��	�
r�B��jh�����t~M�|�\y�-��!-�O�Qb�v
c+��N;�%M��֨S0c�oowQ� lgS]O�[.Y��j�X?��r4��s*�8ͷ�L�B�s��U��Vo������H`�������F<'+���c¨�~��"dѾ�c����h�|�:�℧��$A ��~��a���.4��QdG��4�'TS-�N�� �3�ѕp�U�o��1oT[�){D��t���������&��_kv��<�H�!�	H����u�1��� ��y�\y�S��	o���`"�LRF�Y}60O�=�,=O��'��+�Pǆ��o�������a-w'�����?���܁^v��-���zޱ��
�珁P� ���'D�*j��e7���U@�_h���#��x��3n�%>����x��^"�o����1}�Ϯ��?z�/��_�d��D�?���=�VWuSOrB�8*38W����;��Hg�o�ȭϜY�7�`�� ���<�bB��mX��v)�N���z	�����n������z��#R��Q1� 3��J�3B� īꑜW����\��r�i�7O������CC�f�R;Ҿ'�������Xp&���,z85��)��='��߲1;fq>_��xF[�:��J��^=L&��U`|�w
��S	�Ne�d�d�.�7�/)��6��*�/����&v-3��QM˻}zgF����#:]�M���9e�t�ƫ,!�ha��t�Z�C~v+8��\��B��b��倲H8+�� �qYvE��Dy�{��-|�
@����� 76��뢐o����h霛-R]����tx$C�Ы��PI��:��l/������D�r����Tzi�� �Q匳E�RIn��!�{�eP�>~2�@��Dp�����0քYf����@���^)!6�	:��yp�m_����^��2��s���n�_֖�F��\��Ks�
��;P����k��ɔ�xK�U%��gL���U���|��1��b�bh�����%D:h�0����#����0��0����nZ��lS���1�T,1��X���+�B��[�bjR�j�Ul�k�;�l�&׳��>\pn��'�)'�ʷ�P6�t��9�q'I�3���H�O�Z��^����{}v$��y(���NT³��ST6r�o�*ĚH���ՑB�9�v<�1sx�X�x���5�H ��Qգ\�k�C	�dt�;���
���5^�zc
�fP�8��}�Fďq��W�a�h3�&��C@��v�v�1����KcLm*�J�j8}����0���u2�\E������{u�a���7|cx�`j����ooG��`+-������r{����fԷOc�4�V�?��8�\�� B�`��{�|��(+$�Qg���B*I���}0E1���ݙ/���b��q�:���y�1�ķ%W�����I ~�,}�-�� O�Xz#��J:ԅ�:b]Z����l�]*�m��ʐ
�ǖ,Q��͖�f �G�R���aA��vt����	J=b6F�m�T�ڼͨ��[_Qj�����%�N�b����=�Oz0��<�8��r��3W�<!MH��|]��,E,��T��<9�q�F4�)x���1���  �8�qI�фw{�|~�+�%�P��Pq�1�D��_�=aHG�,Uqe�Y���U/�Aڦ�Wu8/q]ws�V����{�Di^@j�b��Tk�aG��;y��_��?�i{�od�On�<�l�.�btjY)I��곒������|k�؎[Kdr�����v�*Q��y������f�~��������<2-v�^��{�Y�a���:�&`�
�%��\��9���Ȕ`kB.��W�  kF�N���i3��<S��L�t*[��>M.�0IER��5y�(�vs�zIJ!ҭtI��l�M�?6Q�s�|$)ˆq���8S��=+ �<�
݁J�ͼ'	��u�Lە�Ԕo�
�;���h�����>.G@�t�����xP��0O�[����u��Y��NYx_jյ��9��x-���O�8�9p#��Ӓ����|���
E,~/�M��r�hg/����1M�x-P+�`'S�Y�|�X�K�Z��p}�@���A�ٱ��&ы�r�����V@��*�,7%ފ�u�\��?�N1s�^Tq).sQ��ysq<�,��p�g}W�e�^�d�1fGP��4i#�bhG�i2P�����K5�������0��֩9!ճ�y>��{^;l(��:���z| "�3 ύd��"��	���3,5��x{xk�*Qa��/����6=7Z�2S������6������5�	�?'|J�Zb 	;��r�!���Ch�Q����=�)ok������K������������q�G����2�u���{�he|���U���e�T�-f������Z�ƣ����\�j̈́�Kk���i��y��r6�Ӕ�{Y����SP=v�R��7���vm�s.�&�S�����lE�o��#��*{�_7�����~�<p��Qs�#)-lw��)�@|�XEG�+$��(����t��>�5zX��/�d�9�47�s	D�x���)��sX)W���Fx��֊<:��u���܌kf��d�a�9���FR$�dJ�e**Axp���F΃$��ºɦ�����9��t��s���g_w��&@]�1hsw/�@��� ��>����s��'��Dp��"3ad?-�!
N��Q���.!O	��C�ʼ�mB�Ԭl���c��z]*_�H��kGE.~�3¾=``��[��M�7<~�Ip��;>��1�qu��������� L��u��*��feY��?�Fr�_��˒���+��gU"���w݋YDa�7=D$ ȍSt[iYg7	��4	�q��R��WʷDjE\�t�9���1�ZP���Q&����W�I3~-�CCv���V���U��!N�$8ͻe �,�e��莞Hx�'��~�t�ִp���q��X����_4�\-N)^�R ���Zw?I[���=*m��	�8m}:,���=/�nD�|%����YwF�����v��&��%IZ��,�d�S�!0��E��*���a�c���j�����߿��g�~BVؾ!��=�������Zj\�☟�9���!��
�`(�Η�{�{!aK�j�t�2
:�(>dq�Aު�����ɇسѦe�QߗW���ϊ1C!��-stZ�ށ7��:��W%�)P�f�@�7g ���5�4�
��2hS�_�&NR�V������-"�~lD���
����xs�5F��4+��.߷��kv�h��4�����V��rM�p�u'Y(u���(�#��Ҥ���_A�<������g%$��F1�?USEg]�S�^Q��/j���B����q~J"�<�*M�܇R����1�W��yx�?�D���� �����#�`S3e�8��O�'G\��2'*�oI�3�v�F����㧅}�dg��u�9j
�|<�����s���7����q �
�.r,AR���0��%^��6^�q��������3�?N'o���M=���#.dt)��d���v�?�9������%����}�.�����XA4ʰt�����t�<'���OD��z��[��9M���e�K�QQ�1��軠PqA}h,|�m��
hX�?V�M��Ĕ���l,\:ݜ���>�W�Q <?;g�6\�~R�T��cq��r�G�����;��<'����<�m�R'��(��q60�(t�)y��k+V
ͳ���<�&����g%��U�M߲��;w0���d��][�@�2er�=�҆�Xl��$#ZL��9)�-ff�_�$���J,;�p��
d�>���i�v�sSD?��P(��� ��~�Zb�*�W`G�@k�ZS̐b74����C,BRi~��c�K7�<g�|H#��.O�ˉ��.m:���'�z�t�nY.Xn�?;����xm	�İĠ�'�yf�X�
�I�w�Y:����ڕw�׻I7̕����h�1�^+�u�ˠ ���d���3*�ߎŞ��� v^�uH]Fo-m����M�e(��RI��D��� _L�h5$��n�'�.+OW����"�TЊ�+�I��&�?��&�ɾ��`�3�Y�7A�<:�B <�7�ԄO��⶘Qg��%�;%F[Řf�#�1:&�c���ɘQ�tPБ��T]H�����W&�x�Op�����>��H�N����I���H&�,ՑF�ڊ�D��fR�@k���@a��'��c�w�����nm:���@Y5Qϰ'��p�Lm�Y�^��V��ƕAN�H�8@��i&�n��M�� v��6G�\k�8H�s�/��ݫ�'CA�W
O���ƀ�|�-����3�!oW�����$�q:�Q�W�ZW��|eG���붓����.�aQr0�f�k�� �Tb��,�&�\��� ��ILF�QП��tS(�~I��\:�z�"�edz�-l�6W���|q]�Ѡa��ZU�Uڊ���(+N}`��nf9EȐF�\;{�ﱐަ�ܪ|�/#j|�p��w颊7g�������
.�­���n��&�ro�p6�� ^���z������a���|�6yK�L{5�uU$/v҃/�!ŋd�a�`a�2 /eJ����F<�R�P�EX1b�`�;�� ���)"��2r=<���Li��
���I��ixX�!�&YP�ol*�"�F|�17�q.�Am�<�+j���3�Ol�8��6}&0�͐G4�Y*�u�!�1����d"0:�k�Fm�<�؜K�"8�$Ԭۿ�_�q�U�LlϤ����s6!A╯ڄD���6=q��>��8��8��;�18�ҟ���w����±��58��h�]�����8?6qqȣ��)�c�W�3H��\C&�D�䔚����^�K��q��*����TT�Y�^�9�����f�6ɣե=��	�C��Y��"��үQ{�"����tb!���2%���YxJU��|E����ז���`��~���i���?��Դ�����2[?�BH�Y�X2бy�T����n֟z���<����%!Ŀ��M�O2XR��*]w��t|}j�� ��ÊLѮ�S�l�)���*��|^�	Ru��Z0&���Pp��
h$D�D7,~Ug�����:Yc1�#;��ɣ8�j�]�E��x��̽����G
�T��^�ycx�9��E���9�Q
jC\�������d��X#C��jIY%֨���:��m^��D4��a��E(Q. ر�w�g=O�p?�<���md?u���4����v�Ʌ�^��ֳDb��4�8dU2I����H�>'{�4'axJ���5�H�yՉ���V�(S�{���iY�y���z����t��.�NǸB\��4�F��X���8��!<>���o/G�ɒ)�x��J�_o�I�3ʧ� �h
�&^с��C3y)fp���E{�`�
�&�]Ԉ����Na���?B�\*�b���}:g����S�%�o�ex�72��a�2����W~�w>�7ʝj"k ����A߯A��:4b�Ew���앞��h���'���W$rB�!_B�_O�%ȭ��'��L���k�}��62-���T��g鲅�q'6]��We_pS��Fߔ?!Mb�)���h�U�{�Ѡ!%�%%���v�k��i:i]7Xj��7�mW�Q��/*�k�� �����d�,���N'}�9��9�(@��b�_;�M���[{�jˠ@+�3M�╆�\dU�6���bL����j� ���f�ȭVM�eW�ÏE}��OL������u�,ĩ h~=9�j�U�X2S��s�&��$3E'qF[xF��0[gW�* ]6�C�<N�j�#��I��[��ש�fɿ1�%�يa�;cG��ʸ�[#4�!��G~(�������h��7T̩L��.H����C|WW���?��e��X��ٝbv��*�U14��ʛ���e,'1�ɅAl�9�o�6����5y�MsnRkRY��K�J�b������d*\Q��e��|��{�u��q���]�ʳ@��Kڏc~�J��I�?i�w�S��b!�hs�O;�9P�Z���*"�Y!��?z"���7VY>�2V���q�zS�خ2y �t��i��Xgމ���\���gT�4�W�e�9����4U��B��P�|��O������m��<����ߋ��4�l�v���#������֖����L�:�^�%7�IF���UA�ڟ<���;�H�t��m7�n��u�v��A�Y�*�v�`�8w���}���/KN^��:m-	���-:��!@���K�bH��^�{�y��e����SS\�s����1MIuCs:F��4C���&���aߺ�����p�|�>�o�|\������k?I^ږ!k��a�-=I3���[Z�⒩l{��Ҵ|P�@���diS���7n�Fy��O;���*�����笥bs߄��<�ٟ��0D�s��¯����^�����+���5�E9���*�/��X%�$�͋Mc "o��/���fk���H8�7��c���(����:
��Kז���2-�!p�
�����KG9�y\�F0��Xr�?�D��y���N��2���s��$	��	���AUL�E�"#&��YGK�.9��� K���u*�3��=i졍�m�R4�e�L�p���0�x1=42g8�ʯ�$��ŷ��j3*yҤô¬��lX`�|�|�>��t�D��}�s`�#�L+�F�
�p�D���r����:�.g��,�n'�(U�o{��1t��/����}���@�y~8#�6%gG?�j� 6�-|��>M-%;�=$�뽸���������Hf��0^݅s��(vo5��#i9��_���yd��bʎ�s� ��{�^�Y�jװ�lA��Q$$�4@�G��K�R��a@�`�@�F��~�\��	�{����O�J�lA�$2�`#��
��8@�۩oF����щ{����r�5�&!�/u��.�u��=�O�W�+a���;�ꭠX)���8T��U�.x�1�;�b}�@���9y�xֺV��߯��e��6Aʷ_^��j�E/9���Ĥ0�'�w0��sO >��:�N�JK�����f ��*U��U��Pq�)���Mr	u��ڃ���x6��?���f<���j]�_kS�W��?������CN��毄2�[3/Y�4�5�5rU���ǫs�m+HA�X@\�Z��ϡ0��Q$�͘S���5_�yMѡ[�d���<U �'m���+�Q�Vy�^��*\q,K�#�Xr���7��(�]6bA��h�UC��knћFg��*�o�/^f
9�uO�'��/n��^�R�v���|�����U�B J	���
`0f2�b�sV8�=���֛��`�<���G�1���$w"�nG�F>>�K$u��:�q�Q�5Ewt�O+b�k�卛����#�f|�b�U��C����M�O���v^u����{������V���I��8�&]�|�z..�c�����+��8$|d4���T�)��RxK8�op�Y]�!��~J1��6+};"|�N��|yw��KH�j��iB2�%�^����$����ͭ^a��)�9@����=�u��q��81����A��=�ԹQi���SG �c��Q:gn�f���g�r�6�RPv�p��P�n�64�'��EdM�1�yt�@��*�������	j�*$�\�{Ah�n �3g�g9l�ۡ�c���S&��'´<B����Ti1�w�R~=�o�ˣ��_Q'?(�.lȫ][�7�u�n��,�<�A6�ǹh�Ō���؎�����DT(lac���`C���j:��T�U2C#��[r���~��Y��m��Ӭ}ћ���:_N�)$:�|�����-���"��=��s)*��6�_OF�}�M�s�O����M����˘��f����/�MJ�w�6����b��c����&������	c��N��1t��3kT(������h����$�"�8Pd��s�čj���YT��O�B�_0�w��0�2�`��T���c(Xg�ݦ�h���s��ҡ���-��3s�� ,���f��0����_7M��@�(���Y�_�)���F��:�	
��o�ۿp��\�Z��ytD��C�u�3�f)Ǧ��H}`i	cǚ�[� q_�M��D������F��8���7����?����BB��|G�����i���c +ھ��qK��MI.֮z�F4��4��x���M!j�뮟{�� 3`��9J�Gǔ�²�5I[<�e�WC�R"FNk��:�%3?�S�/����eh�����;���>�ܲ>�/Y3�����ϫ�
�L��4�&L��e�X�o~:���?j��g|�$�J�NS$�G��+SZz��B� 5v��$�s�A��1�u[�X���x�aG��x>UɠG$Ҝ�ŀ��ݙM���N��ae���L��p-�6�!���>����6���G,^cv�t6cQ��Ҹ=P�����LZ�l��E�C|~��.����RO�}v�E���~��0�fr�뇠1�M� H����z�j�W������/?���
p��a>���Tè��\��I�g9��~��h��*:n�xV!��MTZ�W���{��޵��|�U�A�q����m�����?;"�]k�u�d��'Ҋ���f6�Bі��ⓑ�U2��|{� ]�!�4�C#��2X��D^w�B�2�y��{�OD�EC��������3�!�h����a�������<{v��D����3��M��-C����|��	�����f��प����Z0�*^A���������F�9����RY�f�Y;t�Z!UZɑ����PkE8�PT_�=Mu�O�;,�I�h 9�utyz2��)�W'}6E���to�k�Ő0�gk��y��O�~����BS��@��B�0��~��I��w����N����ɭ多=��,,�f�O4`8pЧ��r)�ȣ|,�͈�e��_�b�Q�<��e�B�T��7@3�n8�O���A��~�dv$8�����ܻ����v�9��<b����h��i��o�p)cp8롽�D��P�z{�U3�ҝ�h$��8�RV����t�"�35��@��"�	[��0��1�Ҍ��D&$I�Rw6��+z�^�O"0ݺ��B�	�#z�J2FG�۷S�9����r�{�]��מg�F��17[�P��觿�	�#�P�Ⱦ��K�FK^�����g���<y����Љ����wKTC�y�8���j�&�	�<�/��6���9R�	 j~@�,<w��`a=�?��g����2|G\S�f[ߡ��{e�����OU�lVX�x�bE`Ԟ�xϹ�j,�e^Ə���n/���m���U�	��,hCv-�ƽ{tA�����f&!�����9�{��1(Cי,�Ț����;Cѷ,Wb�/��.�d��&0�����O����r5�i�P�i}>���ݚ��_%��y~�b���$ų�譅�3[YP`0��y�eIW�%8�׮w�(�M5�������T����ha>\�l����ԚQb1Z����!���9�T�oU��^M��T9{sM����CvV0kI�R�'���!F�F���q�qʗ� %��E.�#��x5��u1��O�#�뉗0J�vL!�{k�E��*�`�s~ŇFd�NΆ���L1�_2�D�P؄lzV�]���0�%'5g;�l�\n�ptZA1����u�e�N�MW���T�O�e��7R4��4��ee1Y�ܚ:�r'�ː?��x%��&�|r[!v�j1�竘6�V7����D��Ir��y�����9��ݡ��'&s���h�aa������������_qG�M hc��Ƅ�{BBL�q?i]=H��L�)�֘��y�w�&����Dm��p��?2��M5_�#�(�}��k
�	A/�X�P�C�#.�j��X�@W��+NQ��D��� �c~'}����l/���U�>N��~�Ѩ��K�/t�C$�w-��8�P��F﫺�4��@8+�\`��tg���\&!��?�QJ����V�a�3�Edi�Q?kn\��ٵW <��'�C���VGg�~K��F���$�m�=ޢ�OQ7D�\t�mX�IܧX���! (���/�u^hD��#��-!�>�[��8[��K7�����3X{�*����E�2�7t����l�=V �깑n��^���]��=:��DͶ��K��Q���{1�5��#��-*]�=["W]��E8� ��(��[F�	1�1�(��b���8�x6��	>���y�̵� ���Ex+,`�q���fJ���Ge��j�~�1�����:�k�j�u)Po�2�S�<B8N�w���� ����C��7��;���d��~���Rwl�A><�O�`&�3�x0e��d���)A���.���"�>v���~^5�nͧ'��Y'�O�;�T�(L �v���'_vQʖge�}��-����H�Q|cVӣ&��ֳe��s�C����k�pһoP�Mi~�j�U��j��_�48�GS��-cBQ?>�4�[P��W΍�ޥ ���l��%if�eB��nc��	�R5.���|����"�%�޳͙'�T���0�L�R��;��FS
���2pc���0d�A�eٌ��^��:�Ƕ����7s��h��%,�����\/Ѻ�
��,���ڽ�p}L�dt+��SЌ�ei�E���]i�̋!��&�V3\$�f5տ��ݘЦ�*��n�y�
���R۱�:^h�VT�⏓�A�"oZpL&�
���>):������@��@��N�W�=B[3���$u:��B�,.�<8���Ey���aʋ�����:�����UU�i(���KwRBgN;�z`^~�oh:�4O6�bBw	-��d��K#�����rA���<롪������K�i���
z�z�騍?}N%-�����|��LAe��u��E�o��4~̈́v��Ā�oF<�>Rk7��1�x�S�����H��W�W)3׀[���%�g]��C�/�Mb��:�ܐa�h�HW$�|����MU~7�N�@�U���y�^gb�hQ}��2��M���e�D���\@�Y龤J��c0�5T��Z�0�s�躦�\+ZWVt[��������1 �k2��~�L����8$�����	[L�^V�u�� ��O�L���O��o��^�Q�������e�u�T~�9<�� ���;�ſ�ez(ŋ���宥�X��j����>� �p��B:�e��6��S�I�+;E+ye��0�@��M������|HiO2�O�#�)II�9����Awzn�xfBT�������<W�?�p�h:�|_�%�̡�Pͥ�iԕ"��:pS ��p㼥3�����b��LK��@�KA�?>p�]Bw�^����������{����)ls[��F��K5t��}M!R�hH�G���>��#pH����F�3��`�ۭ��K��H��Z��Ś�����ďš�c`[%&0(��QQwUW�he!�n�����O:Dސn��_�β+E������d�]��(ܒ�$�*wr��?:,��!�a2��}���t�TmR��ܾ(���U�����|��$��3$o?i��\g�����ො���Py��o����a��<�i�e�4��SY��T�򊄑$�y�f}��@�|7E���Տ�i�������r_�of�򸃫�[�^�LQ�0O�w �J7v�g���[��\�28p�����Iޅ��e�A�Ԗ2��<�(A#��s�X`?�LHq��SX�YZ+�O�u�?� �B�ݞ�!F�/B.�O�|�e�I�"��TPl�3�$M@����:i~�/0��\@����M�����'��<c/ܽ���^D����S���<Tg��^�MN���]����n��kG#C��6<�������hC�6��=�oj�������� ��S���B�I��ר�2�s��A1@灩XZwz��b�ɑ {r��2α��3�r��#�DN.A�da�p������l��JᎾ��d���D� ���r�Ր+=�u����Blf';���똦�`Ë ���Ɋ�66���^G}0�$��{i�֞"
�j�e�Q�5�Ժ1'���͙���#<����@�Z릍�S����1t�o�|�?[���!֝�px�`�z`�hc>���	��aJ�MՉ1�do��z9��=@��)�!i*_[,P��MOB�h{�>��:�o�;G��Z�(�'b>�����H���(���z�!���%@��g���90�/����<O��b�b�ڽ��+l��Tݠ�فr�%B�޹q;Gc�(�����`uΊ`���r %4&�� �ɟ�R�Wm�	҄�!v�s�����G��"N�.z@��1FV:�X҇79�6�RH{����jB��Ga���]��ω�9OQKloq�'�v��[��y�"�=Ԋa�ͩ��(�m`�ok� ��bC>�5'4��x�H�+�Z3���'H�Y�U�.��zd�P���X���l
��Gz�1�4�1�� BP� I�>�0�;��",�_�"cvI,F���J�c�y3��̉� �j�k6 �z�����B{�[���i'�%�\y����k��2gCX;\�=�:����p~��N[��Y�"!�G�p�@�2*�ũ�e��A�:?#�ܗ���L�x�/�M%�?��Pv���hzPB_���)ظ����C~���f �}�U���@�tN�FA��+v�_��R�:aǥ&���8
��]�\�q#m������0�Y�������<��NPn���y�����<m�Uo�/(*�����XUR����B3D�� �T�Ԭb�1� q��4����f�c-��Q�$$j䤉=:�눶�x��]%�_�k%���@9��)b ��
Գ�H�Y�Dt�׶!/�{+H~�ٙ��+C�[Z s��k6q��B��k��Ի|/ӏ�Fa5ڳ[��R�D:1���xv�����1�  �;+Y6�|����s����k�iH��ޕ�6tR�����Z��l��ܤ��l�7��ks9��"��D�Vd���₹ S�=��/�0�&&�o��4��!�,6^�p���ܩA��N_#��^/v��n��X�bX���<0(�U��!u�G��ӟ:SG��#�����e!zgej�{�ʯeh��|v�X}������M5�Wx�P`]��r+��+BV��h�.��yGa�o�%e�&�,���Kp1"����zq(�'67v�9��ʹI-�u�A��<�gSi���
DB�"����;	�� Vy��(��K��hns�/T��t�`P��.g I���	8&^�����bb�K�I�u
�-�龤����PF��&��e��{���x��z�]��� :�*��8��+o����f�	�&졶�~i:X���X�ly�|�,�S%K`-�t1L�F�+�H���*ت����;Щ�O� �d���ss���ZOh,�zr)e��A� ~a���h'$v��,��
�h�5L�������i��N����T��]����8�P��5�
>��1Y��HX_sq}���>�frpUVa
��AX��N�慠�"0R`>�MXMa:̃�i���3�ix�j"�����O���_�rq�����pR���]U:BU,����s	S���.p��fޑ+�#��O΀�$�ӏ����5�$m���-�HB���Q��[ �1S��A00Ү]���l���j��g���#]�X�1w��W��?1m��!&$�MĽ9W�^)�,�I��l�0��b�n�K��_'���=
/iw��ܷ?�}���OB���KD�(y��}��Ns"�٬p)�^�O��;\3i6�@V�Ӷ��Ă3�)��W��j�E�HA��j����YoU��`Ar�4�_�q:/�w�c�d|�V�Y���ףv�5L ��X0�����*���Z��~�� ?��eQ6����6� 3������˳'�_���H���݀c�?X6¦V�\b/�Sn���EO�hߥ9K��P���;2D������Qoi���I�<M�©����F6~���ދp��-�@"��.��`I�LtH�Q�G�%���ѥ�W}Ď�2*	1�G���p��_��e�)������72��躨7�1S��?QPC$�ݢ"�d%��!l��[�C4Ē���ш���IO�c��L���FB�H��d�Gpr�>L����R����!_�h����� D��N�檯�H���ւ�n!2�B�xד����ޑ�:3� ���/���^y�V�4Cĵt���S��ľϠ���y��Y�e��Ğ+�pU0�Z�nz�♟�4�*Tj6���x�;�d��O���i	��C鹫fSb�5-�E&���KO��	GC{�%v"V��!��R��te�*�(O��di?����@�뵾�G�+��+���F�,uW������f��|,��Q(B
Ǎ�cK��G���t=z=��TF6DFI,�b�����K��c�������^6�u�A���.�ke� #c�!���7��4�-03��tkDTk:	�s���0��.�ioI�rCH�tI�ǾiP��{�`�%6��}��I9�7�����I���h�"T2M0�0ZE�C�@���c{=����Zׯ�A(7]��a
a����/��<](���0��H��`Hq��V�&>���/R�w�r��%*M�/��Aͷ �@��^��B���Q�4����D�qa�X=�[�ڡ��P�a6i�qexɘgM�n(��(M~�u�c(դ����Ui(OSi��S���}&r����z��z�d���8֮3J�;"�t�9�o�
�f���>�7����� I�A�C��4Y���c�4ҙ�|�y\��:�욽��d�\��S1���]�J]�*�R���S��I�&���J^����-L6��W��y�.h���~�t������v�7�`9q��̐�T�������pED�n�y���� `�~xO�s�������1�{�gF;��ϴ�ċ�w3� ��"���ӊ�Ʃ:��뾇�醞�1E.~��R�dn'�T{�=�GP�ۇB���W����{�:7�hp?�8΅����	�@d�>�+�t�8���()��#�B�uA��o�=L���"j�
��=RSw<�ۣb�o�j��./�F���J�.;�)iE�+�v���~q �ڿ�w�<AKq�=��i�3�#��w�^"�1|ï��N�$a���sN��F�!����=��C�yIJ.��'8a�l�c)����q���yE�w��7�wn/�N���Xl�:]S��C��/��P�v�֠�	��/��<^��S�2w��]N[�|�?	ȶ��}#��W=#��g�4Q���g@.@ǿ�6x-�Ym�h`�ܞ�r�p�U)^I(��{.�3����7j�K��0�qņ�ƍ�j�3���J�\�ϣ�Sl�$���ovr�X"rm��hH�2WͿ���i�.�[��܆�U�&1�*�#�'d���h5��%���@�2C-�PN�騖��g��ŷ���L0�N��qo	���9�X�̝'7�X]�%o�bO��u��6jF����۱8��y���4���t���/c�>�Ӫy��������~��%BR���߫|T]���`��d��uO��J��v�ş���(��kȽ*Gcp'�X��� �7@Xђ�w�%�F\�۸���B����(w���	z¶�9oF��z�i>?H$�e��I���Aq�*���`�M�=Ӂ
i�Y�B��Yr�)Q��/���@f��/��e.Ř�˟,��	?)R��ct�"2[md2z��og!�Ҙ����W��Ȧ�n�u��=	���t'ŗ �_�B�zgL"mC+�f��Dk�0�oU���"˺���O���?���_�k_H{@�A�$q���&��EZ�՘��q��&X?ap~ER���>ra�W)�Y�: ��W��%[s�_�ˌ-S���Z� #X#�C�O�虞���#f��2��hݘ��O����o�P_44s]��2�zr��@-j�>h�vA0n5~�kf�VIZ��<�(3���|��I~1Vq@�W.���q̿����b��Q��y����_�����9�f�VX��oٸb,�G@RWS�o��D3�=�?��/w�,۫�,f%��_�����n�=
�Q/�!$Y$V�3�	͍
����`�)�T��ļ�v)�
�d:�*�JL��~3��3���蟾���Vݑ�Z~#3���$�������Fc�8*;���",D�G|�^�Ԍ^O�yU�����g������kl���W�/7u�R�u��ہuZtr�l�8�y�����ת���ϝ��'fKqD$��CE���=�
�!�|�=F{�������p�[�eΨ�����h�c�f�R�Y��Ιo�R\��'UW%l݅�����qS���Z0���P�ΔHk��Qp�L����o�?QB�X�%��IU�n�&�ѢJ*�2D4��ep^E�C����Q��Ralo����se�*���J�'�ڻ&;4�\'p��Ҙd��[I��Fz��v9#�l\:�@Y��oo���b�:��������22�Ƭ�N��O�5����E!���v�+P��
���WLv�`锄4-�F(��a�y�F��HA�����^�gIL��m`�V�4� B�4v��:�Ӑ�x�Ri>�u� c6�c_����4a(�����2wC���3�{������1��rB�F�C��u�����.�W7��6����4(�J�e��CƯ��(+E�N�y���0��2Fb|K���+� ac�SS�6�(�%��#)c���D1%u��ld�x�&���t�C�� �' )�E��\��M��1ߗ�V:$J��Sσ��� ,�mE
,����L�S_�?��31%/�@^Fv~_�&NM�f���X34	B�@--��՗?� ���8<��l&&�����w��ˌq�_?�@������,tex���}����{w�����ݠaI���Y���#���Ww��̖,�1��T�L㰇8��	
�ai���d��&\ j���ҩ��*~+���;�V��Od�13VM�����U����AX��Rm9T���G<��N+4�8�VYi�}� y����f:+]e�v�2�ڭ ��1�t}^��P��k�x>�tB�E��|�]|�B������ma�c��wK����m�z_r�d�Z�ѻI2��s�Ok����`st"j�Hy�m�l�q(n��h�߲�<�sh*�z'�9�.�ę�a+�񗍮'�w�w����k��������L�czB��h��$�U���
��g���U�N�v�ѷ��8R^rE(o�Ak��W�y��P`W�'�����pi� �����8��gS�`6ԗ�	���{����B��b�2%o ��xu��h�ܝ(���,%9�eX\��^!AKU`9�����
��1N�n��gM�l��Չ~9��н�汧kj�q� �?�"܀	�yO�},l?hWy�p��%L]8;<��ߑ�&������|F�D�2�"G\|??>�1��їU�A���뻪�R�U�}�{�B}��XA�d?�˫��%�� ~T[���$;;C�+�k᫝��~L1�	��q��2e{��~ �u�$O`enVV�U�qP1�q��(�!.QyO��m�����E�U�uݏ���^x>F��l��L�7�Z�z+P�$@R[z�\�-�:��=';D}�	��#[+�4薆mcI����I/%��n�������j�?>2��p�G:�V��m�I�Me'Ќ@�6阃|2�Ϗ����Q.��Jt�S25�2�,p��\���������$E��3�S�A`j�a�V�kt���ְ24�.�*�DA�z��<_�G��cƵMǂ�9E���!ZL���~��6p��z޻A�_���+�~�;��s��ٚ��:��G#�D��	��R˔M�.��<꺚��������ҬKW��S���꼐��y(���c�<��d��1ݹ<[O1�]�"��Z���(^q�47�,�ϖ7)��g.��%�g�;���[�K�0��ef^o�E�z%�k�EA	����� �N���}��R�C$�*XDW����]<,V �=0��m��^�x�;Sn\(d�A�[%$�Z�F#��6i��'�?A�}��L��@c�'v�s��ç�d�� g 5��[��a�)'�M�|#1y�*3=�F�o;} 2S���hHB��K�%Q�؇U��DC�Hq����YHJ�.�:-�3<OY̨5T�N.�T�Œ~!TV-;Q�nM�ԑ
����Su#�]
�W'��������HqQ7l@������5^����� w�Qt��#���p�g��/|.���*�-��Z�U�8L�M�$o���e9M�!\
�^H���p�"R��Gv�� �,�P�>�6�)�q�����Y�Q�R#�Ex1�R2O<�2Y� 0�S's+}+dD��Gq�'��S"���+x�E���ͯ�"-��]��� ���l��L��P���9Ά��G���������T�Qh�)���H�T���[�c[��uǏtG�쨲f��7'h%���]@[u��Q\o߇�D����}xV�i�ʊ�ئK��� v`��4�H�;S!�#�ܶ�Q��hl5��:��⩕9l�]2$��đI������DH���6y��GM� o^)��K���@�G��̦d�Kf.�}�WE�L�o��:�&-o#N�}�{�u��P�O; ��_���+��ۑJ�G�g֞�MB5��$���S�:�Y�uE�q�*��Hg}c"�Z�c�U��>V>,m�w�R+מ��#$p� �3O#[��=^��^��G!.91.^����N��r�1��j+��jyS��r�r��k�JO$1ƬT��A��Al�����%<H���9�<�B-,�����E�!w~0�5�¾N�h���Ce�K��/�h�?��R_�$1n�i��O�?�b�dN���yH7MLдҽ��A�>�F[�����j��?�N��G$S�n����0;ρ�Ӛ��
3-�YG7��N�l&��[ۮ����W�/�q�c1c6��7��U>N<8��ѝT�#��&�w=ø���]���F���(�>t��A������	�d�E=�Н(�܈ǽ�L$�Ȼ"�M��a�)��D��Z��%d�*e�nz.���p����TiwNKV�Ԃ����Y�3l�1�~��@,)N��w��bD�g�e��:e�^���荝.2��q5�:=ܯ�3��u�͎�{��@�o`{C���w,�'q��=M���[�eT�/@$A����(�|���|�;�Wne�	̃��j�S�Yi�pbӚU$���V����\;������V�G�R/ȯfGB#���*Ş�f����pU�%�k�t���X�ۂ�����d�F#<{�Ż2.�@?�뷟���KnPR$l�D��W���6,����{ٷ��lR��l�K�/��k�� ��!i����RYO��V��/T�Om���jAC
�UhOef3�^�S�.�Ke8\j����X��,�v%#]��T���"*Qޥ��x;󁲰�o^)u�is�M8P�l�����b�䦭�\5Lj"umT�L��9E�I#ti�<�Ƒ�|�u�2�;�����EEx�]��u����*,���
��ĭ���μ�Q~l"˭@P.�V��r�K����;	_q*�qQX��צ�o���Ӿԏ�7b���E��_�-��T�@��g"�(&(����b��s�F�p}:�l}ژ�U��u�m2'ß�(7W?�=�lv�-u�l ��l?���_Q�qiv�.͒S.��9e����P�?�N��Wqz� �D�|�+{�����/�u�,��Tr#AG��]�b�'���ᖘ<����>0�?��_��m�g	T �:��KI���M�q�a�eQy|�A\u�r:��3L �K�C3��J�<Ӽv�Qa���D�?�lTX�X���{�#p�Kͯog�HW������%����XN�A����t�̿�xQ�U~�X��l����T��G^��S��u}c5o�L�V:�}����dR��g�	���)J>
K_C��P~;)ޔ�Z=����$VYܽ!�=Q1��+�>����j���E��W��v�3M�v�|`8B!���fp:s?��K�ו"u�ZK�4�,62���|<��=B�Ĩ�E�eČg���ƶڽ,$��6cq8�.i�4!@v��ڏ�M�>�C),aj��%���z;����x'���-z��38T�5�@�;�E��zT��V���q��/�H����z�� ћœ ��+9/��(R�:�"�Ev���rh&'{{���Put����<��t��S������v�*�n?6�&��TJ�OE�Y�J��
�MI{�\�>u�Ħ��=�|�G����@)�W4`�P�tB��KCǊ�͚��k�y�0z�#��?4�:/�kVcm�����Tc)+c��aa��H��ͷ�]I�?P\��3x��''��5r��_���J�O�LYَ�̐T��� �V^M�r^�wLM���iu~V���Q<y1�8��pp��H5oW��w����V�G!��B}�������@[�5m���7�	��^9����*A���]ڰ���^�������P���(I����F���|��R���A��+68I���n
�`�![[�~zG�/�ȏ�!���;�]KxbNL� �l����k��Ӝ�Ce����UU�~��:�ώcL���5�9��2�uیr�}3 
�'>���>��FL�?���HG�)�ۑ�st����>�
�+@����0�Z�F-��.�B
��Xy�1�W����1y���dr+�M��R��P|�E�b1�Z�'[�p}q8��o��n����b𒳻�tGv�J����(����+X���:wwnRO�/G7�U��2���x0�w9k�>q(m�b�i���M�b3"�4F�B���)�����:lR�FN���1�	D��쌻ʗy��U�mP����P,E!1N@�V''YT�Z>�ZVN[O�-��zW�T�:�T����AV>zsi)�f$1;^-aO]��L[�F��~�f��@ĚJ�1�3X�:���+mQDҼ7a�9���"�k����Ʒפ��0�l�3:���D����4���>�����`�p�P�'�Ǻ��B�P4E�`e�����-2
C�Qc���䇮.�	�����~��A�֧�<-�7(����kxkL�`YXn	��'��ʉ^-���y�*W?���Sa6Ӛ厰�q�iZ`�b���S�|I���$��_ؐ��Z)(�s�h0�l�_��S�| �����Xi��9������}�mܭ}�w��`�R����Q3RB�x�Y�#������U���.�)��Q���(�\ik˥�'Ś�H����zd��*�i�ßn!@���72|)i>�csg�R�������b�/��|��)]�Q>�\T�"гݳe1�ږp�)@U�c���CsO�Oh�j��ZSy�.�&��zݗ�E���?z�MK�8ԙ'o��6T1H��6/.Vuv�̩��Kz��9`����_�/�m-50�tP���ݽ�a�(�6�-��=��&�wd��#��ᣛ�:h
�o�Uq"E�Պ� �,tZ}�D���d�_�-h��ٛĆ��p����S���o��f
f�S}��D��=J��*�x'ic��9$�X9M]���(E.�	Fıu�-�g��g�g�G7��g�F��2�ٲW�F'��WC��	_��C���-�����&�j�J]�~�D�zWܖ\��|x?�ӳ��6�Δ�x�z?u~[��҆s�v'qп�4���A�2S��^r��^��xeU�wT��nV�ֹԔNW�g�0�<W�&�=lֿ���=J���g,U�5�/(J����0��{!J���I�B�"��BD�8џ�V� 8�f�6����]G<+�{Ȑ�??"����f�mOf�zu`��? I��$��qJ}�KCŖt{)�`��O�u+E�@#$3ũ��f�'�<��D��@��?�[�ɠ��uR�zn�����kB��S�wˮJ)��A��;�$=�G-}�={�F`��Do���ڂs�_���M)�d�S
�4Gj&�d �����~�E����*"�ʍ�7+K�̂K�i1�12O���c�~�8^�ЦI6�:�N6<��!��L�%6֊�i3i�z8j$��J�z��Ð�d��1o�s�CVlj�)7�9Q��؍�C��>��K?Ч�m���Q�!;��Bn#�Hg��f5_B����-偀����gFf[H��G#�-�7�1�D�3)��29�U4騂�yg���V6
�q*�a�0������Q�$��w4ٛ�.��c�vu:�6aV�r1����rC�N��!����e%2�eb�᥊
��4ա�{ *��K�I���<d{��n$R"�X����a����p�ix�)�h�z��G�@�	��S�d�8���F���� >	� ?t�7e��Z=�O����#C؁�0���J0訕��:�-o��������2zŷ�J�� �	�>��5��7�7T�$Z���Չ� qw�yF�*��do?��ǅl[%�(��K >6�En��B�����S�1����� �����
��?1�T��E���2CF��3�cJ����E�-�p?�Z����p�����)F�Gxj�ZĜ�"Z�r����ߗO�G��'#`�Tv@d��[��4��[�m&�4��� T5�Cθ�d�l�'�k���n!�>]"ı�0}����9sɸE��,0�c#�f����Mt��s�4��6n�~�~���M��3�'
��έݹ�$����T0b� v~@���K�$�	j;hrE�E>���@�jt�<e�7�'�@��)�)�,��JU�^` ���,��œc|��b���x�#󷙫SzH{<��C��]�������z��)�Q/ ކ����F����×C����^��^�Z�^{f��/SB�2�<�K���}���C��aO�x]9S[��:ԭ0��l�R��u���'ѬE�%=
h��j�s��GU،�k<��P	��u�O|������t�kꥮ�a��Ǐ���a�,
 f�i[��>T�2�h�M�끲��{�e�6�@�|�e�qQ�%nזq^u�JR�q�ю�v��}��� ���4>��]���Ɵs�:��)��.�l����
GB��`�;8Dk*������M�
��نH��̢c�U/��uܷ��A�)@�<W'1H���䪏#\�/�u1g���{�@Q�XL�#�Ͽ��lg��o�1����'��4�X'�-��8�ߧ��Ӓ髦G������b�ԗ��G:�C����<�(�=��j!<E@�󆷑�X(�ۊv�S力U�ď�o�;#�D%���u���zUx[A�-�Aev��3�õ��&
'���X�Z��d�+�%>R�y�ob�wR��<���4�G�tK�U�ޝa�C�R��cȇ=bke��F!�y�)[����VH��B>�96�xV_�VPC�x�M��T/w8�q�=o;c`w>G�o��Q=��2S;T�i��o���R���SJ?�Ա�fsݩ"E��R�\8���n>�]�lc�?���[ꈇR�K����މX�#�YR�S��\�t���mL>�6����w�V ��4?a�|�dJ�f\�K~(�$~"���k�"u�ܶ55�O�@Dl���mDG�@û�mN&s����4a����q�Ė�fCz�e9����սf^還���a%8��?���M4��3���,F;]y���p~����A-�>�s��	��g{q�}^`-,�9Y�K=��������"�!�u�Jf Uk��~�-�*�ב�z�hj��W)�7��&W�u���	��u��m+xd�'��~��櫷�@����a&>4Ñ�Q'���+�.SCm�a!;b5��m�`���W䍡#!��\�T:�����
�$�+��}���� ft�Ӧz�zE��]�6��#��#lf�9�ed^h�%:���x�z�i���T�CfH ll�vP�KG-���b��r'�ȃH �}�x���(exʖ�ْ�b�ȿ�r�w�^�7�ë�Y�|G�_�i|u?�W���Bhg)j���pG�'�>#�4��%c�:���0�,�o�-D�%�U6~�l�f�DzXm�Jմ� �&��?�uh�/�l��7�{��\�Ò�=��#�t���`ꝬT@�<���=]Z'�2�1w�	(�R'#�U����ހ�s��^jT{3��H�5�Ǚk�<��?ͪ��'k�ڟ��;��ш��(�?w(�](�J��kVیw�5r�WD���]��\���:B���G���k,����G�~7�MG$f�Vr)/P���H2Μ�љ�I��?���Eԡ���]�	��.��QΞ�9'_�r�������Q�r`,t�! �a��T��!}N��գEҲ��j=1"�q����+�m�E~\�aw�MF ��H�߇ ��JJ`�^�9��6o�ҞJ�SQ�9R�tz��#��2��Gþ�]
;;,}32-��%з �W>4���i�Ww#3(p
Ӣo/PJX����>=���7^Q�䈤�$--�etй��5���(i�"�r��.���}�s���;�m���%M�lU
�U�2�|��~d��+g#�z(�v�a��`��	Z4}�.8�`�_4��s�c���H���~�g^%����h��OG�h��Ν�TS4����/���ԓA��I���7��}�e�+���wã��q����ǚ�C���<���:�������+���y}��� �Ch���0�9��J�dܭ�bF-���Oɨ��j6ҙ<,�K�}�$�"�����B�O����Yg�d���Th��o����\���Ad{XbH�3of�s���:�'��P?�ڣ��'��o�&�dt��P�(�(�4�8�$�	�UU0�����]������02�rN�J����-K@���gc���d)�MfA-XY���(�۟׺� �LD�x"�';�I�<�8�[[j�W�:�� <�WRR��CZYv��/&����BL��E�A ��˴[���f���'P�<��]�O���L��x��g8d�]�����c�5�����;�r���u&㹼IC�	����Q,�$��I�|R��<@)�T �~;�9��^���U$�LnA�Y��t�Q<ϔ����P�����D��X��#���7t��!���e����I9I����o�I�W&��� Xg�t�0�#��b�|�𨃵�,�O��f`J�,ZNP�ݔ��_��! ���#,�.X��fB��PS�w"��ߛ�F����$DW˰��n ��}r�<Cp͈�ꐼ�����nW��_�(���!�yQil��\��N�Kk�o=�H��/���	,NI��0f��=��f?��}�����u"�!l˛#�GR���U����h�D�����\�xΖ��0�c�5%&�o7h���(�Ƒ�a�?�c�F$^�#�9��dU%�:dH Sτ�@�N~�YTr�BT�l�;�G�v6 ��#�UÜؗ�ZNӌWڃ+r�3v�f�+�͈����$�H�-�}\ɑ<�<���fV(�N���������kqi_���+�F���+�Ԍ�,�dA�T��f ������6�_A��*9���@��TIT�d�Q�&Ǘ���z=�ph鴑�����䘘kwi���`�e�Ǭ!��q�d��S��[�_AL�̭
��YDiH�C	�,m��n	���Z��5Y>�Ҫ���=���'eq�9�f�W��������各+P��#���R
��D�U�����z�`"k��y��5Xt\j��ƴ�4��Vr�G�j ?�|���m�f��F����Z�v��{��jQ�-<�z�j}Cx�i�Hb� ß��F��"s��9]�_1i�{�3�#�%0r�I�Q�8���������5]�W��������-��\r����)����M��B_�ZG�uA�Ёp�,��m��
����/i����<n�&,�Sp������	e�} 5�5�ҝjp��|�ӯ�(2�`�O3�������x��x$@�g�ߵQqƾ�r��8�7��V�� �3?F1�v�o&�	���ӖL��b��ݽ;2+�z`�y�4�f\��;V}�x�)���<\A�,Ѽ U�q"���Bb���l�(���}$�Y���d&�b�\�H�T[����)ϸ�k���B��gԧ~��z����1�xxS/�';)cD��I�amE��x"?Q9���x>ǹk68�9������s$���3e���65�e.�0�C�!�����Z��Rm�i��q��P�Q�U�z.��:�Eُ�a�d&�98s��s�k�\Dx��ݲ��
��~۵Fۂ�y&���"��_^���=�߸po�x�`�� W?�,��D��iӴ����̓�څ�@!������!��]oN�l�6+[��b�J��?�n�᳡�w��?�H�.y�7E���9��0��N�ɻ��J�i�}]�Gs� 
�ic�^_W��V����+4C���8���F�P�l�ɟ�A-�>He�:��ά�}V�f�$Xoݽ���ȷQL��t�G�\R���r�2�L�r�ځ�#/���e�ɜ(!��x��V�@���|�F����� �
nHʊD�3V�xYh,\}/Q�����>�5�JU	��!ɀ	2n1�w�����q�Y@���^�p����-�A�%Ϊ�.=̠�G�y��*�-�;��b�AEq@�{���PD�,m�'�T��ѥR��|�o]�;�G�RW��6� �0�����o�;��2�,��B��������ˌ+k.�K����2�����l�6��^�Fﻌ���c��% �Ӯ�JQ� �5�����|�׈D����cfuԽ9^��s+rʽK0Uu|g:Zn[l�g�jǷ�M�*9�t�1\�$k�$y�.Q�讴�;ֻ�T*T �x�-'��2a]Q4�qDV��We7��=�i`�������'/2<���}�  ����'����MO����S�w��B��w��I�8��&Dg�-Yen��1F 'Y�L\V�;J��[4�r�Y��8�a���>�O��Z��p�\RA5�3X�h3�Oh8�"LR�y�e1�[���'�5mC�,E��o��b�mq��+9�aH@hS�͡*�):?��/~���(���Bg��@��up�6�x�{��L)��ѥy���Z����A�s��(��2<8��H��[��z�5�xZRN`=���-���o��s�]�M�I'�>���Vh�5
Z9&=Uw�CF��Xą@�h)�����qĒ����]Z��ݠA���M!�ǝ@5�G=��*��rM,�DL	�wq�'�z3����L���U�'�a�0`�*!ʗ��+@|��&,[�O���@�v��7vv�����:���͗n�Nփx�ɤ�)��ʭ�0�d͹:���k�Y�ڷ-�G�N-��,q#{�����,���s�Pڟe)i羜Ev������so$t�"ʁ�E�#�lѺ����]�Bs���ͨ�a�������F�)%�K*(��hC�5Ux��k�+��rU���(�u��KM�?Q�1*}�����M�@Ղ�|���NO�#�j!o�6��y��՜1t�1~-�iw�u�>�o���#T5�{)M�%
���m�-'���!�Vn)��u�i9:�p�TbL �wF��fY��z�$�n�r��א �Z~�A��~aL蠛m�Я����b���J���"w�?r&-1��\���	~}^Oy	�D�a"b�ˬ8�/�S���ĕ��U����NL:J����4�.��� Ϲ�P\���M=�m �z��+6m �T�� #C��* }`���<�����>�ŵi��*$�<7^��JŔ���i)U ��(\�) �8� c��w���V�M�?��T {|ܺ@�8�����>Ȼ�uѺ��I��_E��!��Ζ�w���_���u������� ��~gU��;(wK��� ݰ�~YI𠑹��ͷHw!1�e�\>3R6����_>�#tIʐG�רg�L�/��0RɃ�wC�����HLɳ��� t4�)Ź;��록��ɢ%af\���PxM������X�%�T���x�ޢ�����ɰ�<\썝3����x��'� V��9�F��<�[�I��Vo#����Y$J��h��SN��%��C��O}3G�W�r�}���;�M��=F)ռNgyjy����.��RdrbV[�oqQ&�<d��*h�W'�>ԡ�+��/6�Dd'��_k�
��4(�o��(dg�A�����6�!��2�ko�֭�u�	�iߨ�qL�Y,*M� ��a�F��L�k��:FG���UkjE�b`q�?$V����I�]5a{i 
�CR�AEB#�bE����4���X~��:ы�"�G�O�(Rl<ث�O���
v�*yN9Z��5��u�u��P=�"��o�-�d�9�{��V7	oq��������
��!���yf�~��`N�,K%峪��F��	0��-�$�)\y	���)�;��B���4���K���Y����FD�h	[���{�����S����-���}�����ǖ�
C�#N�M(�U���t��-�莓+��s���切�����G�6DK�o����@�V�%F�}���G�_��6����Y:����$��mOD1�0(�����B7��u�G.sh'�lD��G��3��HL)�CPe�Ȑ-��ܢ�xy����t��<j�q���n7��(��s�%��i�)@9�����k�o3�t�7���{��s�Z%�ls��z&�"X��ꙥ�*l��p����$�(���m��1B'j���,7���Ԑv��Hgb�� 9�|��sHȍwާQB��&O�Х,���;g��B:�@�7�U	i+6ad�����9iG�:���_+}x���C��Z�P�Ŭ�#��J��*:�?i���"�dO�g/�`���LB�9hw�_��B:ׅ'�w ��0W�8.��`:�2d�[��+yYY2������.-^Gl��}�`��$Em՗��@��φ�l�(�\E���p8i`Uآ2�� �!�&�d��5$O_����I�Qf@�<��X�b��L��DN��nC�"Ic�\���1�O��\Q�4(�1?�w�;���6�15h���H����s�7A2���ŏ(���l�4�����]��8U%�k����G[�uZ�rx8��'a��\g�����9M�C|'D�	(���'��j���P8�\&��h�*h�"��ʀ�|��F;&��Jm�j�@���@F�w���OWj���ǀ�Y*�M%TY�����kW�����[���iI�I]�C3t,q*�6��>hy�d���g:$e�� P.q">�a\h��4�> g�@���R��' ݒ;��+�x�����'_P��ӝ��h|H�3kx/>M�8b֑�������t�Gx�I۟�����F=����y���t�+�]�0N�%<�"Nk�/=�׽◮�#^Ȫ�3���="�R�MAC�if.1׎By� ��+h�ɪ�_C���;~$6���҃�����^��P���O�`����F��ۣWNE��#�5"�C�![s�١� )���y��ҳG���-�+�ڤ�IH7>��JD'w,5bn=��P�U�G�4"�zȰ����w)R�-�,֛��g��S�'����M�'��B�W9�˪$9)�3�Ѵ�m�������1|�n�����c���
X$�!"�e�UK���{��md���Ӏ�<�=x������hw�K������e�)}`y�W[�/�cZ��$1Yl�rT^�ֿs��O��NQ��J�2|����7p����8����Y���ȑ�\��=T� �
6�	S�?b}U�#|���&fO=�rY����"
i�z�p�u��		=��	?>ߍ�������FZ��ț��.!�W"u�F��|6۫����W��q@>s�*�%��\�+*�7�B�Ht��C���̷im��Xe*��dy�?01+N֔e�����=P{�N���9j�Y
�����=I���1;���c^�Y W����C���G�S����	a7��%� L�p�t�D�g�@�`7�os�H}�G'��L�%���H��j�]o�=0�Y�GO0-H)���
�.=}Vpҩ��^�)׈:�hM����̊zZё����?���;-r�F֧�68�m�r�:9:�"rB�� i3Z�V
�c�'V@LY� ���1Y[~���	��j���Q,W_��Π�1t=J5�"��n�"  �B����uA�\K*��v���Lk� ���WW�X�g\�B6�{�i�@����4�5,�������@pA^܉e��!k�L��XTN:FՃ�k�)1Z�X��[}"�R�f�&�(Zw|k�_��b���-a���а�E��3"�d�PdE�FE�s�2lP��Bu��Uo�!�6���K��<�w���T4l?��^�6g	����U+�jm�i{TLk���z�����������ZRG��hsw��pd$;�jJ�2��H,��a��Ug�H�qĩ7sm��Ѽ��P>pB*Z�>��p�����0A���$�j�L���~����!���vvp�<Ϋ�DUg���֟�ٺ��f�i[�_hר۫�8��!�陳�>��΀ŏ|-�sG���MwC��'5\����f�&���bH��yx���/���2�m*Hv��Uӧ��q���`��.�=�M��Z��r�ք�юe�ȧ4�޾��v93��2����/��1[5&��	��Sq��䱀��+؊~Җ-C���/��U�VF~�Vq���=ѝ�ڃ%����<�4;v�(��z��QL0���%���䎈�TR[�kw�l^�W��/o��-�y�k��%)X��?O����i�D�c�e#��qT��*��J�r��ɣ�|�;�#��ݓ��K���ֈ��丼t �C�C2�o�A�}�����^��^�b/}�8���NgZ(�l@����2��>@��l�>�^t�^CC'(��Vf�̯d���^G#[�^��!<a�9��%�Qn��*2���&󉻍h��j��O�?���Fo�_���kq��ÔV�w��r�2!L�tL�Z�b��;�}h�7$���L��z}Or1�ξ+)�G0�Qʭ��?1�9P��G�=G�^���?mR�`�0��7��y%�j����%oŸ���.?y?y���Q#[߷t����NצG&E��SPI=�����ǘ<7>�Mڹ�aw����a!�{n�R]����+|���!1�-e��Tue�r�f���#+�ã��َ2���B��Ҡ�h/���:��!���V]�4lz���ߠB_#I��Y�a�vr��'p3��g�?pga���O����lhŭ��D�+�B}��	��)���>*4��K���)Ng/^����(�Y����J{,�X=�K���\�7F�g����R��r��7^�"���C��5��[K7p?���N�j���M��|�zJ������r��E���֐��o�^�2?�%@�"�����J:�gk��
w3����ea*������#U��,��]��Ԋ�E9�~B�f8C�F*C��>�M�����	v@�sa>��z1$Nͣ�l�5>�RO��R2y��O��oUф���-�|x�!��!����l%�MG_<ǀ��M����W�Ƃd���m>�;rR��@*�L˷�H|�;�Ϛ�	;�{�?f�E�꺙��j�X�d�71��)	�pdT�6Q�q�|������]c�t}�٤6HtE,�!'��OГH'�V1�M��g`Ʋ`����G��b܃aKe�6��-?K�%�+�i肦�}��sZ��T��#[�#�f�AG�JO)$"�]鶭՟
Uf��������01���ˋ�j�c�c܎:�.~���*kިT�1����ዙ�:�8��$�ެ(,���(�[ @���:CH����,ĳ'�>��V�&[f�3M�^����<z J�5#04A�"��K�WY9���q�o�Gӄ?�����r�1kF�7f�Q� �kG��q���~��s}�Rү(�Ϥ�$lC�!!~e{v'�[$R�=��j��F�Q#!j2�i�����C��7W��w���9�k��Ο���� �+�t�R�������n��/R�kȶC���|�R4b#ÒE�﷎,J�l��zt^�U���>?����w�G�Ix���y-��0'K���5��>*�e��	���l��'I���� t��8�߿�h�!�|��5�{��'�<������{�� �/�ڵ��kr��0"�<����K��qh���f_����_��k�J�{G��<�T�]�c��y�YsYV�����i�z��Wa�(ƃ��2هU$�ʘ[�v�����Xm�ɔ���v1I���Z�j����B����sL�����X�1S��e�z���2����Qё/\[���A�=�(\�Rg��u���5��i�E+�IP��D5�/+v����5�DS�ǛM�O�@!2�~�)�;(7��p� �����E�����՟��u��­�P�y��~�4}>\��
�K�A���X ��{YC�G�gX�B�8 �L�}j��+�+�@�Gp:M�c)����c��c$<����<=R�������;%孎ö|��К����Ɵ�3Să"�W��A3��/j�\G�Q�7,}��}� I:ﭝ��|�0�1Z��PvL:���ݛA[uE���EGe]��+�WlY2Q	���c[�5��!ઙ��G�lQ�;��z՟�:��z���bn?]qu�WJ,���(�<c0ny���A[�p�:�ӎ��ͷ���_��N�f��Ñ��N�O.�@��
;���~��YO�q+~gs�_�M�l>Z����LK�w��m��4��2(Ǘ�#hQ�zO SfBpD{y��KX�����!������!MYn I�;a����8����>K�w$u��Q%N{;Fy���{�2NԤ��r=y�1��׻>���J&���ޛE��&���<�x*2���V��e��Z]�><B���˖$��ae��;$f�҅N]�Ijo7��P./��ʺ+���Ho����R�ӯ'%��^��#��/�#�xf+���9��ǎ����52�?�x�8~�~&��#���#y/I��b���R�lWm��������ņ@����	>�rc��_�Q���IQ�^���s�;�4�o�~{��eI(��4�5��bY oA�`�h۴�dԉ^t:[�=�����nϙ�`]�da)-��\8�nс��xE03~�`�P��n]F/����,��̲��52#��k�؊��Yi}SwZ]��gR;`����ߟ�2BU�4.%X�ۼ+ŋN<(����XS�sa��/*)��$�/^TM��z+���?�"��N�Ӑ�	�O%��u>�_'iǞ��ךx���?�y�%���
G!��������$�Џ���*���@����~���r-�g��6��,��x�%�x�Iw�=<��z���J �~�)���\���z�(�=_(��qY]�X� N���Ɩ#$g�F%{R��uŕ��%�uW��(#Aufݮ��PR �xW�_K�ˠ^$4jLD�}����YN�?9f	�t��*�'�-��6�� �4ڝ�	���Y������*`�B��=��9�����q��0 ����M�ɫZ~��CXԝ{�]��{�)�f0��o�Ɣ1���!΀ ��L�0?y,�"� �I訮[�����#�fSt� 1��+�ǣl	)W�F���HQN]?��̈́��~`@$�+AX���ͳo�+�����Q�][��x~�ߣ�D�;|0Jv��9[�<�$	L���HF��k�l��u���<z�A�p��p؄�V�����i�ͱ�lv���/�Z��{���X�:Y������w��Z��\qT��1I�g�E(�i��@�\�`�B�0���{QT�TҜtD�T�!�1���C3ӥJP ��,��4j~��P�s�b	��k��	��>�� MM��k�{�����#Un����A,�`r2��^ܓNT�B�R����lq��U,�2aG��.�$�Ii�>��wV7�s4��b��-�C���*���p��K ��hڠ%`�����^��=�8�	�u%
�d�M�،����Z&r�#0ܩ8Au�YRjc�]z����G����%;=�հ�,��h�?�"K ���E���Q�Q��D�t3F1�}B! �W���v���y2z���x��˲���DR.�nu�����w��v��ސ�;ۊ�nt�Hh�τ�w���,��t��N��r���B���)"�l�u�1�#Ng���� E�:��Z�`����;��R�P�~��{��
��Lą$a���qB��P�#0�V�08�bf�Ai��{!�p ���g�P:���6?�,�|N�v�j��C�Gϕ���q.�G�y*٘�:�6�&L�()��k���>���`Zh�����-FY��lc׊�A3��s�{OG���õ����iB�.�c��D
���KMgf7-�k����"�&�1R�ӧAKc����k�o����� IE~�g����E7�36�t�i��Sp��ټ�&A�6�G ����]�ɱ��{~�HoY���}��l��N��F�H����j���H*�ϖ��Y rLf%b*P��|��GC�1� cË��_gIc������j�i+��7��r=,���}fb�#�R��P�6M�Z�<ߵmݤ?݄�n����6\r���M�/Nfnőa��5�o5Jk�SH�Z�:V���Ȓ�[[�O�5�]��=<��h,d
�6H�Ejb���I=��4|�i�������u�������$���q�R݊V�0�Nh��}0�/mA�E��S �C��� 	@k0���<�U�wG�gs�q�w)c�7@'y�����P�'�2O� ���}C[�P�c�w'��>�ѿ��	�p�S�և$���Z�3��Z�J3��G.�h��LUp���ʆZ-	$�2j���4�&n�H�C�<�J���H�S��+����V3a��Ø��O�b�j��|\	8Ax�6��\� #I5֢_樲k��i8���;}uQ7ƨ�T��JrolQ[-�.�$wm�y��Zΰ��<K)Dmx��wͱ/L�E#�f* �[>7%yq�Z\��2���: q]�t�=+E�����Kx�9B/<�E�f���/�:�T%W�	�-�ɝ����vݗ�A@�Fcd�&�E���w�S�~����+V� ��&�� �2w�i�e�,��l�w�} �7��θ��xd�Dn�;<]�тf���y􃱷�b�P4��q�+�>�Ad�S�l�@��OVWwB�p?��ߝ��c�dn]�ܘ���DQ�6<]�U^re���F�A��&�#.��B�d:W��G}=�]5k��D���+�#��NzR�P�V[i��}4���es����6�i0!s��o�]%q�# �j@~ۺ�I�i�OA�	�`aӶ�ʡFm�����[�JI�	H
�D�U7$�2�C���� A6�Q�p ��P�z�X*�[��>aFp�%�<��lf�%kX"��۷s��7a|d�	�̏?<�}�Y#t%���p櫼��*ymfCNe�n�1�5�bM�oT�D��]���6�j�A�e0N��֝K�3�㻁�u4���F>T��U��î�%�r����\�m�Q�KZ����$��M[��p��� �����9�hzi���<����	�=��=p�:='�(���ɇ�
h +"�?�S4BP�AN-���9������W�F�}����?�W&4�b}DY嫘Y�N�%T�J�_FO!i�K�O�a�wv��j���e����qy�Q�Hp�}x�kq���9R�/�&�I�Ch\����_�!3�T���@e�w�g�G�,�������%�B�h=>�8A�!�׵V	����i}d�iOX]c�k���T]�Lt��Q��5�����8"�T�y�c�@HF���6�{Yo�;t��߃�(��)���&e���G����h=r� ���`�wv���!�;��'V�E>��K!e�~�R�S�D4���N!fJ
	G�sɗ��f o15"��`q�qv\L���y}��}�q�i�C�����0o"��r��� �'�fo���(��s:1׹��4=��V�ly��XK+tš�`���1���o��������	�J���H��V�ӓv���hE�}���ʱ�t�t� �V=���N_By�1����=�U�E�+��o���������:�50�xK�}�2���ݎ�Y�]2q��Y�����v�L&Ƌ���˹-�����f�) L\�x�y:x��ZU�55et���(��ocGj�݆���Ϊ�	iه�p�(�LѹF�K첵ֺ�бn |7<����l4�8U�r�M�"����U6Hca��>W�bĬOnRs�� �YN�|8�-�S�M���L
�����?����8R���UN��ɱ�@G;����|c�є��*'P�z����&�X�*ۊkf�p���>�:�������Zz{���f�66VW`�ɡ�X�R���j���{O�y�a�;:bH*Wqs,�u�������K�t�/+�tC����[o!�Û	_��^K�aMH]��G |j,����㏚��?�s�G����yIj$?` �2_j��d��G�S��"z�,$�B_�������8��<�cTx%0s"��S�j~�Q�����\R�M�l��<M�'MAE�VU��Sb��=�C=e|h�})�[��ֲ�J�1<ɫ���t���q��$��T��,6�i|R�fTe�N�Zad����1�о����J��*������z�^�=%�?Lèm�a_���W\�3���c�PA�#@:�F#�؄�2@ܗ�'�喷�6ݹ�����x���x�,�<�0pr�Y��U�%L��DΩ�aUӉ��Xy"J9��l�^>�L1�瞡O�#Vp��V�x�P`(�w!AWh��y��Xy;|�q��U)��*RRl������P�P��H�r`����xP�##��i�Sq��"�L1J�D}����f+S��朻�&0t͚ ��1˘��j�=�<�� �:�Bkr&B�t����=5C:�.4*H����t�~��-+��v�QjU䴣����"��4خys֓Ѽ\T�Z|JK!�f.?��� �X��2�Du���iEl����ՙn�3hC��Ql��������;i&D���v���{,*����Y�G2�WS�o���;�󗽩S�*��9a��J$p�{1�:I�̣�l#�*�<kk[#��E�f�_��
1�@f��%�:" �����*WR-�sR�;�"�2L%AG%淿�+����[^���ay��ѷ�,�"�x�u��\"��~.}��p��I���P��.(�S��r��S�҆��!���>/�L%��_ݻ+z|
������R"M�I��A9u�����L �n�ڶRp5�7�Y�ܷ<��r5�pSf�\@�^�2�J���j�Mp����у���z
��VFPF4����p7��۾َ+e9-!��gY�JUQ�j�ɲ�(<�N6�e#�iⰘr���2�v;��y4�zk�Jҧ��x�㧓��[gRʘ�ޥ|�� Z����.1{����(k��mR���@:��0t�$�(0����L�bOz�Y�0x�af`���Λ2��p���Q%�I�9��vl�i��Jc�>f	�0d��ì)�j�?�S	sB����^�k5�2��������Cg��\G)Ɵ#�BA����;"�v�%ln�z琦��ӎ	3�1ʊ�M��������MC���>���������[�pv(�.���(^�>�����<�#O[�z�Zf�<�y��z|��J��9|]C���^y�s���N����{��T��Y��H\�B֊�����e��DgX'2�3�c��gNx��T�"��Hi�#�hwTl�e�0�Х�-�``��@ �U7tY|n�2'Rg��"w�lu���#��b�>��\��EX%���6�:����n
�%���Rf"������*�<Ѥ��C���1�c]gb��g�G�� Er/����鏂*��k>�"9���u�a�ݐ��?|�z!��{�����So��1_K+Q��A�����n��wzz����4�U��<0��w������l(v �|M6+�������ڒ��ʬ�B���R�j�}|��a���2�'�ڠ����}#��wU��
��
&t��(�.�-�^�0��ED�|}1�Wh���|��u��.X�b���0�و���u6�R.�"��ߤ�ZlY�347P<3-X\��� ���&�ϭ�;��(ц��5!$J���
����"�o���(�Z��@�4�Ƭ�8�)d��\�����I��ۻu�>}n/ �Ǣi�����q^]K�ì5���+����[��9MRB��~b�,��N��GuR�Z�aaՓ%�L�#���aq�ьDsGǑN����ω0��}�j,����K�񲝅���a� �f,\���̀O��_g�-cPfu�܃���yx����T�3�k��6�{^����0���Q�\]g@I<)/�����s>��zTTQG%"�W�����畫v�.��M�-u�}I��_k!���O�#�f��7�����&�[�T���(��3�#���W��Ȃ��n�t��?$�[��O��b����K'�؟p��+�و��W��ߎ7R�:c�e�{��Ml�?KG���;o;�O�0�B��Q&�vF��}�}�� Q���콛�NPc`,��tU�^���	6��l\�F��hc���8�=��/��]jbƣ���[��JǤ��yn�|7��G��p��K����C�J�i\m���&4��6����b����p��B=�����g��#�o���4�o3M�U&!0��wk���E�5Oҗ����V#�^�;v�i-��DV�fbe��8A�R��%Ī�5����}�V��f�g�Ifp�ڟk���ڣ���V��:la�����D����M�J�8��g�ЫǢ�9j��;���;�8�����酑 j<���糯7)�B�#j����sU���^�Åݩ���߾����ʤQ��N�_�#�!���D}/t�H�`g���1�<�����RC:v��r@%#�e��}ȣn��;��d'*!^{���*�vUx�	����K$&!���}��[%N�$e��y�_
�4���`q�l�7+�n�>��ޙU�}~����5uP���,��:�jꨵ�w�>D�i_�ً}:7���c*�U�xUU��WN�2H�"q����$��g[6�
��:���6���!��������Z�t����҈ErZ)x�]k�}ؖynG�u!Xl��h�K��?tx���\ӝ/���yYYy�������D�BgCzd��S�' ɵ�źgږ�$`����s� 6�?���fBr�>�*���\����F�"�x�'`�冃�W�b�v�
�l�������ÒP\��b�Xkj<=m����^�CD�� �~�]�)?�#����!q6D�|m�7;���7� ��».M��2���3Wθ��d���UR��=�4��L!�PúaG�f�%f�@������$��:$��A]�Qj/�B"w�W��TT{;73�B���f��凭��+�7I5<Z��#�K�7��J�8��LS���	R��Ȩ[���7PӢ'01Z8�׆�����ɱ��2����)r���x�,�y+9�#m�|��@EU�~(��U3�<\�
q]���%]�d~���P}���Į�F��-���i�-��lJ�r�����"�mKG~�'f#�	O�Q|��ۭrI`K�=��ۄ�^�ﾨ^�E�z�6D�:_�P�;����J���]�sK�R�:yجnH�Wۧo����qy�!Tw���F�)��J�5Zj��=:����yU�A7"��s؝F(��Nvz�YmF��8���1q�h>��
=˙��g�2�T\�d@��K���ȁ8#�Ş􅛅ӼǸ�gz�3��C���t����N�g�z-
��Npe��C�#��['*W&�@�_���q'xi6�.UG�k�:D	1(��f�@��[��@VA��λ�~c���ͽ���4��\OW�@���O����4̭���᠚!��FR|x3@\&C��1Z7�S�Τ�.��I���D�م;�2�8�深m+������k�Kw��ւh�{�r5����Y�{@�|�Ni����Ah�u�,ey���^�$�=KF��j�wyr���r'3?�Δ���6h�����d�d�Guc=ei�%��3��m\h�,Ls�S�Z�]P]?廌�_O�0q� ,1^52�V~��ݜZ�%-������<"��Hes�]� ���8��0�J��Gki�������t�qa��0{8�
��v�v�k�ī#�NC2��Y ��Z��:+��T�Cy�F����r��0��:���F�_⒭�֓�m�,h�r�;�ЫDg�^�(y	���Oآ?ޫ�+�o\��-�)��$~#������X�r�i\��Wi1o�$p� /��>�:(p�������M'�5�]*­qMS��vgX�ں���L^�ᴠ��������_��'���T,��x_�z�kQb=7I����IE���C�-�PP���<�Q��8ŗN�(d�aQ*"�'��j0�II�֫�ۖR�q�����h�p��#5l7@,�ڬ��uFPX�-G�-{�Y&�:�:�n��Vgz�3�x��)O���m���w���x��C��~���{4���1����Y]� �����f-�����5	9�f&L�k��� 2*���]��6��d�×V�6P�_2 4��7�5I��2ܕQ,3���m���я�[P5l��9�j۳#�Xp���&waeF�"!����^�LO�Y!&��6�
�>��?��M���@�˛�z2~����pE@�g �e�Y�	����]͸c'���|b)kCb3dC��e�l�qZX܅ߍ�?��Z�F����5�O%��S�tl��_#'Yx<�ޅ��?6\�>܊���C�����h�{ �	2#7���݅�&O������ap�A�
���?^��=�v�z	��X�g@?�N�Try�]�%�-!r����t�w-�X��j*�������FnG{�Cs�L)ZK;��s�������d�S��1شt�n� &�@���qa���a��FL�àu��o��SΪ��vo��/k71i"L
�U�8J�$Åjv���ze�dn"�7U��]a��Q[�eԌ�
ұv�zw�>+��)LjbpO$��W5v]Z�^��96͚V��d���)��r����h]�U���g7�.�Փtc<�=��u="����ď(kB���@�A
ش����kJ��&a&y�^�s������^��^��2v���§aC��n-��ݲ�}���//-�}$&��ʼC�r� �ʎ����Y�F�_C�ˁ�(��l�>"�}��D��_�P)i�d8�OȈ@mx`"��Ʊ���"�������s-߃���W$*�dg0B֖6V����%�z��OB��i1��VJ#�P��Zg��܋��FѨs��~�;[�}`����L����&/�f!�[��� �[�Ӱ�fɶG�q#����Ƿ�(rM�&�m�/�����~�Zu��
-�T^�B�:)4߿���'������A|~�bT�F?k���������oE�NR�ܗ��jB.3��K x���K�#O�'��.���h�T��f�	�&�^��MW�PHZ��e�0{���5x�4�b�B0���h�2�D���4��`��y��\m�b��q{z[T�������1)���J��R��A�����,I���`��]ƗA8���Ev�D%E�(���rꀣ',��S�G,l��5�i+�x�����B�ܿ�*���8MW�g��XQ�\�3��>5ʥ+���	H9�����r.<��Q&�SS2P�q��%؁r�L�D�\@����h�T��ЛH_{a�;UUdI%����+V:�V�gU��{OПB��2������tץs��v䦬��B�^�g�x��Y�R�梔��J����BlȊ��c�����Â��E�s�O�\v����4x 0���'�������mn�Q�kpA�n(m�7�zT�A�6�ۆ9>�S��� �(6�`�K��JBa\s��؍om^�����P�ۭ���B���e�t�Y����U�B�|��#ky�HS#���Q4�M\���"��+��O)�.��Fn� +���L�t'��K��eat�&`]^{'�`��Ͷ!�M}��d��O#��*T��'ί1�����/���D�7��Ɣ&<�6^��/�����Fcl�J:/:�J�R :�k���q�{����X"4�d?�H����(-���+aG� C4B��]y[��޻�n��w����K�'�|�/�S�eW�	����&-A�y'+T�-^?�rj����c����`�!ai�Gս��K�{����CPdA�������Z��O�y�j���l���ִ%�Ed'������2z�\��y�-�{�Lڕv�3V>&Z4�NE���)�賥������kײ�	�LZ��x��Fb�i���q-���Ah$�=!�B��\��cbd��V͎�GZ[�|��T�K�}Y$!���ж�U~6��4��b+�|�~�T'�/�edL��'9(��;[�5�����(�c�XB��jz]�O��Q��*�?-��7O���:~G/-Zݭ���iVo��<7��Z49���Z����7����hP�WL;
����1�N�p@}��/	1:��\�-h�����ܤC���B��C�D`��I��Zy+`�
�:k��T�h�炴}> $��C��)/(!hš)���L���*%���Cl�A������'B��	8�Rm(M,�f�<wZ\i�ȂjPh�=�ʌ��C� ���B/q�Y��z��axU"6�b��*���A��^;Һ/t��CM�Z��	����>@B�XӠ�|�CO�1&P�q�l���0/�'2��BC&e�J����ا�%}7ӆ���y����dU�\��������h�}�x���7X�1��k琯`�]�Y)��X����������劸��k�:���]��$Nu��A��[��?gw���ߩ���kX��Pj��j'O8z��C��q�b#�6��,���bY�e��!/�^5̞b/�qc�!�ib�3�.>̤`���j�j�?�p����n�rr��ceV��b ��:����WO(t�6��V���y�B�V6���fVF0�T��Ү����1g�`���1��B@w}5Sgir۰3�hE$��2���,\�8���~���ɱ�H�قpHp����G?�-ڗ��k4����i@��Z�Jl�cF�r�eʔ��a�xk2�/<�� ���K�xrւؙ�Xh��-��`���Ps&13����¥%����nE� ��_��]��޽����G�7�ʦ.��/M\�� �\K�����ȇ�14��x�$���#�k|����9���g:�/0�I�Cq��8}ߥx�����;��1~��"7>���߾���)m�hѲ��Va|�>�5R�f�F��
��N��o���H&�zI���ص���WRo}��Ì���.��ZK�U=�t�	��EĄU��{Hj�q��'��+�'JRjI�9R��]:�t짔W���Km�p��lNPL_�GlH�Y�踕���e#)�e���6�G�K�<�@��n���m�#�=�t������ �����S�-����E �O�y�%�r�k$m��wW3��Q=:�����Ee/7��Y�SI�UG�0�4�c���"Y�"o硄�0X� �]��\(����� ��Z���H9�C�b��߱�"OH��!�2?�d�TZ�1�ټT�"�/څ�^�]��?�ؤD�y�}�w7+Iև7J��䇋�bз��\�_2sN�,��a�.�uv��:1n�yb:�T׃K�.��*ץs�H8l 9�y":&�����l��7�C��D<�5�m�!s[4p،�F��Z� �ږ��heW�jҁOG� r��ѽ`���󳛯g*ru�TQ�Z�L!�͐���b<?��Y�:D̆PIZ�4限�C�3�����E��5	|�Ѽ�f!M�X[��ۜ*h�����l�"�x�G�:l~!ބ^_e
c�I�:��E؁�X\������'{��%�(ļ,zzCg4^n�^̗��1�<e�n�T?�|�bW�:�(Ε�X�j���#�h<[>L��.>�?[@�򅂹8���Ŵ�d�Gm�[�	�5�' ���]�y�W�[�����g�b���s��s��| �����Ā�:�v�^��[l�����2�)��K��}e\���c�Ė=�:��eW[P��gO�{J�&c�)��}Mvl,�� �Z�4*�%�������P\L.�mQ�>I���U��A�����AS�����$"[,7oLl�-���s���8p��;m(���c�L�5�Fx�٨5�8_���5�ѡ+;�w��J7��b
�RzE�o���a.s(AY��=-RX�q͸ȫ�q�${�I��m�z�-��	��4,D)�!>��U,x��Q5���4��F$'x��]�:@�h!��£/�r�m����v��}��Ҷ0ۛ�$;�����-�h���r�z�LM�P�f[*��=��Pq
.�!O���+�P3��o���p��m�Y�@��E��>OW��K���OӐ�������"��m�]�nz�K�IFW�O�R^������l���.�4�� ������9pH�GW �R�Ae9��� Q/Iz��+Y�@LϮ̄���F�'�[U�z�;�̬u�<$S�nЛ�	0P���I��L+
�AZziL��q��|`�+AY�� �H��c�^~�@��f4��NP�����"l������]�K{��lι#P��B0'*|�V���q����R���[Ɍ����	�<�hhG����(�XI^�5�N`3dŒqT-�^���(fP��M���y`�w��ښ���FU��Ǘ������=�s�Nƌj�;�s2v/	i�^b�n���B�� ��ݹ�1�b'�u�Kg���ә��]��ѥ�b�M�_�y��о%�7�g�U���H���\>��p�'��� |��r�	l��v�Q�vň��ׁ�GΠ�`�R5Rɘ44�d���sBEΧϤ�N��`ˎ��h9
\Z�*���ե\�C�ڣv����5�-�WMYeLR�LV���{!�9H�%k���Z�i|��iN�9��m�r��o��'�L�J�OqA��������`tGZ��UH�HYm���.�+2$���G�}���.�p�IaGǑݳ������ǿ�<j�/[�Q���.�*;�B[�s�����!�g��f�5O�U@l�$�9`�
�#T�D/v�{���x���.YP�����E�@�9�:M����5>]�vx�����:��L޹1OޝiuZ���3�6�vj>PK��F�����Z�x��BoŁL�S�I9�/:�I8)�03�v�1��_�_�5x�/�<yr��ه�)�«w�x��tzL�V�5�M�tb_[����	ci�
cZ�t����<(1bp#�O����� <Z����'�3���C�E�L���4�{v�{ع�۩���@_$@��y`�+���ح����\�?�F�J�'�%���[?yOF�ƊQH)?:��]@����a�B1��j
j�o�������"5}a+��{�����a����\C�!^��,���$yy�J� +O�Sa���z���FeM�d��G�d��;�yh�w#(?Dc��P8@��E� �jx\�<�v�r�;�����U;t���ݳ=�[o�KCy�1��O�����V�8d�&4��!}/����*�P\�G������7�ښG������c��8�gIY|��'TO�I�Ǣ��O�Z
M��S�m���6�����A�Kn׍���,@�x ��i̋4�e��f��o��:h zX?2:��=Om�NN�'���=�n���3ͮ�W��mf��ז����qW�N�7U�0�rSD��2YR�s�-�Cxfm�<����)-�o�~�z�<PHŷ5����L��Md<� =鞤>�2ӻ�ڗ5.�����jL}w�A'�F�T�?�S(|;z4�ǒ��-�
�S�*^U�RgF�V0�:��~�1N�X�,�i^��I�}wh:M�i9�[	���u�=��r���'�%��s�g��6�����E�$�Q�W�ޥ~S�[C���C/�
��uXQ��M�&����R[�z����H�d��N[>�f6f.�x�6�)�\_(p'�^�
h�Ô�x_�X՗�x��޻�y�}�o��2E$��XLK�btT���7��b͠�T��	�+��D��㟺�	�?i)��
_���Q�5�,1T�/1�#�B#�#��XƋKi�(�hva��9�R���8\��
���E�Y���'�\� �ޡ�����`5�j�B�K��3�.��ߎ�js��p�`Pv� 7�$D�����N���8��n�e �l��{���V$��AQ��)/U|�T��^c�R��>���;��������Zf��,ޖ��)B1mP����˟*=J�v�v4�Jr?��n^�{�<�h���΃!�W&$����M�tjQ�+\��d���\��VT���a�9z����-�?l@z��U���+Pʼ��:82������9��� ��Lm�o	�������y=�������E�I��p�.2h�+R���\nY���Ua�'��9ȏ���+��BOD!	~wT�l��<Q^b�v�#�����/;;q4�gr}��a�Ƀllw&"��;?��}���#!�1���5�ˡä����O�	gN6܋0���%�O��}B$���JF��th�&]/T����\�=�F��9����X��3�Ęv�z�
���ؔKg�U�?��.��� g
��놄	W>!˝�@�L��5��b�h�z��B�'����>�A>�� �j�b8}7�d3����6��.<���)i%M�܎�U.�`�o~�ٶ���l��1��o=wG��K���#�'EЛ��X�����I��y_�y�^*e�)���<6i�:�C�UZi-�?���Z#2 L>�[~#?N�%���kB+�3|H�}4�06y=R�pk��2օ�z	�T�QS�d�|=�´tԮ����R[�����F!(P��~#���w�1�.+�4G"�m�^RH�D����W��ҹ� ��*�P?��I)�����A@�Ʊ�7f��m����1�t{goGJ3Y�S���T6�\7y��Lފ��a~z%U	Q��H�*���fp����6��i�*Pւ����{L��b�RJ�c'29��͵5]'M���`�Hhw���%�AZr��Y���̲�@�"�i-���,��;pg�\�efF{�e09X4�#�m�]k�Na���g�Z����tJ�/�Kiʚ'_��}���n&���&>�i��Wbf��?�B�'�Bxt,~!�B��Hc<��x~Ѽ=w�^��[�ܿ��fx�K�/��JReXp��`"xMN��Rt�+
�x�N�C��+;�@�ja�=��`T���+����ɱ��^N���e����hnC9]q��Z�XL��:M	z�Q���jVvȁ�N����|`3IĈH�hqH ��hhX�'Bl���V�C#�$��h���C�o+J	j�U���Q1`
�-V͠�a][<���(ӓS�+Y��l�0�P�p�?�9ʰ���U���8Os�R~1���0�D���.ݪ���R�!��T�]���\6Rsb��A���13N>>�u�wx/��K���)�.�'Q��	b _ޅ��,��Pөv�Ō�Am�3�����r(NS�p
�����U6�=��=��a���h�!ZE��� ���~g'F��=l�_~�m��7j>�p�����ܝ|t�Qa\ڌuף8:܂�&I�M�|,+�0=�]�������YD�Ĳ�*��<���{��<��Q�S�b���z��3V��4n���t�1"(�����6�wv��H���O�<y�e9�Or��v��D�f%����{pj�Z�Hxq��H�E���H���!B-�38��0�$���o���d��԰��}���եl��Қ���n��@4Q򷕽�%ME��=��C"���O7�nd��eCG��f�4݆��^�`�)�p�)v��3��C*��y9�b�8y%�ڌ��V ������=>�[��K�A{2K6�z��F�M����_E6Bp+a	q5�rד��������T�t��f����{a�5�����)�U�R	�T��-���"k�y4�3��L�tV�zu���F���C3�%\iYؑ��U�>/o�-�mj5G�P3�~�Or{��6�B�"g1�[Kģ��@P��RN�r�&9�&�����#���5�:1�������ba�ߕ�-6��6~L@u�X��������W�2�8.�3��m��I�C�Yu�g����0�n���T�*�+E�����k
��0�lc\9�q���Q9�K���;'�,
W��nѴ�\A#��T�$E��lK�	���Y/��Ӹ�h.�p�r0N|}��Joy(yKd���Ɣ�ŷ�wfX��hN�v��̨F$�eX�e��ø�_n�2�Z�i�7��@�.z�	�[����|�U*�B���1���?�z{�����DA.X*�kN�~��<�9P�2J��`�X�w(A#��#+���'�v'�p#]!�ER��� :!��%Uf�V�*N����H�8"�|X�4bj*�Zx́_p�͑�gO9��\n�R���9��K}�SKᵬ_'|���@;
�w�p��ֽe�n��I#r�I�xD�5wF�/q9gh3j���� �\N�9!�1=^�����s���]�L���0<w/�%�ͮ�k � T��zE�� }Џ'w�TY�{��{)C�BJ�qUy�������5��V�,�_Ȓ4�4Z
3_�}E�'p%R>��v�t���%��-��U[M�_��9�͓A*��$˛��rŭ-�b�f�M�>�i�̕#L.r���,?@�8�#?��M�D�w���;h�I�G>(�&����!�ӛ�
E�t�C�nW#�@����'�S6ySH��f��c�s�ۺ
� d� ����������wM��}���ٌZO�oF�:����� �2����U��[�a�JRȜ���;j�Wu���m��`S|���0&��e%G�^�q��=��%���F���Kpd��d�iǯr�s;-���N[�'Ρ���dg���O:�����;�Vg7�OPIF��A�0o�O���AD��XM��;��-�3��yZ��D�D����;���J�u����d4p��s��]]�������`B�N��w1��������>ٍ:f���1�R��ʭ��E�H�0�y�X�'0[�cԷ7�U:�=s�����#G��¹!��L��@v��v�!�����z���Y���7�Y�?��!�*�����r*-2���>tE�N_�%GP?Hdv	���E���]�>�Y��?�܄m������s��	��H�I���[o+�K6#s7ŝ��z �r���'�#��,�����_-h"˭��2Q�!N�%�T�e=r*��U���wc��'�n��s�}�0R��DՅ���P�d�5�+�G­d�N�ώ	�@�6�I��O
�k��q���2{:�8�#=*�T�9X\�+�$%��J��V!��p�筣oZُ�����ľI��V4�-Q��Z��x�o ߟN� �5���Q���|���9iևm|���e�������>��.!2�}`qﴯp�(�[pl�����F\*G�	��]�2�U4"�ݫ.�^������l�*<� �>���1+ a�/<��g1�Req״�9�=�=��,�P&�ʓd�@s�AN��R���E�"!w[o����1�'h��w:��t�M�[D�������o.f;Խ�1��vB��UF跌}��5�5�E!�h|���I��e�"��$�v���t��5�́Y�~��o���Y'�i�=�'��z�"pjKĚ.���Q�HsA	fʂ���
��/���]�S#�.����n-z�! Y����͘1�Y�%A.�z������0'��,��q���v���H(�k������! ����<����0�E�n�Vp�V��91�㔰ѳ��A�Ct�9���=Gb��w�<��������%�w �X�����Xg�?��x҅{���S��Cؠ��+�v�d?��!����nƌCҪ�*���E�����L��
������L��̇,�& 1Gf�D0���=��`s�G1�e�G/G���tYk�	�1e��\�숭���@�AŲ��XF�?΅&�W�"�8��]K�S�W'$���g�Y�*�$��d��?���Ok�o�^�i������^&���a�y7�ru���0%�Rr���uډk�f�r��W
|����K
�p̫D�����8�e���G�����Яkj+�xS0�Nf'�J�E��ŗ#����AU[���0p9�
�p|��Ϥ����6�!
R�?7�$~���#=�w��Z���9r�b���W���9wÙwNo�a� �S�����܃��MB����L��s���=�k���4�tT���@��RT�X]�[Od4g��	���|�`1%�~M��<:^�$6��dTw�~�ع�Wq9��S���,!�q�� J��03��rE���S/]�g3�M �e�3��1�ݧqh}b)�=p�JC����M���R@��dĔKC�P�b.X/q>y��i�@�t��f~�!��+D:K���l�����m��>�U%[�w8���U�Z��]z�i8Z��R_:m��Ue
@�����h}j����!�j莤b�^1�z
1�-=�{y� �/��EԦ�G)HN!�f��ܪӧ'X�{�ڱ\���u+}���}��6A�FR��h��=-���Oʞ����~��2ΥF=l$p~d������l��_j�Q	�;dG���a�3ن�X�
 �яD8���`9 b�P�$� ��2Q�?e�7���Ak��H��r�?Z���H��~!qwh!uKU$y��)��G�@ƾλ�*s���-Pq[SI��W�yn�Ep=4�/WR k�<r(v���<bS�h�(Q�}^�:��Q���p(ҡD����<�-��R�|�6W�B��8+8Ҳ�H/�q�
>��]90S���pŵ�Mx��L�z[�Cٿx���UfE�<���~<�U�%�ϓ���=NA�[�S�qH�D�7�t@��#I~��i�߫K0BR��n�b���1�����x�tk���^��*U��s^:�%lQy("��
~K�[��z�@*��3~�-��޲jɿhf�Jk:f�}�ꨫ�����M�w+K&�g��V�I���Ҷ�"t��;)�Ա�w(o���F�6rű	Q37GM�J��Q+8�U��F�\*#vr�������z��]�7�c��<�2F]���w&�.���$�����Y�C�~��{���	�5��]ITWXfm��g��ݘRmN\���þvFr̖�������%��)s�,����H�<�a4����'E�̂@��=o��̐i�>S�u�&KL�O܊S��{C'y;`P��]/�f�w:}���è"��tj���a0I��Z�Kv/;�Х/�)�{�O���O�z!�R���9���lM�P�KS�\�OP
"Y`�рi�))#]���Nm;|ԉ�d����}ocB��Ĝ�Yּ���Xȃ;@zWŬ����N�I�z��z%5����z��9/r�5�O t�cbZ02W>M|�[���d/�����zG7U�-Fb��15�~+�L�(σ��`e����%PIJ�^�����!p�
�`p���yU�l:�\��U%Sa�K�r/��d	��[7P��
���M]�zg�	�S(���5���d��nb��z�u�2�S����0dx���xk�I�au�O��/L�G��"�����BI��9�:�y�f{Ƣ�M�²;��"�P�ZO+yr�9�s��h�Ň\H(�z�&��"�o���;zo�r����h@^)�٘9�I��+#���`"C�����J�B3�i�(.s�� �+c���?[k�v(�Rj�����ds]%������*�q�G+V߻�L���s47�`X@�"l*��w(�2�j��M�@Wa���Q�k{��~��*�%��9������xNQ�	D�����;��|���'x�oXwR��ԁcq�*�U^��

p�O5�"SX�/-�2�3�p�/�j_��Y��QL��P�8�(��ƈيU�4�HR�6��
�$�2��1�c�p�:��2�*�.a�(w ��匑]
�9�����;��a��i!<	>�HMG8��z�g���-e	���t��
A��^a��#R���xaW���<�Ϝ2��+�i�־"H�ƿ���8̍m[��آh���hۑ2,f/� �^�-	y3fs�7VH��f412E�'�{%���,��ž��iVTC��~[i�?+�H��v��t�{W�I u�JI�Лљ@��֞�ќ�k��jOR?��.�gIYyj�ЭO�a��B����q:O�@�G�_��z���?�ju���6P���s�QǊ��8L ��.��i�>?�!:jV���?Y�l���I���d�"�r#�(��?DmI[���@�ώ�M*� �>�kU�W��5���/:M�e$e�׋�{�RQ��I�b����s4[f��N)�*��j؍�T��*xJoʃ���2�*$�"*�=�����d��4ubw,V#�5���b<�q@KbU=ڵz>�����,���v������U����/z9���2,��NW��_���7�z�+yC�[EZ0���|�Ƕ,������)���<ml�d���3�{�ș�c����sj<Y=w ��K��В~�&+�:�]�R|N����zzԨ�������~��a��Mྛ4��;~P-��w
<7A#rJË����"�4!�Hs�莁�X%�+�<�������-�O�!�R�.�oyQ��5.�������=K����fT��6|�C��>�2K��d�y^r��]�S��V�˽�c�xة����CC�ߡ�|�6��<dkܺ�\ƃC�b��?��I���p�럛���2�S�R�f{����շ`�j�"S�dt��E��~�v"�:wy��~�xٷd�M�o���`[��䄲]��l73���4/�)d�tZ��f)Jpǌ�	��[�>ts�1�{��b����U�A�6�\I������B>��W�-�؜1�ү��ػ84�xF�,dE�%ލ/�ߨ���2�'v��:i��[�����p>f�;/��-�Iv���
�����X���c�f��(7�v��W����1�T�K�.�&�]��*�h[Q���L���9��j�����E�kk;	��><�lb�ݨ8��#w���XB�~�nL�Kvgk��59�s\�S	X�s�ޢ�F�1���obk�\��L>8��S��y3�9���:k�Nj��sA�p&̳́Q�$Q>89Hkp�kp�V:Bd��ݵv��F�e���E?�)�o��%�S�<�slV��,��J���^ܫn�K����pp�3Wm�ʙN2+d�GcsǢT�ɮ�-U2q��k�]��X�E{�&a�:�1�ۈUp�Óo:��O��F�����e��)&�DdXŐ�����ﾹ�t�@W
��t'9z��ڞ�ݲT%��N[�YǩUK��0j�q�{���]c�E�'[qB�x�<�5�,v���];��t�U�����$��S�ͯLl&��EZ�xYĀ���$�:���{����������k|LtA��L�8�'�#���}��C/�Գ�޳��j���$H���v�a�A�8�k뵧�Y2������0���0y=sbC�%��bA��AnW���e�Ċ���4��3:�q�:�O��)L��{��$�����bL���E�����\�C<�@�[��8̟ѵ�z��X��c�{ۢ?�Fi8��~s4�&c�n�I�����ߝm��%���%�P�b\Z�2�B[��Ͻ�ej�Χ����~�(���0��R�!\^�O]Xm
����<rp-`�ZG���Z���}x1|����ݙ��m���8W�J���>�=���w���!�}F��j1�-��Z��K�fKIz#�6Hp��&��]!9ع���~o��|a�A.��"�L)Ď��%2���y�ևN�.�P�|YL�#�)���0ɨM%$���Y$p��Tv0��?
Ͼ�5,����<��%֍��X �*G��na��l�Z�C�k6��;7�l�n�m�(�C�������h�:��{�¸k%#���a�f�^5��r�`6O��<�s���N���x��i�[^��n�r�آ����к/ D�K*�o�b�zB�P����"#~��Q�l�$�<O$�yAeϵ�+20V˖D!41	��z�]�8�=�M���'��&&q0�����.����<7��r�F���d��`��D�8kX�wd�tڞ�f��O��g��[kM0��AV��57C�2>sa�)FDB�+���0�[��~VzC��$-7]�1P��D|g,�e��r끰y�<ƛԹgY���Hl�4l'd �
Pd߉�����r���5�������@�n\D<M-�7�t��Yq���?a4F�.�Dlvb�Ȓ$���"�^%*8�*���C�0H��O���1�J�ޅ��
�@��I������B����7T������&�`�o��^Г��N5;6i/��F�)�M&J����}�toi���o�[	d��\<�@5Rn�~Ø�Sf�*�E'�a���q҉��8zhs"��P6�!����տ����d�y{�|W*6��FT��;^܌gb��Lo�F�����{���~���-0��d����]"C?x���s��Vs>��±�}�@鍚��T��"lӏ��%��(���SG:� =���"�����#��M�|;�O���D������	�0}E}	��2 ��&�z)������.�"����4d& ���\R�6��)Yܢ��%�:�H?R�S�q3[��	<w��W8�Xِ�?{�3�b_�T<eb��6ǌ�%�'�ٷ��´�V�,��۷!^��h����R�B
�,;���y3^��x��x��;T%�&I�Ng�֦U�ݩ~�K¥ON���@�ѡ�H/:l�D�&�s�[U�z�5�2l�w{�W|C��\O����n��e��ࡘx�%����� ���Ւ�{q��u>?J����;hLo�v o�ұ�ju3F]�V�s[h�w?��.nGiAk��ñ��@N�IwB��1"��Sm�oU04�і�t�բpw��؍��ݫ��,	��篏1k��&?���tk�yݰL6���Ŭ�T��{�Qe�s�,��Ix)8�q�ԍ��C���hS�CS�(�@�=0^ZT
�N���H/#��;'	��N�#��4Ul�5�Xee�p���/����"�p�S�c��#'3�$�y��6���^�U���0��Ǵ��ԩҌ�$�k�$��@O������ZfZ��DT��t��I'��G.�~	^i���Z��ב�n:��u �PnIVDɱ�Z�}�e5�A���>���:_7��4M��c٪�H!����vh���pT�6e,C�Sˠ1D��l3��>hjա�	��{�����"7��(МeY�M���һ^�ȍ�&���U���]j]���$�c9]As��/֜�������U��HW<=hS�/��<wGj�X�@�ӫU�=:-ޡ� >�Y�0q|�/��Rl��"EGS'=�x?J����MA���DPU�+3!9G�m`~#@����`{Gp�g���ƥ�Z�k�48S�EÒ@OCLJj����%c/���}�J�-|��aoE��5r
R���+�M����ȷҷ����8<0����B6'O�M�r�Ȋ�G��ȍ�N}���?3�WO��_�T������԰&�R��aԄ!)�-v�ُ�����o�\H��p{�BȲ���}UDz�?%��m��b!��RV�y�yFl�l�[��]�����D|Ǘ	Gʼ��g6���cD ��zj�nr���M�6 ����	ϾI�[3�_3%r4�8;�n��%ǧ�Z�ߵ�������Ɵ��
t:d���>wAWd����M0.�%2qxL�hI��b;�=A@R�cJ� ��[+�)�! ׳L��3�-1K����f�M��ּ�ZL�B�$����@4x��[�~2։��(�p�NNJ�uDb�ńy���n�Q^�H���S݋�D�r��r�*Lcڟ�b�u"7��T�>2XL��o����e6m''C'�I�)Mn�����E7�p��=�3[���ѺQ�t_�ш�lD��El�w����*(YRH�N�3�p��g���0��&0m���/m	�:r�W�/_�㙽�F}(����GV���X��E���E@��?6����1�|��6n�u>#ތ�iW|-�njq L_fO�k�a,69=o�#řJ�`�@���˱1u�QQM�c>�����S�3HU�
r��=^�i��bPQÔ ��E^������~ūw�=|���lL�I���a� e�E�=��B �'B����4��􉔵��$3��|��`��W�d���YǦ�E��}N�x�pZB���c :'�X��u�XO~ʜ�z~�$­�Z�J����͠�}p�b(N݁0�����:T�p��%6{�)߫�{Q�i\�LO�꬘n��I�Z��w,$�&�W��
�/(�N@i���5uP;V��j2Ǆ�5��}�zey���R04x)4rF?���@���A�D��[Ya3�c�OU"�q���kV�j)j팺��n��B����\0WZ��e�<sN�l�]���;�_#����!~�6���m�<Th����?�^��J��hPg��V*�g@��)���h��ȱ]�4QQl��t;����	k���@]+`�X}� ���ފ�󼢜x��X����͌z}��;�w����=ă�u���mB�`�z�\F������VL�S�/�Q���8�~���Yci��N��
c`؍�	�_����>�ȳ�CY��e?�ͬ)���ag��x���sY��	�ܪ�� `����z�7�Ӗ5�X��SiYJ�H��O V� ����-���\�dz8qMu��b�a.D�,�U��c'9X�.eu=�z m�5�� F
_��&�CYJ܆.�圪�^����տ��a;�8>e��uEӛf���9U�T����&��X�F�{�*�kB�����I�=?�i�k�U8ݩ�ʲ� ��AQ,������Zpr����4xhet�-j�VNm�����ݱ��e�]ԓ԰�f�����og5\�dQ��N�T��6S�2jll��G�H��5��3��۞��xv^H�nɩ�lC:�8�����w��B	��`k��J�Tzě��(�[U�>Pi�U��y���7��ѯ�o��U�18����:;�KJ�e���J�"�7����X�3 8�tK#��z�;a�IU�G&���4�����wVc������Sg	�_.������� '{���21�V��@�$�BQf�_g��D$�=p�B��$}L��?��4��i�t��A�%�.��1.ѓW�f�1�Ͱ�^fCJ،�;O��6���1�,$b3t�2�鬢�nJ�Z�%ajuF��^� �<�i(�P��y���;����],��ߤ�p�w$����ޜZY�kY�a�V�
��H��Hr�*�o^s_�~&�(u�ˢ^��J�ۉ���C��58���8�b��,���ˤ��'��T)���9����9~�y#Y�futʓ
�����5��>G�K.GJmrj���q�M.,�E�-;����\�@�W#>=�l'W��\%�ڋ ���Xߖ��R���  7˂Ι5���,������q �8{\��S�C��ڗ��(��jy�Q����^�q!��Cc���X�X�4R,��k$N�C�/�Qi����.y�ޛ����NNx��Ĉv�F}��8�j�z���҆����1�V���Cg��1�r�R��hem����=�����Y�=}�u ��r �1��ꔕ�3��eA��=�p� J��Šo�!�09�k����wn�ݭz�����.�K�0Lr#�(�u07-�!�Բ=;�J_��0�R�i�;#IvtS�t�Q����"6mRH��9��N
nb������j����τR� ��b�[�>�k���w������ݣ|�˲���b��_Y�\�ը"���Ӽ�D��ḿ��V�S����I(/m�@W�����B�M8�q����F<��xSp$��]�.��Z�D,���{�g��'^cz5�17�>��|桗��7/_��E���+<X������GY58z�:��u�(���^�H��sc^�k*�,[M$�9u�D^zA��L��2��B�s���\�%�h�jK%Òg�����F�b��߇�f�j�zqי�Av�ٓ:"%$*k��N�����9!K���)gp4|���Ғƶ��� ���r�~P�`|�<���x9=�]].Vu�Y5�$n#����B}Zg�]�D����TsĎR��6h�6���pݶe�м�.$b���:â�S �{��Z��ht_p�Za�ݭ!���͹VI���d�h��e ��Ϭ`�^�bt�8eK܎��W .]�)��΁w?�� � ������d�7c��./	�z�8)M|����.﮷Nzqo��y�OY�)����B�tg�e9X²#�ܽv�=��=�#���3tgMV�0rd��+��G�ꖼ-VlJ�ީ���=
W{��u+t��$2��j���,�՞�g����!����?�>���h`>*3!�{�Q[���]��ťÄ���7C�U�]M\��~4�ef]��0,� �	�dMJ�ֱs���:�=����SŚ�F�sx �Y�)�*��d^��<WiSH(�-=��e��fX��E�ݿ�� |�iB�$��]`��09��C7�Sie(4�ۇ?�C��;�3D@��pTV������*�N5�rI��$�M�14��+���
�8��ke��N��aSƔr���O�]+�IlQ:���R���I��Ң`�'�\H�;���P>�@<[\8ݦ�>>��2Z������.�a�F�%���T��C�������XQ�zO�z�`���oe�^�z�c��c�D*o�w�m�e�+,�}���$I��i�4�]�鞈�;�,�f�n��!���feܨ`봀�X�c嶉dX�h��^�U/z��-�sM���O�����Z�/����1,���=#�8mh�@9k)_H���Μ��w�=n0��L}�W[{����	�\��)���+�|:N�Bӭ�@�eH�ѯ{�X�� }��WW�L��D�~,E搫��������c�-�p����m��(�-l��HOc���D�T���L/v�ӌ&Scӟ�#����ХL�1^��G��x*�����U�>U{��:����z�l(Ռ&�8ܳ~�]qں�P�������a5��t��xA$c��[�Sf�A�2g��b�"�a����z=&/y�m0����Y�����N�0��$�J�R������Ѐl��Vď6�AO�'7T���V���awfʨ9뢂��Ҕ-K��7�q���������;��r��X���c�}��{����A�����9<�"l{�8B:p�\��A��X�v1/���r�B8��c9iZf�Ň.!*�_א�Q�h�V,�6b_$���2:�WX� hˎWl��V�3F5�.<Vfi����_g8�q�P��ZL���L�'�64N.]���ߕ��b˗ֈ��<wA/J���o���#�ǝc?���wj9O�9�Dw����~8���9&Љ�	�wS+�c&]� �#��=���~��[ۄ��s�}�9�ׂ�MD���*3��Kò���5Im}���\M�uG�)d�C�3�Gp�Ȝ�� ���A/���p��~�ya;��s�<	��Ŧ��z����-cU��E�5v�ϸ�=`[�!�Q�u�kߺkv�����O;��l�/'{}0� ��&�<�u��S��Ҕ �Q��b�
���)ڢX�R�)Ќ㢦�%�>gV	$$��MMJ.L�ub+�&�6�ų�U���X�4�1����R��޺S�2t�ɷ<A��Ip����.9��Ϳ�Ɋ	d��4��0D������[gh'$L�14�Å�x.p�}���aL���4O�H�h��&"c����]����o�E��0������3�Ԃ�4��;�|s
0��a�����nJ�<���R^4�
'�d�Wi!��};�iGi4�����J
�r"�-I�b=��u�Gs?�z�����<:$�hlդ~\���Q*��04��!���)+�j�*��ϪաAF��4"�y�RC�V)��_![�Cg�A��[���R�o�-O��xM�_��s�ΫTo1o�u�Q� @|7�\�'}�oD�~�[���#n��~��|p��æqA���;�V�氊5Y���9�z�y���	f��f`r�D��A�'���a�S=�� ���:��`���#���,nTH9"�Vۈ�L;�9���*&�z��P2��/��)�n�9��q��<��~���:x�[s��-͆ȓ�����~�CW���~wO�zP����!�؅�����c�:]�T,�3LQ��dM:�p*LӋU�j������~-�'u�T���K5q^�AԢ@���;��L��uMI�.��;���!�L��^�*@��}w�����<��eC�g@���q!�oϽi���^ƤS��~m���^S�	ys����1H�ڰ���/���a"�^f�n�.���8Z(%\s_�Q�j}_C9��U�ۻ���}�9��#����{�����g ��4�j��@ʎ?��y�������9f��|��譏��I�oVjGA�D��)
K���56��ø�B�����ML|����.LC*޻=��-���BJP�ʒ���Z0[(�TØ�.�*���c̦����*7�CtY��Ѧ�'�OI<���?���:���������%��o��g��kʱ���U
7�)+@��\�hv<9js���A���f}򬀦zy;���E�	�jz�|[<X�3[2>ij�T�ͤ����I/C�u������&w*�tپ)�+܊�ޫ�a����
�'��A�낯n��1V�@fw����B��u�V�x)V�C���\<U���	�m4հ�Z��UT��- ����.��wv�x�s�f^11�D��� �	�]~���Hٿ.��|�T|В�֖��BY�¢MrD}|�M���uۖl�����~4�����c��:��?3I�_%/3����n��;�j�1?��Q�Q-QW�&c[IB�՘�G��<�^�!�S��\��]z WW��d��5�Ψc� >��y�D��������(�fF�sf,n#��R��抈<�l�����m����q��9�D��[�c�:��~�� v����r�L������`O��$�}?h���Y�Eq[��D�fS,x)	y�Wq��~�����CwI� V��K.��ڎ!�m��'EB>�C����p/�O�[�(h5ݭ�(��+,rCަ�=�Z�
N<���!��խ�_�5Ks��7-Y�)62�Īu$~c��y�<���KS�T�d��<��Ұ7�U����E��&��i�Y?�]�m��ћm+Jr&��r��'��C���8��dwAh��ZVx�]�v�L�s��z�O'Q.���_��1��������<��&��i���8`l,9�{˫b�ɰ3�`�$��L<�P s��r+ϳ�qU#oV�-^y�P����*#��nm�ECk����]^Mi�7C]����X��4�  FR�]\����"���\۠�;r�;C���?-^/���x�%53�#����H�-�o��*�0�e�-�9�`S���͕�<���n�ԌT�	):��V9�q2h¥\�͌�j�?��E}����n�ԑѣ4��cY,R��i��.�Ta׷s�%�	��\�[e�>!�N�n��r]��L��㮽T���Ƴ�����d�a�����9-�`��q>S)-�B��|����V�hj�}�<��w���Y�4�:���A����ϲ#�D�;	�"�J�9�v��P?a����Guѯ����x��Z���昳���9��?�� ��Te�iT����j/9ڪ��#���F+�޻,�|0I��m���D�M��JMؼ���&���YlG[�0���Zg�m��?��%]6��=vu����Dr�F6�ڡcX``T�$R�������D���f{(Le7�?y����:(����\�}����������3������TE� �P��B�`M� ?~7{�~b�#�K��ߍ�+r��b���S~�~;0xA^��,�9�<�����	Z%����ruyx&OŴF���>)��|���r�֧K��W�}�G�$�V�~1�K��ҍ�m��5�܏�`W�x1V�#ò.ғl����y�w�˻
'ݰ��"��w5��=��;��j.U9C͵߬�'�8&#q���p�#��*>C�7�%��д�f��o.e\� A������X u��qm _��p���8��)XL��d�}���W�k�x�j��+ �-�n��/e�f�
*u�*(��1	52Sw:(� �}6`�!�gI��D9���[�L�G1QY��2�_�v����a;���Q,uX)躡/_b������}]����=UZv��%G���j��W��#W���AP�x%��h�����x�GNqaX�: *Oc��x�
���F,]�᪖OHj�ӄ�P6} ��+��&�����E�v��UR��vt(�����Η����bVF��,�B����7���om���n�+Bs���+���W^j����z�z���m�C٦�|)ATY�TR����l��_���^Ci��J�P�uvHP��OZ|w�����*��+�)O�r�]S���)p�Ţ��;B���YޫJdc�T �Sj��֮�!K�ȡ�:Zv��Q���c�����v��g ���"�	�7�?vzc����:f��G5�aY=K1�����Y������D^Z]�?`z�6���P���K�y\�'�.��У�A����W-?�=L�(���ɼ� �Ө5i�W/�#V�S4��%�Ȓ�H5�] b���&=ۘ�'���1/�mHH��&�6���U���&~'S�B|�0�2�(0Zy�d �_]���?��X �c�'$��~���u��(��'*����4^03�����y
��-[�Tϳb_�sJ������\S��Y�>��f�9�oℬ ��2���s�_ Sf�-Wp�_��T��~5�Y�S��{���"���i�Ix)�+b3b6?�8��]l����D�jo*��S��C�6sn���/��?
�#PD��:_
�&d	^bg�I�d#��� ��0h�+��8�(¥n����$/f��Pn^ʏu�\��
��Whߢ*�o<�4�NW�ȓ �xV6J�i%�>���+(��<���A�G��9	��j7Yc�S�3�̣�3f���NW��Gv����1$��c���FL��Rc�4�Ϧ�������k
 ݗX��8Y����;��MZJ���R�G҈0j�:��d�F����d��p����-� lѱ��D��\��_���^␽\�O$w�(;��s�P�+�|��h]:6�)�X}�����
Ԝ������j��h�#��\��]��r�)�����?�bUc��0�7��G��X�R}c�yY��F��dϲ�a ;w7�vx��l��8�	K��A���a���5eS ��Η�U� �Jx�`Փk�`����r�8�,�p0>�����k�#��+i��$Ӄ�ji�A����N��Γi��3��cs��V�vaꤌ���T�x��ldM���gsa$Qc�/s����z�̫�r���#���s���`��2@��OC&�i��SN�mdm�rJ��:�@�p�YJ�y�� d��Y2��Z����u\�۸��d#�q-l�w�a/���TR�m�������	�/g��lK\�ƺ(7�p��+��ldu�^cz�x\.ģ��������V�\j�8�/��r�Lf'dO�K �|����G;xfJ�!	�i2�D��,�X�@��SUGa�(����\�;��3�.���{k��tr
M���&��Y{�Op~{�t�˭�2>��}Ǚ����%nԽ.���Xܷ���L�ï����}w�]����e�J�Ţa|��je�5Dw7�B�U��gYj;��A����7G^�u�_�[�+I�a:\LQ�+<�ꤒ���5o{�*v$��(�=�G�^lk��n�ә�H������=b._�~<}�_(�#��/:���b�V,�jt��1ȹ�`-ox�!;�L ��Y�R�4@{1z��ΝUD�����\�`=Wݽ�x�����ݔ�K���<�e���~!�/���b����\]�v -��
6~�4���6W�	(�1�$��Y���R6Ҩ;w�S����`����ٹ��*���H���"	��&�,+-���|������W
l��J-����Х���S��e+�pK�y�l�I�1�b՝!:�Pw�����k�m�8Y��;�;5���;+F:�_�+�����7�jXTň�R�LbY�GG)A�5 l>��/
!B/j�ν85Ke֐�K"as��7Y�,,�ї��o>2ִ�*
�����~�%�B�	�V�J�'��Q���{���tGvH�P'�S+�I��!���N:�Y�ow"�z��b"�o�}�ф �[ݿ}E�Й<=�e$�����:k�`�������I�R���ا�f�8աFzl��K+���1힤�'!N#㍐X6i��a��t������zR� �2���N���~��E�K��.i*R����CI$V� t!��	7�E�R�>3�6�1ق�`2����oN��|�q��0�V%~�0�Y��ĸ;��}�:����5����ooՠQpU����Xut�f��eM{�oj�A�������h/	��8����zu���`>w�(Y)��+2��o�w��.n3��&��P(��?���i�Y[��E �2���D��Pƻ�G����<:�ϡ���aS~�42I�� =��0�U����<z��ޣ��O�/*<��	�%�tp+��3SEnu
�HE�i˟al?�%����&+0H5��2�����v�&�o)f�O�tt��/�����{����k�zb����ă�k���Y���椋6��D��K����8?���a#}�b2'��:�dv~��
�����Im���=&z��d��uJW���jr`59T������Rĳ7���ሮ�cKp6�E�V�S�4���4��n�ʖ��%z��脅�����Zm�a�E�dn����*���+�;����B��.��du�]mA~�R%T��̋�竉���˿s�X1?T�׺�y���Μŀ�_*�[�%k	9O����=���ܭ���G{#�V�[�f�����>5���'�Dw
�l�C""c|�7\��\�Ӿ׼���@��`�:9v�7`���>`�Y�iA5	�*�\��5m���m�Ŭse��ѝ`x3�@�9�k�V���/1d'i�p��=�˲t��c	�sݵ.%��ո~�sǮw��8ً/M~T�Q���,T�Q��r6/��չޚ�\�О�c���T>�ϻ��ͯ���z�J��Gʭj<��7��}�ۊ9F�)M����|��?K[��bN'�=��\m ��dE��T���wd�@����Rs �56��u���][����d7���ɐ�fD�]�  R���*����3�?/���ŊPUз�������������w�<��k�/��ᱢ`���"�OC�c]���P+Բ�u!rZ��	*�=yR�BD����G�[�Mb[#��Pݘ��ą@��|�J��ڎ�Y�F��&.02Q.�]h����ē|�ș����+�x����VMhb��~T���xJ��|y"�\׍�Jl�qG)�	����Qj!�;^	�]�}��`&��]� �L?h�oќ¢���y�Mn�3�T�s1g�"]Quy>�c�i��Y��C�(���l�=�(�z=�gak+^<M,��F�ifP�./�|��*�ٷj�N���o�Q�&�{K�SZ  i�Y���7tΦ'c$�E�ƫ�C��zF�G~<����ު�M:F�8���`��N�y!ߝ�	*�h`����vIM3��ͷz�o4��M�)����^�_��Ժց�tzZA�+#�����@ޛ6Yky�P��J�0�$���oV$�kn����!N�8�N���GK@QǶR�����u���c<���u��T�v��X>I^Ke:	&�[L�o�.H�"ܑT|�S��ܥj�\Z�Z-�J�Ī�����t_;��5I�"s{(+j��PQ釺��m��	o�+�B1Gm7[��_�x�
\��*�s�#�����]���J�?����WB�����% ,2W��݄����	�vC��5-�����O�N!��f5��4��M0�Rj��[-�JG�1a�p]?��K��o�
;'J3I�e�e2|�} H���S5��Q�4rq��`�\��KU��-��$mN���C��3D��*˴u� CK�ف����Ge7�/�>�y����VN_��B��YFҬ�d.
u��J���s��Nn���k.��.�/&Z\t#Vzn�ho&T��A�x̫���M��@R��~dd���t�d`OM���! ����)�]�"x>m��}��)�h��"Y������+��W4��~d������reQ��Q��tTh�QI�8+�N]S�8P���Z��L7�����!���f�����7�'�p�p���v���7����O��''e)ә���|�7�_@��*W	J�����$��;+��� )&ʽ���y��rR�}l:h���� �;UXR ����4�1s��g&3�BH��4k��|�N`��O�`C��i��Ń4_p�'�Ds�l�1�6�_�@_�2E�"�;�8�����sN~��%1oEY�������J�r���cE�K���l���G��6bh�ڌ�:wܛ4�S��W�Ş�qT��{1���\;)}r��ʢ��ԠvL� � 9��ҟkH9ɶ�׶���`�ͻ(R;���A"��ƹi�ޭ���d5Õ��n��(h� ���D]������f��Z4��q ׉dtD:��qC"�
�����^�	w��#9���j�1��G��%+wp;�Pӆ�j�[/�O���� �H
� ?+�v��X���v��.S8j�r5��Ӕ7<�./)�Ǭ��X|,��NU�ӄ���}�:Mi�5_��gB0�OZw��WZ��)Q/�z��d���UO�\�{4��Em�ff��U
٫�E�#uS���O;�L ��۵�d�£Y��#�H
ɬ&�*�̌�4��g!���4���`�i#Ъ�i$3�h�!��Fl*%�~�b�剟R6����֋�K쎬t]��:��%���l�,_����OȢ9p��t�䵑�L�J&�z�
'�a[d��3$}jIj`��n��Xl��
S��� p�~���l۠=�Ho9�e�u�@1�N�s(�MIu4����v8N��!	��U�w���J������*���T����g��HU{��t����f�9 �2�1��AL5�랤�mcp���I�d�K"ٖT�W�C[xs1�P�-VVk���� �@���s�Pk���=�^��|��a�3:��)�J�3k���S����c���IF��_�]k3��
,<�.�ϼD+~�Dv.s���濒?��`�m%'��-�R,[nYW��nhSbp.�@�?éQ�c첾/� �B�u�Ip��ų}�� 5�����i����]�3��5���3 [�M'����Pc�d6�j��ܞ��r��d���O ;��1G+�@�A���&� ��
�Wh�e^�ݕ7v�n�>�p#�-��I��x���8�	.:��i�~'DN�f��FZm���%a�t���E�t���P�]{���!�y�Z(/��<}6���u;�bf�#W����`uI�4�:�aT=�^�Ar4�u�k�������E^���d�cF��hb;�ݛ Z�0 �B�S�[�υ��	#ж��;�V;�c0@Md�w�� p��g��j�F;�����r�K�0��#��>@V�'��8^���)�_��>�w��+�]=�eK�-k��Kp�׷��?�Ĩ~=�^Q�̝�+tiT2���'���!��R(d�I&Qh�C���X_�ج��{x#�b���;��%�b���$�g6Қ��x�Y��~Ej�Yぇ|�n�]�^������s�z������w���zR<��[1��M ��:y�p�8]��'�{f��T����9g�4!k�I�Zď}��𔠳� �� �����_^�\�"�.��-4ƘRi��N��ѝ�j*��΢����� �x�t�i��d�":��k��L�Ij�Һָ{�������@2��To��!`�T��+�'��}��"ӌ��L�m�����'�޻�A:0�9v �Hi��⪼i����K�����}�a�9�&[ڜd�[��o�yi����� ��⠭�`� n8\���S��֔�k�囵����{m�Ԉ���#	�bCZ$z���:�1�n�%,�8�;�AԠ�#R��Z��Z��P��7f�e:����[�{cқ��LN���w�3�ROZ:�`hCi��u_~vj�
L����l�f��(�*�?��;��_A<���� `�M���8�E/i2�)�������x���� ³q:�����K6��˖��*Yٿ�y���=�!8�����%K�(Ge�`Y4����?j��؊FI5��f�~����p<v�'��%c`�n��P��v�6ַ�~�6������`!_c����˧���$���[21�:&�!����oe#JP4�ۗ���+Lem�q�}{�*C����p�Y�9,��`�&��l<���ZFtЏ�	����9��l���+r��a�
or��t;��Pː�-�������I�a�ܤ.��ĄGl�r2��9��L1
bh��J��t�5�.}�����\O�c�q��[q����^�#⭉AO�x�ƽ�zQ����{CXd�L���}��v���b�qQ����ܚf0"*�$����&K����Z�Wa=R�B���/@���z��ý5�R���12c����dC�x�*�� ���@e)�?������<���
D�}���_M�m�7.�7�&��^�`���L͜4�ܻy�W��{���+j�O�魾Q��Y�?��(��u>���L1J{���vi�/P:Sg�`(�g�uÖ����E{��A�,����U�'q�_-��Y��{���O��<�d��0GN�1�,��#�栯���2Du�߲?7S���7E��̜��4"m����u�y&{`B4e�|/�M�(S����z݄5{��
��}Hx�T�~��6�(�뉖�]K'����W���։��n8}]�pq�ͅm��{�v�gp�r�R�`�N�4�D+_
����U��XäbM?��Dz#w'�[�p�h��(��Br�W��w��9K���3AB|���`���</ ^�s���Fy��4c)�2�yQb-\y &�l�jղ�oD,r�����,��'�zv�?�ھL�ŵ�ΧuP����gm0���ڈ�����X��w�������Jg�^*�rlB��\K4g�Lb��\��ONȖP4��EB��:��,�I��d/�jN�p��D��N��彖3�t%�|��o���C��O|ӷ6��bV��\����ڀ��eTE���lrD��⤡�e"/�@v=���1mT�������d��~�V�8�����=��^>���ǐe8NΨkEv���R�DKM6U�ے����p��4e�QN�`�v6�:��=y�tש��8g��L#��m(!I���F��o�]yٵr�� ��BdJ�F�ְOur��K\"��-aG�� ���X�g�C{g�����-}�\�/��X����σꔡ;f(��d��G.�O�,�i�H�������"<��D9Ws�q-��RCu���N3��}�T�0��3WC0G�����	�o����6�4����"���=�2G�ܮ#��^T7}pþv ��eI :��68>;��j�j�&�q�� S��&cOOr�5���wzc�[����e{��y���[m�#�T�|u��׀���V������ũ��*W�r	�6��8��y�Al��3q�M�ξ�">[�y�[�|������Ȝ���w��*�*�tc��'��Wd��ĥ������L��Ǟ[^���MIzv48�.R#6U2�ꄪǻv�[*���j���S�I�=��Ѩ���'\��;�$	��o��Y7^�����0�P���rIB�I�n�-h��þ�WU�f�Ө��Ju�wa~��f�d�C�]��C܈]���pE$"�~a�6�^&hT]��{����B���x��j�����`������B�S¾>낋������i�U��5�b%n�27S�xe�ن��ŏ�����M��J��iu��1 R�����p%P3�|K:]�?��V�=�~m�͌S%�M���t_Ǣo�O���/O�� ��@p���Ju�$]�=v�Aׇg����EI��p"Y�B�F���Bш�.El+�U9[G�O#�ԴV���$�h_L��eR���*Z&vx28�}>�oi�ߨI��	�:�� �Q���3W^=R�z/��H�68 T�yFk݁�ӶXSE���X�����t�q-'Q���nӶ�~;�'�9�ӯ@��L������P�)89&Z��RcT`��Q���w�G��շ<���+� 	���5��}�����p��ݺ�t���%{�ˊgڱ����߃k�1��OJJ��Gr�BSIv��V\wD]���Ca�dy婕�@�I�A�&�J��,e���މ���>2�H�?��0�O눧��n���u3���q�V��O���Y��$�J|ɝ����R��o7W��G+�;�C�,5hɊ:	Q����IF�V�;,ZL0��p��Ǆ.;5�fD�7�&QZ��4Т���5�tH� �߼�DK&�=���3��җ��X����7�����J�|�C����էޫ�7���d����ib3]�!�a	��_�8�3����B�,�T��o�!c�e��!5�*y~��(W{tK٢�iDC��@;e�yxb�y\_#�8^K��0i~IgUOWE-��O�$:u[T�S+5�81ʜn�s����"�1T�w���Ǆ����4���K�VH�i؝W��cCV�m"�� ꌐ�a��J���T��A��q�p����F�!�6ql)S��M{��+��%qC�d�Ba��ʷ��$]��5�"}>��BEJ+�*R�m��o�F�%U�1B�r��{J�5���륯���N�����W�"C.l*��I5�D~4s���;C:��H�MGQ����"���}K_b�%KKSe�ڮ5A
M)<U��4yK i��`�	h�h�ې��brΧXqm�d6;�����dgUZg?�qՊ��6��Ji7̶����:��e��.�=�AOǂ�TB���pۍK��̌A�����X0w�Z���<�Z*�F�jlJ�ǁ���!��{1�z��#(lOaD��v����;`"*̑+�=Gl�z��^��+]>/cS����.�z:�n|��.Z�X�'-> 3L�z�)rne�{��b��0�~Q����������bQ�����؞�B"a�9q������oSg�(�p��S��0V����?�
>;��_`3;��n�#N��W��+|�v�`���g�����0��W��=�aH��!� BvL:�z�C\��3L}���:_Uq�m[S�y;@���[�U�E�d�`�C�v�n����(�_m=�iҾ�D��� E�PL�5�f�n��MY�U���Y�%N�h�g	ׯS���88��1��?�э��e�q�?�T��n�;�ܾW��3)���Q�r}���D��Bw�7��4f�yZqW���i�V9���:��`Vd�V�N��~����>���Q�֗l��w�rg=��2��iJ��*��0�����+�EEb��g4�U����~��ݣ�Z�YY�θ^͇+�Lþ@<�y����j�9r�2�M���&�`>���h�M{2-脾�Ѱz�ܨ5�f�*:3zh�"��b��0缽j4Y7�_�>��R4�V���#�Ҳ��̆�x]�$mh7�1�4q�յѢP���}֚v�u'f�gQsx�	k��c;�\��v�_EEwiV�>`S��X�Z�ƽ*r/������G�:EZ0���Z��+G���RI�K���R*l4��� ��U������C9��G�r"��{��֐�FY�Qc�٪�"6�= �1-��#���#����agC��8<$�5�]6z^dO�g�褐��vg��s�D�lf���`q����p�(<�;᫿�k����H�j��K�Ԭ�������� \��&m�}�E�9� �l��^�Ʀ�t�	id+	�g��Q)�8�\'�v��Z�N�z���瞗W�q1(�ٚ�F���f���A�Y�5��!�g"�?%���6�|F�����%b}$�^�̖���۟o2�Ƕ,��*�O;FtGr���*�Wm� ��p����j������&ۗa��tƪ�Uwz��5���,/�c�y�e�fSԋ�֜��vL�.	���A@��`�6 C���c@�x���_gc���mU�(�U��� �V�$|����A��+�:X+_.4�g�'�Q��<�3�Ȫ�ȋ��}���솅a����#m�P\��ii�sQ���
-"eZ�܍۹l�F�8�I����1zD���2cl�Z�i�>�>�>0#�0���ŝ)�H�OG�o�Bn�3DO�$�����w���2��GF�,�V8�
J
,�_U]r���#�=y�A��3`V��x{��*+vj�(�ҵPL|5���E�S�J`_�Ñ�C髬�*�h.1��s��CRx6�X}	�)��++-�xo	�����`j�"��+R8���M�t����(7������a������-X��U�\��^����s�W� ᘽUI�=��鏢��C��Õ�`X�S}
�П_�DQV��*ؐ��[d��<�^ٗ�Ôոko^�K#/�2�x������4�����j�4SJb�R��#��V>�H,j��/씆F��+X���P�N)s� z�ݳE�&��^G�q�Hdkq���v��k���x�ϏR/��0CK��ND�H�ba�����_=k��>[ߋ�%�6�@>�|B(��|�VN�&�׾A:��b��=A��>_۞�ѐ��}���1-ˢ��60!>z8��.H����S۩��7@���-��;�6�r}�OnLH$n�s2�!��),���#�S�g���#�;��s�N,���r+C� 
�x�{��`+z.�1�L��(ReI��¶k�Sf\*t�[f����J^�}uUM%��"A�dOq�.g1=��!�3������$�ܤq�����cOߚ�����8��d��;���8�㙦�W\�<x����j��;��f�������K��_�u��i�0��_e�*�M�K�����0��o�E��qC؆���#�?�3�(��/�	�	���u��(� M�)��U..�hv�#�`_�ab����*,	���+�-i�h
�N	J��:~���h0�/$,�=�{�-����B��I��-lX���-�I iׂ&�9H��ϛ�l{�dT�m_:�̵�*T������t��%"��%���=�zq���&<��d!���r~.��R��A���*�C�m��D�[q���R����[XM Q,E��E�Oh��wFe�pu��V6�Y���=˛g���;t'�-��g
��GK���|燘%��2E�)�2�dƋAC*���P�`Ϫ4��8^�Me�����݌~���\����˧r[yM]d�ދ�B]��I�4>b��G�L�D����~H�����G�'l)&c�ᕦ`�r�a\����Z��m���x/�0��:�G �;.��������oa�)%(����.a�#�[K�}DJ����H��)�!��\�hʵ.��&+t0��|��vl&�ɞ�����o�� �(��z��e����jQ�>�Փ�=}�����2§5�8�r�DлJz����5 �(]�zo.���\(m���-�ZT2�f�T���(������jAC7	ng~�%�-.��Ye��J������+�O:�2����R��K
���T�o8Z:B�L�\j��yiv�m2��L�\��#�]1��ԡ_8�T6;�֙?^�z�1]�����Q�<�`�h(0�:p�灥�|���K��ȣ�Ư=��Y�7�B��l>�YZJ����0R��X2!)�(�T!���[v��ۼ"��i�[v��>;�4D�S�`��q�B� O�N�ar���Ep�1wb�-��枢�������ѫt��'�go��F����^��9@ƒ��������ȦC�]"~���2	��N]}#KQ#q�m/���#�����_��+��d𭲺�=��\K�#$�]+�0���խ"ŗ�֓s�(��6�v�_r�$��{�[隆�����\��T�K��z6/`v�\F���KS���P1W`�f���㲡Q�O4��œ1=�yy̅��}���C;,owQ�9��QJ���~���5�������H�~��̡�?���S�dM���Ir=�7�W1���tl��H]1\�f

�����MY��J"0S(��'�Kh�d<��G��� �^�m2$��eL�D��霠�y΋m⾴���������a��I��i�A�PRc��1���][�A��Yz3�Oa�gi��v�U[Ux~�O���
�g� ��NƠ��2�h�u�ǳ}�w�7�?�B��k��I YU6�m�:8};���Zߴ�1���XV<a������M����kh��m�|�&��!uCo5�ܦmv�j�GuHۺ�gXՖw&�k��1�ѡ�eKGԏ��ўиR�GM�,Ф�VY�	�x����t�Q��.�N���Gw��-|$��ٲ�rt�)�u�l���&�HZ6G���Tn��*C8�7�~ۊmiAc:���t�웠�'/����u�@���������6{�G��@>��=w��l��k��U~���q,b�Ha}���U�$����K��P3q����H7��y����*ܬ�63?���9�n�ڽ8|E'\17
Cw9ŏv��o�l��g�,�A�]L��yx7�V�#-��5앳���I����Ծ���n�
G��#��vaS�/���d�+Y�ߤ$[I��$d��- ��dD�/uZ�5]q�9	�ue-t)�4$���o�R��h𗌗��I�jrjG�~� .�WA� ��T׾�K"���7�\�������eXܾ�\	�ګ����qI�Α�h%����e	�e������2��O5RCJ�J����N("�gG�jmϸ����C��S/Gʝ�I�!jJ���_[���ΰJ%���Uљy����@�v��l[��u��ky�f؁�+I�>q���F;e�~��)���f"{�t��O�85Bâ�r<g�=�Ч>Ȱ�}�U_$��"��d���\ƻ���&� �=UQ���?h�m��U�w�z&����Mkֽ�@,�R��͚1~�3Y���hP����zq��Hƺ��1Ȏ4h�F�����I�zL�/�@kXH/���Ăi�Etu�� �_��Ǹ���������J��Ӌ�^�؀U"��[W�/S��!-��e)|!�!ٿ��"s�c�Co�_��j�'<���G�̺�~y�9�,z�w�-$�p$$[��(�g:)�ےf�DYvH)�m4f
:5:2�>O�rI����]�5�=�Z(��YK��
�*�j'`�}��Q��C�W]��a�m��l�6��*�ֹ3�v�ߤ�GΗ�BO+��8D��G>�D�xz�WN�EcB���X�UW;p�r	� ������]㬁N^6Ÿ��h(L[����Ꝕ�څ&o�`F�s��^�xE5n���ŋGX͝u�9��������ؒo��RS-��d��N�� hF���M�u������G�	�
�Cǁ*� d��4��s����,S��導Tv���ߦ����(�^��jwk��0�����
h�����H�9
���W�e��Ѡ,Œ~xEWZO��G-�����>�dN7SMz���{yxo �]a���m�IݻG3e��{�NU�����#b�]8�E�˿l	��&�t	Q6!L)P��c�ٝ=�W��o��IQ�dԜ{�X%��c�� ���6�����9e�޼��+�A�W��;��)��pP�2��?�"��,&r�(����������;��F!ꞝI���C�ت�C��
m�����9%�X��BV�}�;�D���I\�T`��V�� ��� ��5�������������G����7���H�{B�Xr7��D�#U��^&��3Q.~Ws_#��<�{f"�P�G7ƭ_�2%����!>$���075>����c�CȌ=�=@jٱŖ�����8Ƕ�MUtej� w��h䒼ë�,�K�?�׺� 
�A����C��X����O�FUz������j�Y�c��=�8�c�##���P[��T9�Ik^c�93A��ܔ���O>�ҌǛ-)��/f�s<��Ix�[f<%'��g�E�/h���|�d"��)��|��0���dfr^S��2f���
V)�s�5��I�e�[����8�����ަX~n���|yGə�X��l�1X�W?@g��Vx�g ��x��1�M7w�	6)�HzV��g�G��ȁ_�㪭�$QiJ��B�����LrOV2���O�-��c8�a��gH!����q0V E�#����5|�ūk+��8�����܈���Z8�a�2g�I�>.���*q��}��OG��%��ػ
����nG)ޱ����%����܎xd~/@�2Y��+�7�U_�������_�Z`�4�9���0M�̇[���d ��HIQb�w��<���ч��Ȯ���ɳ��%�Z:�9y⍮�\��U��M�y,A{�G���#\�����	ȏ+/���G� p�h	Eh����}�@ΉG��H��Ae���ʘv����0~��1���vi������z,I'�Y��Ա������<�MƞgIq��ό�ò��:�f_�.���vxn��n���ӑ����w5������^���\d}����62�@�$�桘�\\G�u���y ��qO=��ڮ#%o����ty�^!D��#�ǭ�I�
�CF��| ��kWn�=�{����z��,�iq�[�*6��,�����T����VJ ���w���z;,��<�Db��h)貜�"����da�m�>b�J?6�����v�Ԧ�s���h��Cн�fV����<I�����&���{�/dMB�r��O�^�i3���n[x`�[\���x��n�-	���{)N�+m�+S�Â.�'.x��p8��}��+�tY�	��<�ix ,�xU�<�7�)��K	� ���N���-|��&���1?}�������b��W8�R���h�V���R�j&N4��F��R��#��:�L�cT���i�m�q$������dB 0<P�K3��8�IL���ҫ��1���ޯ�XS⽞���r$ӈ׷$ò�p�:E �ǿp�[�X��+��$�-\�_��?�q�3k]��Y��D��Z s�aA$�Ju_6���E=�x�aya�gv�#\p�ݣ��+B����, �L*:��i= ��P�
h��yC���Ԅx�~��K��Y���d��5�a�bsG����3��6<D���w�
Ԕ[9ͩ�xyQ�8�L�]�^m��5��/�t��g���58�TG�윣_��"��=}�r������by��"דE�&E�����{�kfm���O���%�ws�I;�@�����̗���f%7}m��[E3ģ��M����!P��X#��U�!�s���#Pkx�푒�A��d���x���7K�E���l<�I�6&A}���;TI����4.�`'ǰ =a����Z��bVBO�k�Q�eB�`G��%G�X(ॸ��;��A=���_qU��u��4�Jf���N�v4ScVE���p����S�]�zU(l3�Z��8%>�\�gT<y
�8H�oɟu��"�c%���>M}D0��/��th��U�7]�6�}eӀ��� @�n7+�5�ӣnuw	�i�1[�$A.At-o_�9����б@� 膳<$��W�^��x̓��ޖSS3�]��Qx��SYtw�9�ЩR�j�?b)(=��A?��ʚ���T�����*����$�$�D,��m�DAn(�S;�� �+��A�N�I&c<��.0��|7><����� #���o��l��VUv��� M�������n�i�i@L1�����ӠDS��� N����
͍��O�ڱ�o�>	���G�9��Ǟ�z���0
j[�\5�_u�ɱC����_2��w�XχZ��K�c�Ϭ�j���Y����0Γ'k9�����4$VPa�������fEnE��T,���A��7q�H�`��/�ԟҿEc���-�>SO`ct������Aj�;��Q�' !{~�>��g	gdt5&//{���t�'˫<��u�U!�K?;e�R�(��e�Ѣ�,�MB `?��:�+:ֶ�<,C�6�+����1����˷��1������'5�a�l ����y�@�{Y�� cp�[x���H�0�Q�|_H����Qc�3.�̒*'q,b�οu�r���v�Ȃ�~Q_�.�k|9d��&��XMVU�����(�`���s���?���}`ڞ�?���N��DjC�����wʮS���G{�>�<~�z1>ae�u����w�l@�Q��S�f�����a�A�b�B�K-�7Sʏ�r^5����������z��U ��ﯡ�7޼��_JL4A��%�r=�YcK@�3���Z{�޷�7�;V
B�j�^pX�b�̵r`C��e���}������6H����1�����H�2��������۝�l�#TVw�����v�꫗Si�/3��9Ü9�zn�U;��z �HB�8⤫G][�	N�w�����I��fg������},�|�[��@���]r�^H����&i~J��X5<H���
�ƶ#~z�[A�X[Wk�[_0֡˨-����K���.����4��g'�Y�>����v`�q��L�������=˝���	{�q�i2��3+�*��|m�|?H��I�<��W$��Sv悳�.���j � ��D��Z���6����J��dx��j���
앧z����տH:O���,f�]\{�V��<>�l0�uy�X>g�PA�C�L5�Y�Y
�15�b^�0꾻��@~jR/�#=���X�aM�<�L�)�Dk��f�*fߌ
�G��=�>�Ι�p�2Ģ���~���n���R$�a���C8v=T��<@������
��� ��U�i"�����lb�~(��1wVkA��b�]%ܛR$z�Fus�"o�J�8]��5���<�[��C 	��Wk�o�� �Né2~l�=��\V��kK���ȼX��OL'�3m!Vs s��^��e�?�dn �2p�(���T[ڽ� ��o�UFX�5YM@7
�����xH0������רs�{�n�H����*i�m���ֶ)��`Dq�䊣o�B����ɾ5��VXj@�;�S��j�)d��`;H) 'o��[���d鼻�.���r+��&�����\���d��1����1,:�O+�����Q(������'XW��9��1���p��ޑ8F?M�����OEw�s�2�M���c�,0F* ����m���r�]�bW�K��=��\W��ܻ%���ƖOȑo�/qz�Rn*6�m��0Mnr�{�	;�9�[��V�W���)���UqΌ!�ɡ9�
�m-8�/~��⎏G��.Y���ʆo����c�=?
!Z䇰X*!��vn��$�i_�la�0�GPh;v��[�m�3A$S��Nd\��H�	�uw�#�.;���K�~��B�?Q����ٔ`U섬��r�%ՄT���!<������@`3�� CO��F�|LWbb��г�|�
_Qt�-~|�雇 [�k�盩�L�h��5�I��x�*a}����GH��F5A��a\�,�>�>.ЦT��it��i:���o�x5I����)=J��P��)�*�'5j�V�I=#R�� �h�~�/�����t��~q�\Iu�����[�A��7Pv�Y5��
���r���Н��?��X��D��O�~h��l (�������f?j��
�~���5����f�ʡ�->%뾁�G��n�14�Rjj�b�3Άo�(��Q��2� �/]�p��g��{�YA � �g�<#�Ī�n�Z��jY��f~�2C#�wĸnE�����ֹ�vkH���>����+WS����M5T&X7��f��v�B���X�nL�%k�[�̓ǋ��7�KmU�#w=������!R~��$-�B~�˨r�-�����-Q���I��NA�}��g1ǔ�s$�&-����6@�k���
�){��G�1�gn���I[����vN˧ډ��[˄����u4�ea��)��gu�:�ܘե��G�ɽ�� �D!�߱݌�������2�W�]��	�坝e���ci@��x�W�yK�kUt�
�ežB8�3e��i)��}�Y�hĳ�(�chz3���z�a+����r'x�����2E����@`Y���|g�2n�a+�PG��0� ��y5B�m=x�| ��3�����?v#���h�.����N��΢L-��M�-��� 0��M��碋� }?��ƒh��eqߓ�_��.�@O8���q���12wM���K� �:�P'�|�r\;����"�"���}�%Y�7�L��7%Z�}>z���]�66��x�X�`nư�������'*n�QDA&���6(��Z��5��✔.F��.[�Uf�Uz�����r�� ���4�{
��� ��s�CQ�0��:of�_�c�<�;I���kL�i�
��=��0�bN�)C<�)Ukި0�S�vDbmi�\f%w����}X��.K�R>�ަ��;"�+uI��U,#�ǖ�"W�P�������\�/�7m��)�Qf�Zk� k����6,�և��6�c(����������߉�OM��Y�?S��{ʤ�V2�rlGoB�	S6����0h�,� &%���3(�q��K��1U�l�E6������]�v�/�"��3�?VI6��/�)Ɣӣ\i ��c�˼w��7����b� 뱪҅�+��hXK�M�J�)�'_��>F��J�V*�ÚŻ�/~�*�jņK)���u�a;���u�2nH�t��!�� �g��wn�{��7�<�~uMDmZL�O�5��������-�뾺�I�E=�ae���h=�c��.<hDI��dL�G������`�.���M}0D�yq���IN�E�࿢׽���"Dk%ڇ`0����]���ڀ�w�(38V.�t�������۳��y��c�V�p�0�.Zn�50[Y��;n?���:D�S~���3�t:
��2����[�K )b̘��[�t�%�i!Ȓ�g�t�ϛ�	��5�!�IW�m���t��y(Yb�Hw�ܨ�+�+��o�rOq��
����)k�ڂ=�˗��OT�����&���
B̝p`���{J�	��^�k�V����ׄ��/L�������Amز�I\�d�������E%�Oc��b�NM���N�2�ԟ^2�l���m���rF����ᢶ�x�NLi��ú!}k�.�J�',Q�o��l�(	7��n~��60��]B��3��~gdh���@����iC�jUP�f��t�V�+�PJA��¯�3c؉��� �p���4=�ő��mf'RT�w	ڷ\a���´H�2)J�;
*��U�ɧ�ֻ��|�������ע�+0��R�^��+����b��εs��/O%�K�d�N�s#n��Xlz�<���r�E[�ନ�LC�͂�6:���ib��˟h��f�Й��Z>�8�p��F�"ș.�λt�HQX(�myƔ���7!�Li���� ��
��Y���+�ӑ6��t�iXr���V��WQ5���Ə&��7���v*S�0���Ålm��hrp��9���-xġ �@�W�Q��8�.����fk�gޯʨ��v�7F�U�M���b=�	@x\�5N���ߙ�1+k6Έ���"�PR(�j�� t��>W5��3�����P��yD��:�Ƨ�:��%H�f��ᇳ���p^���/���|GX��0r�̑�
#r�{ѵwͧn9��:ᩏ����_�|��l7�Mc����QR� W�&���z�FL҃èF*��.���};�$:>i�ҚU��	g���}�	�0�ī(�d�����F޹�ՠp���µ�ړQeeю���4d�� W��;$�� %�'�l�>�.{�A0��S�T�*<źB�!A$'��x
�@�1�*D�����i�Z	���6g���L�4�i��t7����?j����p�A����q��R��:��g�-] �T���x�xQ��>�=��Sg� ҙ�<P�#��J����_|���[��?���=��+�(�mK�)�	36�Tf�U��~�AB��&�c�#�|���UxZٻ�?�[/����.��������6*H'��>�0�CD�fm$} �#��lEĲ��`j�����BSM�(�01a��I�m���������]S�E����>ę�����>M%��.p�v��n<���^�}�I�1�]�:�2�iF�����-���Ht��o�~�t:	�#��b�1�;L��*C�S<�T��_�d��g��l-�fN��C�3K�Z���B��R�h�a/�L(p�Q�ș�P؀��^�xV!�D�b�$��b�hL�{J8�6��،���М��6�V�QT_Qd�w�1T�2˽��*�.�l��Ͷ���o9��Y��M�yY|�?瘥�Ǡ�2CU�{�92�8F7��s�^0\���F��ݲc4PI(c�}�>��,ygκxV�I޵���|l?c?A���S�@�Ù�m�Pպ�@I�Hi<?��D�j$j��d�|ܜ���!�m2)�ǭ9>pE�U�z�cr[ĤZ�eU]�,�W��ܓJ$`d�W%���A���2�q�L�¨C%�T�R��s���� ��67���*zT����p��FsO��:YEĖ�̼cN�4��z���I�"���L�F	��vs~���C4��2��r����ڢ�!NVXPY�p��>���({%�3�S8u�K��A�F������4,D�Vp-��7Z���(͌�=��,x�[�A����Nӕ���}�$Z�7��72Y�q�B����<��A�}'F��q/Zp�Z��>[ �{+l0ȤAX�r��E�8B	��P<�(�^Iz*�CM���`D
�_^����Fqu�� z5�!m)yWn��FD�5O��hK�'e�!3����tQGH!օz�~e����xɂ��Jp̴�c@^���HoG��/FH޵����(\^�_t�%,V9�+��FEk�Q쯁14�h�[\��OA���F�tm�y{o����jgى���U��9@��a8���47���2B�:��D��Rl����A���[ P�Q�`K�0��d])�n\�D�zv��	zV�Q=��`�(9�B�����;8vt�Q|�/�a�,��~�V�����s畑���Ս[���X�9M`�.<|{@+�@:Q ]�C��L}�K<H&ˈ*����SCe5b���7�d�$0����g�g�K`�A��k���)�\7~�c3K���шx����CX[�Nãޫ�{�^��h��+C"^Hz��k���_�s|x�Vt�Du�;�,_�h�"K����'Er`l�`������R`֖@#����df�s�銺1&Y�����gd�9?9�ד�6���2�L��>
��I���*\y:Q���*�ʮ��^Ї�_���>�_�v��IU
3�h�o���h��d��Jw����s7t�*WV}��]g��N㤆���T*��ʽ!�$���y�'�����Q�%��U����"��tV�i��
z���a���9��{���:�yAF�<�EJ�� �y�w抏2	r(4k�ėE~�9#>j����>��Ԭ�_˚�T1JW�S�;��O"�ޛ���������+�m��,�^(< �G�����ߑ��rPS�<�'�oHv�)n|���ƹ#�����i�pk�>��D+eB]�x��EQ������,M'N�$��6X��<R��!iAb���`I����燨��f��ű٪Aq?����Z��LE{�{����Sl�k��x=4�1��d�N#��"��R,ad[���N;��c�P̜�G��F�;-��OX�_�V��yp��~J�1�fX A�c�Ż�))�9RL��@>��x�xĈH�<A�];�FLe�p繫:��#����~b.US��?Q�7�X�e[u����u/��oMN�A���_����]���G	���B�o7G}��f|�{�NG[+�Ӛ5�-��Ԁ��f� ������3m��ˏ��?�_.Hj6D��}9Y�D��~�o�/���K�NGu��2�*Q����v��ҙ��<sS���R" &F�x@�d+>n�HBi`�1��޸Gv����7�����e8d�}ye�mϺnR���p��]���r�3��m�Q0!a�m!;o[Go�<en�э��E;��cR춺���>�%��Vڂ�zxu�n�;HXq�W�` �������Y=�C2���b�d��FM%:�8G~�����j]_�[�3�}�e��qԞwd�p��;�
�b�=?')SϚh�FfT� �ז��j,�ް���U�#�aAzL���0;vÃ��Ή�o�q�i���Q� �X�"Q��W(��ҁ�7:r�UfĂ���$O!��Lz�= ��)D�F9�u�������yT�O�,�\_���W�5�um��
L��y��F{�g���k(� �P���gK�4b�gz�Op�&U ����:
1�-�<L�D�q(5�o҇�諥�u��	���"��M.Gl1W�V)�=�Ͽv�F�8��\�i^佭���܈�8B��@x�]��\�c��;�,nb��P�K
>C�0=��L'cY������Po�S�k0ux�ڲ�0��|L���ta*��s�V������ �����u�0�-f��sC�3J�æ�sb{
�����HO�vY<��K]5��Q�.�/'�5I���i<�]-�;#��,�y�Τ9}]��m�#W�K�ˢ]
J���q�LZ9¿�b���JGn�F1:I`�_�*�8�Ϝ�᥏��1�?�lj��j�v1�S���.�wn����5կ!�)�sp!�g�y�Ip� �q;����9�6�[�ꦞB��?���o��O9wڜ/>�\���_(x��Fe�#jx7��eG�w��I�i]�X�u>�W��yf���A�/y���yI�F�
��f�(}6��d�%GV���	�m��%M#��Z��)+N��lsd����$r�pg������P*��0:�R���
�p��Cv�5�E�DW�ɓFY�$B�;AL��_�hx�85*)D��d��p�q��Z��w(�[l�.�q�ؽ�,�v߮{�4��.-�ZO����&"�%���v2��L�$6|��nHOk{:��@�yL�I�(ͦ��¦$Y�_��)i��lB'�����9܂�Ӣ��cW	2��zy�Z�FNbHQ�}��}�ء�[.�[���O@�~L��x6 ��@��%��4�N���J��L>��MV�ެ_d��s�� @�oY�o�K,��ٙ����n8uKH>M�� o&�sY����3��l�a��~\�A!�e�fEr`�����2^sJ�r��ps��3)�ͧH_Vĩ�j���]��l��\��Mqp����ֵ��>$[�
����=��3� �?C�^kֆ��@b����K�Z(�HJ���m<2�3��XV_I3*��ݢɎ)�z��%QJ�ݽdkX����9��o��N�����a��0��J�|�7�6<��AhM_ؐ��d�q�'��������Eع/����q����+J������L�*4���W���=�٪!���7+z�H���ϧ��TP�/G_��oP�n�(1��({�r�����Pw[S���F~��ȶj�J�L��ӈ�;c�6�)M��A(�ݼ�/�������J�
0��+�)��~��!Ǚ¾��g1����K����Xة�ٮ��A�*d�oj�y<#��E���t,���W�#f�� BD�͑k2mjQ � r�I^un�a�Tyi�����&+�)Q�]fتw㑉TT�)`|<��'�ܲ�6J΍�u�#yG
b)��-��D�^E�t��5Y�a��s9�҉��H<H�+ug�Y����~
ot�&�M��[�q�ܝ���@��LK\�A�-��_yx�UPw�Q(8����S�@,B��������2p�fUW!VZ��`��_LS�Ş�&t��/�z#�!��A!�J�B�g���S~n�4Z!�����{ *��
vaMک)>"��@s>������:$��]��e����Z�*����%����� -G�J��&�q����U�~	�DM8_��-�n������2�d�)R��ʅӴM�H���w�Wo#�*�mL���;aLQx9�	J���x��,r M|����Ź�P��F���>&��\��3�D��Y~����$��Ju7�O��W�T���)Ĥ�u��4�W�1c����>ѝ�QS��Țr�$�����N�����B6�s/w#��y{)=�j�$8˴|7|���506��~�x`��r� ��q�WVk�;TB7g�AL��_����)�^���i�+���FL2��T�闆E���w��&+!%�P�N���
W���:C���0$`O:WW׿~g5m�@X3ڨC�h�?�Ԡ�����4��vc¼���cV9u>��8f2o��h.��k�˒=���`n���\�}ٕ͌������|׵��cO�ϓ��p��x�\e�yZOC���CX�^{M����e7��qi�� ��������[9��ܡ{/ƿ/�����<����ڍH����q������ۈ��ck��q�� *�:\��9�V�@L����4�RO8�,[��CDn����l���P�X5�� ɞ�߼�w��$�@sb�5YAp�\��Jש$�YGdf-Y̯����d)�pf�����<����,(��:C��&"եFF�s�l�&#(`�\\��肰(�WF�7K�����nΜ�le��@b��>^�4���.�y��7C�c��5�bNq���Ԗ��t�H���n�Ul��J��G'97%&��M��29� �1�3�C���c�7"�g�p�	k#����h�!l�)�s�8VԩU�������h2C��yˡ\�w^�c�M�6�b�ƚuSAHඒ��n��vi��=	�x�MUVf��{�Z#,m�a�b�d�pS56�U����	(C�z��ߢ�,!`<���I���9�6I���xӈ�Y�|����10�S�a&$O3ىT�͇���.��;��-�Zga:\� p!ѷ�7B;<����}K�{y��x)���Wwox�Ğ�D���=�@� �,_���/Je�!IC؈?H�^�s34��Rr+/��U�ճ<�ɐm�׫6��X�"������%�9�0F��Z&>��]<B����?�n�%�,9�͹c\�GcI�2��|�8��= E���n�E`2�K���af0o8ؐB�c����UW)��� ����V�ȇ��Y?�VN)�V�I�䞕��awr����nP<�(v���O~�<5#���1�T����ԅ�}Iޱ�cVv�?ٶ���<��;oގh�	yȡ��*��z�v������׉��a�_cN:���?p�;�. ߴ����0�T�2蛏���5�J�<qo%�MM�/�zu&���tk�� A��r7�F7���-p��^�Ȁ��'�x���5��0䱺��"r,#�Q�%�h�^*��^����I�mf�{ˤIύ>D�Xs�Ju7�y�x��R�$#\���m�,�nN��ȴ8����B-
�W������$�=�הV��:?_��Xu_NSP�er��Z�u��Y��7���y"=����?e
2�/��$�f&�cL��Y�<�����@��2���4�P���2ͤ[(sJ$�`�=f����1^c��4����|�����j b*�nk6��\!��<��`9���xSʤ>Q�,�~�G�_;w$����P�A4������x 3+B۞ ��L�I�x��?[<��n���C�m�
����-���C���ԜC���u�,�@b፹Ҵ�g:���#��;�v�y�y_|i��� >mg�-O5�Yt��P���s�	�!Q�����i�sv�G��7��wO߸|�.؆Yk��C=_�o����%��&P�������5m�o��q+���g�r�у��p��,�C��3C����\ӗ�w�Y�U9�ko�����zgG��d�C�J9Ò]�3�+p�B�b�>�����9��-3!UJ�ajf[�ek���[j��v_c.�~au]=��G:�Ic��za�Ajd����g�6%�.hDj��&]-�cO"@Ƹ��L��c��24�|S<�M�+����h�����-���a�2:iI!���ի &�	���gFF}{�����DQ��\��:PW���2���盇���	�@.>�0���h�x.�ænUj�����_Cg�#�|`��4`��w�1S�?1�L+��o:k��糣�����wɡu��紧ҽ<m� O�,�5�G�p<�q��ُ�7*_�u�E�4K�j?�|�������F�r������n�Ƹ�N&��T)��Xe��R��ʧ�����(v��kyE���m�!U�)���s�)��|�����m���� ���,_iѕ�XN2���[)��Fl駛�^��GG�d��G�Zlzz�~�?:���*["��P��;�TC�!U����;{�?�p+s�
��ݿ[��c[�J�)6|@OϺ����#���<r���{����U���C����E��O�;T20X�Q�v���f��D�p�r�Ֆ��aF5DJ�
�_V���,�C.����W���㻔N�!A�m%��g��|����1BTͽ��Z��f�z|䪼v�z�+0�\s�b"��ݥK�Bk��">�VL���(�D	�d��sO��f�
CHz	��oY;9���0�ߓ��XKG��87�w��"^�#<)��F�
m7�̰ћ'��N< W��eڕʗH����S�������ы��v<�VvF��(n����xhi�9��T�@�-�|�N�{M|
��R�b/�c�wQ��D=٨���8�E�f�����{Ș�x�.��[g��� ��(����׵J��4��u;�H輴�1�Fϣ�f_�q$�S���b�������ӏ4f�:F�t�~D��R+�zgj ���xe�{d,�fÑ���bo�5����Y<��X!q�l��h�$��n}�Y{�A.�t#��z- jm��Y�m�}X�dԭ�R��C��)��X�]o��b7����Pw~�ѰLeNS����4�lg;�|��GŪא^
�}�B���I��������Jϧ���#�Jl5�����\g��6e�N�x�+۲0^�W\��6�l^��#�"9���RBQEa\rs���=`�U��x/�J6���*�=�'B�dDw��B�T����X�`L��P�������=P�_��\-� #�Umom�d��0_�����Z�C��M"��_z����ӡq?��2�� �kb�C"3_e�b����߭%R"UK�Yh�MN��)�D�`�O	ס�h�6"^�?�d�Q�~�x�A&{�I�{�m��rc��^��z��[�|�N����b�;��VB��2N�cm��w�����xgS���[X�_%�/�d)�)���иpyHG6N6?R7�`�/��5FSg;�E��L �pҼ����+
`�e�3{��_ꕺF_A�;5�W�
�h�&�,bQ�(l�+�LW�������u�?�I�"�ՙgT��q�eZ���Aj�&Z{�8�-:b!�~}f3�՛]
,��A��R!�ր��Jý��'rj��XR$N������d&7d)�Y��C\4@<
�	��<��%/�"8�dϠ�aA�����!*�O�7)3��:1��uDZ����S�ݼ���2����`:O�g�FX(�a��/��	��̆���������ԅbB�Kǣ�Z[3��u������B�g����Ě~��� cΛ�>Mc'X [�ue���!u<or��V��b�i�]t��^3G,jɵ��EmN��>(���_ gɣ?�}��z$3G7r�]�x�IC���j;#�M��I�/�u^G2���| ��J����ѱ0%�*�Q��d͎b�3��O`T���VnS�𤌼v~�-����l�K���H޳MxV�hQi6S=��cx��!��''-����G�&~ʭ�!�ڙ��χ�r·�3��cy��xJ3	̍Mq�R���fr^wf�V������ �qL���a�]L-��67#��ĉ�>�{��k�y-m
�l(�5��B��2�N����ӿ�p�3���
��;6#4�br�����0����!��`,�b��Y�6�+�4��焧�\���^g[Qwx|I�:�~,�|�Ll����ɏ]���ʝ6�?��p�qOɁ��C&_^�7�����ŐV�˾���T�
�W�p�������ܠ��,f�"T4���荪�SV���޸$�¹�c"�:3ǃ�DD��[l܍��H��87�WҊ�D~��3ql���I�×�@+���҈���a@C��ţ^��c�vN\�X�:�%(� ۧ�9��F:⯨���%��Ztl�y��5�k��7�(������%flR=��,�e��=I�a���3i����o��Ʌ�UK��Xi����=�N�ʏ�s�j����2�L]6�Q.
���Ԯ�&	Դˋ$�����CJJ,��&_@}[�I�[���!�������W����/:i$XK�MǾ	'�J���g"���#�|�w���5_�A�q8�ߘG.����H�Ej��n,��?�9ij�ꨡ�o�7�<"@����p�K���̌&`����׿��oM���8&ӅRt	Z}��!N9�-��`��J�Gͱ�����!m����;2�f���=���∕�ZC��uѯ�6:�������S�� ��§֧����u����`F�߫���6��ZLNW�%_�k�	�w��=�/Q�w��
��@�0�=e���Ypd��z}I��0�rsk��m��-��F�э΅�NG��^
�����q��_z�6V�E����/n�ƻ��38�W�~(����픝:����p�;������d� r��!��5�,�i�ө�$!#0qߚ��<��	�H^ӿ�fAG?��
<X\Ɖq̓cr'^�0�?|��ASv	�w)o(JtI$i�i��>�/�k)'?}�z�΋�u�u��wMZ�	�j�\�O���>F�M�r���-�v!�c����2=]؉������"N��\��zEݏ�/kW���΄���t��Z�lg|Eb�����VY��)0� \w�7�*���b�X�D���άc�0k�H��{G�biNW��-���k��N+��o3ߖ���b	���7a|׻��Q��k����nM�H�N�
��S�8��&���0��)�ɭ�T��]57��	�y�U==F��E�!ݢ&@��#.ʆnHik�b��a׷�s�w�b#��:�U?�� ��2�}���x�1PV"�=N�++�i��n�oIB�%���0�u�Yj��Z*�8�8b��Y��K.��<���2[��.�������S�T���w�y���KT]���M�y��S��D���10E|�qF�,��׵�I�
�c��_�: ]�ז?1�t"�D��4V��	���XS:��[\�Zדv+�_��6r�r��������ts
 G�Igj��k�ܲ��vD�p�z��Z���ީ��	�K& �y�$�"�nQB�� J�D��f,4v��������=:�^� ��&!��T6K��6�
�?Ժc��>��G(�ア�������=�L4%J'�V�����ca����>�6��xv�&䋡�-�^A*R���dE7i:D����x�)�(Cb���x��׻-��>Rl�O�ܐ��~$�s��	V*Do]RV��n��$�nà�����vc��,�V���yִ�Bv7ǅ�@�r?��y�uَs�;�W16��ݑ!~��M���t��Y��T��J�o@��0�쟏k�\j9������:h�������xY6�s(��}��`p+XY�xL|ɝ���Gr��>^6׭.-KV��*L�=��>�e��kf��R��J�a
�"��=Suoq�>�8�d���]���W��[�3�\��/X\�,+g�.O�V<z�l�B�D3>�+�R��xf��DO���n��%V�Є�D�/\�)N�#y�}��(�r!K���}�=�ϲB<�p��#wv�1V4�+�5�������;5!�9T��s���K\:��u�8�8��ǣ��-�f��C,j�d�m�`s��4m|��,$��x#��*�[/���2���¦jRV�p�����&d���}u�D���J��$�9=Z�0�{�ض1�4�N���#�.>#��& ���dg�`m�F�9X��?сs�#�CPC�R�����W�)��"��q*�ӭ�֟��>�A��G`H��"���~��&m���x�'>El�*�y��ѩH"����ve�E�
�U�hN�h*A�_�S���$����g@�X�6�3!y}��B4��շk���s��/�VR���W����/*/��a��B셮�9�6)�n�h���F�_�U�ǟ�-jM���U�5���
��a�^Q&��A�n��.,.U�"|�I���OD�pc�r#Qs<��[]I�g��'
b�[Azk�^-}pY��"�FVk+�,q�ءN����d;G��'����RP�/bR��x�u��1C���o�O��?�8�-#�Cd2�
������i�8}M���Ќ	��z�Er˜��	�y�lp��{2
���big⠩T�ܼ0�ُ�^�����M�m&=�3Z�і��yݪ+�-��"d;���w�A�ѻ�h��������4��oj�f�+{�n�/9�������\�|<�A��[=��M�J�ݥ�
��#P\~��5MSG�+_��a�̉O���K�g`����4��K��b������	8j��kg*l��3'�hkD�l-�k���S�<c�Ey.6[В�~������1B����c+�ekU+rU$����l3�<4kV��n�<��j���r
X��h��^�4�f �̳�^\a�f^$�h���|�j/xhh@�J������ܸ�<�Bn�m:�״O���>�o�5Yi�9��ܺ���1�!�|(֬|H����F-?�8�ܹ��-QRn��Ń��	w��@[�!����М*f&���ΦN+?������DZ��v�[���P�����!wB����P3I�]�Y��n��6]�}�0�����4c�zx��$�5���߮Xy���3��AX�gN&�mɌ�_�x�����
�WI��� ������w[�p���+nM~��K�W�i��(�3?l᫢
�k�4

鸁.��$o�W�z���a�^����j�k>*�%/�2����T�u�l|/�UpH�v�X�,�mpdW���\b/	,O���	&�j,{Vm���(:L�dh�ȳd��eE�)�ڻ��MlV�7ѭ�6�W1�w�ʪ��f�Պ{۹�NOѐT��l�����q��L}!P�&�쐃����z��5߱]��Ge5�6���.2TMx'��R���^T!��ut�[�C�`�Mz<7�7?��)��ԲڹuI|�vJp��[f��b���B��7�ց�u d�l�Ə/��|?�V�;C�5h�0���,��VP|ᾍ��2t<��@���d��HTZ�J�����M��)qMء�X��֦_M"9���(�d:�~�t����hÜ0��Q�y� ޸�I����r�$�4��F�(��M@��*�R��r�(o��W$��9Nv@�)Ăc5[kA��2p�c=�X�/�!�/���*U?��Uښ�C��r� l��H;t�zb���e˯�B���ʨ+lQ=%^&����;�,;��M�<I_̻#+�B����v�*m�u��_��9K=��d]�O���$���-��>���߅U^�S%�ye8=��"��
f��8�l�E���Gџ2��hÒ5�Ͷ����R����9P?V������޸��������l$������	U�TϹ��]
��o��䎰.g�)���	�n�]�Н�ҭ^)y���be57�/��[ـ�������E�;��"��#��"l��
�R�A1�d���x��O j`_�2<����8�M�+��;���z홺��i^',�,s%���Gi~֚���EJ�Y��_Д�6����Tg
�"��a��լ�n�ۊ(����u�9��Gnq 1���F�#+�<�O=�c��(]��d�W�o)���̋�[(�T��a	�:��c���@�����e��/e*B����?���J��F��s�G�-�NE0�Ï8�\���E[�/��"���A��l����˄�#�ig���2��\�a��ߦI@�Ľ� Ҹ r�i�|�ѝ�z�b�UDi.]w{����	i�ܕ
/rʔ&U �?�Y1y�]�*��)���}�6A��	�l����źe!��+٪��+�U��`j����;���u���-�w+�/��VV���3�Q��|u[ vC:)� ��Š�A���<���aP��r"����G5��C��f�������J�hi
2G<�.j��Cװױ��<[��;8i}�H�����X�\�D� ���� ����tw��)�'�A�J�N�Ƽ�v[�&v���jF�z�J����:4�B�v���3��
��� �n�ɝ �9���-C+s��;zsǾ%�+(D_E�vZ���7�N�Ϻ��R����
��ךE�Mvӊ�j���@p{�_Z�%�9t�	���/�/���&�y���K��`n+�ì��F��b��'xKblv�����x��e�O[i�f	���#m���d&��[�	"m{&T �D���i�t��X��T;��B������M�PU����J,�?I_t��<�M����L8����7��i��&��\`>"wb�I���s��J,����D�z�k��t��9��&��Ob<�p31�.���|�6�ԸȒR����]��k�u�`-h�*oIS>kS��ڂ:�����T,�Bv1�H8q.*�Cs�7�i���Z^X��ҏ�e.��蒷���e&���3XeG���rQS�=(����_��4�\��`�@�h�oӲT�4��R<�^�4G&���� 
3F`�tg�˜P�'���B >�/��A�R啾 ����r)�	�/?V��F��myn���(������x�w?(u���J�A~����F\��e5�s�g�=8O"F���N����u�瞑m$̫w4U&���c��W!j�0�m`1�euZ�y#6��c+_R~\}ZL�ץ��yJ0�J���:�󨒦nF_�N��G!��5��zd����J�"��N�'R�|�ƞU�k�D���]es��m�^�]�=�Y1�Z���8�27uu(�>��B�+�6Q�rԆ|@$��Y5}=��l���=]W���V<��(�	��!�:p{2��>d���c�'�&i���|Չ~�6<{�΃�L�)��:��?�P��\�n���q5I^:H�����!��b|���lFJ*��u��S��|�zm�I�1�D�
tߦ�O9����Let|�>eOIO�5��_�}�3I.s��(Y�lG]9�����[[d
w���f6Ϭ���EϏ�bl�p�T�Ϸ!����QA���.{�w~��D�b�n�JO�W�9W�_-j���%�h��0(�pn#+�oi�V-�%�a4+�z��������M��;l�W7iE������[�(�Q�#��Ϲ9UV��wu\�3�Rʸ�C����k����B��Q�u����}��q�([*zT����5�B	��@8�2�r�2��B�&_�k,�Î�`A�������k�\r>�_#�-��z䀗+�!$�����F2OG����*�7�ť`��=:�ٕȫg*}e�fM��{X8ye���<W���j-��xaV�������-��S/���YJ�^���7����b��y3'=�\�7@�*7�1�*}d�@J�F,%��s�'�0���Y���.
Bm���-�i(��++3H��6,\�3ɽ�֏bȳ01�0�\T�ղ`�=+�M #�mJ�^�Ŭ,~
��C/�j�w	�Oo�
��~�Rlc��Jt����(���<�$��s�w��n�N�Sݜ���j��6�xF�-@n�t��!�b�7k�t��]`�P2�ʅ��B
1a�Rq�����aT�ӳ�f����6�k�>:*Y��
�i(]�5���'T��﵂��F0���S��Q�O����o�m�����x0�C���]`��n$�ϒ�
���n^
q2��D@�����7p��]s-����כ�&��nH�q ���7}�K�j��^��؎G����`b��n�=�tdN7z)S�$�b��[��q����a�<���´jB���=�Q�<� ;����Tf@o�'�M3����$�9���X;�I��̖i��[�ņ�+�p�� x����.��T�8VJ��n+������ɣ����4c*�"���ܻB2�G��%KU�����vpBp�I�C�@��Ҕ;�� hϔo����P���汤 Z�e%l�<F
y7�Q;��R!��i��u��]W���{��x����% Q�іdq�l�1�����
~���]�}�^h/&�9?��JM $�
g��5���D6U%���n,�VQ�VkO��R
�½����9�B��%E�w_���c���lUY+حUho�+�����ǯ߬�'�r�O�uEU��^�����V�4�1H�yntnu�)��N�g�Hn��\x5*�E�B��Ɏ���3��m�z���c�P����DZ�x�t�|��N� Ό��ӦqJ���b:�b�;2͙d�����擕����/ݤk�Q(�`%�
a:�j�u�m �����X�~bU�O�HZ�5�r[��CU�t1�fbiz��mA��O����/u�#��MՈ����.K��dޓƖƦ�)i�ݕ�o�A�U��75��iJ�!�ig9�����SM��K�r<�q(��	�[���x֯#��٣����t�����-���xv���V��z�7���ܑ��]4�E�B�Pr�C�#�_<iS*�h���Ȟ��}�ze�p$�uKE!�J��Y��@��׹I�%P<�륜�p4g�狇RP�ܾ�1qmB�t�����$UE熢&xgL����D�7�c�������+S.�R���D~T��bL��t�0�G�M4s� j^'�}y��w�����ھ�c��҂^p8��>zj�n���W3�e{TU"r8�[h�h�o��Ϗ&SQ�N�4�띱vd�i]I��ʩk��!�;/ì�E׹��q�<@M�ቍ����hX� iTهŀᓴ<���xh_�!/�mR��S�99lĎv�r�g��2����x'-����X Ǘ}����5OW�o��x돕��G�*�H���^.|���3`���Ԡ�G���AgR:K7,�w���e���W��B��M�ǜ̃_G(��/�;��/f��l��L'�nx�)i�{�W|�Rp%]]�UA&�rxF'�6�L�V8�(�0�E 0�ßc3+�:དྷ hi�����5��!g]����5��˕`��o8�����g;��CM�������%NU���]��~p��4����r
�yn�H	"��l1��sN�t�F�dz��.�����^ee�ν��	 ���<�6�ID�O=�O��<���s��,{/��H�q��|<�W8�Vю�H�`D�ö�r�8@M�8ɗd� �Ws��|B�f�V�I�cq�y��Y���8�.�st�ْ��7��%[a���f,l��c����|e!)���͌bw�f�oo�

�'GG���лV�������-&R��=
�֠. �2�-*Gg�pD��G�FY�^¡~���a!�b�nN��g��	���9#�p��-"1��_�Ġ�0����[B+5���l� [n@v��O��uw^:�~��	�@�T<��:�j��A�����ÇX"��g]���#�����!!��������[���xC��OE������*S�jb�����A[��4��G�q2�[�>���!�#���~+�P� �iY&p�@��-����KD��6Kӯy���"��	��qj��:To�?vq�|�D\Z��&vdP^�TU��h�Dk�S��'��@m#UZ�Ȏ�j$�0��(�,��x�~Y=�CF�A���S�u�������7�ޡ��LBq����Ā��BG+F�8��o��s�'Q�@�!�m��}d%\E��f~xWn�������GR�`Z�a0��
���z����h=�"�_|^j:k�lC�����D���^F�]�֓���L���o#����+5-���s���3	*��vxOZ%lK���j�B+PK�����]\��\�sx����#N|��c�;���yԜ�~ToYC�t4���+�G�㸄U��2s���Q$�}8�d��?.��C�$�"q�V�7m�?�)����	�F���	Y.�5��x��ZB��??��<��ZX(��CX7�s9^s�"�r�r:���K0�ԟ5���]X�﷽+X��`���ʧ�8<Z����}�/T�l]�U�4A7�ѱB�H.j�T�K���͈�v�:�#/���1~��ƶ��B�`Y��Wl�u@I:�¸�R	���4��Q� N�^��V�v�N�C��P�*vH�(Z��s&���<�3���!#�_�sr�cOP镥2���̕�eu)��l��0СZϼ�9t:�R'�x�� ˧���8n�q��-+� Pw�V�8e*���-FԪ��v^���{�<�UÎ���>@�1�0.��e�e]þ�=���`��u�I�J�h;����h�e�^Rw�[��^oN<���hx5Ԫ�B\��A<	�^ѿ4R���U��iS���`ӱ�����8�M���M?{:�g�*�r#�҅�x΍��=jG Np6�LxJf�P�.jW�w�M�wu�i[�,~W�҆���������f@q����/�è?�����P�+�gr�d,�bd[:����&�����XF�;�:u�T鯧a�2[�?Uh��8i���cQn荕��u���<���=�[|g_m�5�"��6���l��y��nZ$c�U�$����VZ~_7�a�F��ArF�4LA�Z3)��؁5}�� -��zAO�4�
�A2�:
�����N��n3�*A�."���)��Q�c��O�xF��s�g�(5��$���3��>�Ͳ�Sq���g��n�M��7%�;�,�s>�&YTq�N�A�T�Y���/9��0���G��N�T�P�����rZ����8>��J--,� ��B��İ�h���������b�Hw�+�B���"�b���,��kە	{�D��	��Q��T�@m����u {q�[�g �׼-\$P�]�����N�e� ��?��W�L��}�>(������\�vq�%.��q	�:D����y����ܛ���kн��ϲ�j�zA��{iV��w�[��T�`���&���4*: ��)�qI$>ץ)���tJg�q0�6K_�;�>8��a�'I�>w�@�M���o��}����̽��N�w+���+���c�M���ֱ:��3�	����5�Q��W��!���_w8�Z�d��[�	;g�v�I�!��hs[�eUz�$�={��E`#���}Q�CB�������v̗GT�4��k����M)�d�0���S�̱p��-K��e�.�F5?Cq�5E6ԉW����z��r��:�*m*��_h<�����^�0��o��.�l���;�̭�ד[�/���d7��R��"ͦℱL~�}���9���3Kz�Q?� �+`�f�);���r5*��@�y�i���W���i�Y�s]ww�N���TX+kL�	D�EN��SnZ��X�i� $m���Ix�{U�UfmPz��MD�b������Ԍ$ዢ�/���3̀\�
��8��D��.��K�j��������ߣx��?�K�fe������;��E!`}�~��P�;��+6�P��RH�9�����({yn@�{R8�Yӈ���ڃ!@3ڤ�nq$�kz7�y��a ��v�YGP�b����%g[��m\C�m(� t���nm�*9{�9�ӍdV\�#d]�Z�T ���g;c l�G4Y�G����������X˃w
�?���+�!s*i�(׺�����I1��X�=�!�Q�kF�zŝN>���c������A��4p�:Va�����/+��b��݊��Ru��۾��|Z�*�)�	�A�����҂o�b!>�NŞ�E($�!d!�e�Fw�WG�D����0��WW/~���u�Y����*�!%��H�d�:��Y"��0��Zx�4�ѧD6�q��n�1(G�����?�c�ĉF_"���L��)oG�������ge���k�߿�P�{,� 	�MK���r�3����Q��߭�5~ I�$�"�V��$�ςi]�`�9�mj5���xL�w~��@�֧|�n&�;��� �U*��A�(�x��;�O�Mu���2�1�n��J}l��-t�7��y�5	q��H[�v�n��;�h\��&�2g*��I��b�ӱq�4��^��� Up��m�zf���Ν��BZ(���c���{��}��O��*�鼘Ѿ���9�����]\���޹=͵*����-��ƥS��]9��,	� ����@IpJ�K�����>y@4�>t�"DeV��&k��ҧ|\�"=�$nQ<ʓ�o3�"M R@���܏P ߔw�gb(��kW�d��L��t�	M=О'�5@2ߺW(R�lX�x��se|u�+p��Ń��>��a���aB����a�v����q�a4u&���C�}�����	
�1P���x�~z��`���n^dK&q��ccVDop���H�4�����6�#˰uͬ-M��9�i͚��U��N���P�؅���¯6� ���|�r4o����4���>@ �۴�hf��N�yI��>���ɓt��U#��������9��K�~�kFY;���6X�U�?,�'���5Vc�
���-#�W�<c�r��?�U�����3�rŇ=y%�d��,H���2�Uj[6�Xr;9�s���	�O�:2��9m� ���5����Ix�)2��iہ>6�����L������ҙ��.~�
^2�d�����2���|�� ne=�&"��Y��$�}!Ų�c+�@SNg�������H8u�F��[��=��FTS@�W'�X9�#����rY u�ۄkm�\��<���YvJ��rkݲ�!���4���d��w�	ަ��\4�!�F~��;z� �����������њ�J���a�x��T�+
�6�*E}<��O(�R0O����u�/�{��ȅ�_��9��a�r,����{��=�{�o#C��N'o��{ғwݓ�>���:4��~vU�Z+)��襅J�����ʶ��iяc�j�<�^�%$C��/b?JM�:Z��}����Rk���}�r�]dR�h�By"��p���$0�`�P�ϭ'��Ջ!E1hv�3wO�����9h�ve*�M��b��S���o��T!�E��Th8���3͌��/}~Q 5S��3Z�} �	��)M_L�RF��;�� A�E%rU_���}��򅵆%�/;���^�5�dg����D5��� ���#6Ī��ݟ"Y�N��Kd�<�_HLw~��]$fP��"R���G�in�a,J]֩�#��0rh�E]7p(_c�����N܌�s̻_p
z0��q���wYY�<�Ih�n�х�w�7�|�\77n�!;��NW0Ƈ�^i�c"���mĤ��L�l���}B5~
<�[$Fp�+΅���M���/��]����y;��b#��t�����m���%�b��5�ا-GhG2h{�̠9\R�Nۇ<b|�,y�K�i��/P#�6�=��p[gv�W@��|\S��ƦYgހ"B�d[��cN֪,t7A��_��g6��&=�.<ݨ\�37��$24�u{Zާ\#���ץ���Ѡe�\��u��������1��2�����Gh�g4-:a���f�i_���?�о,�"�ָ���N�ө:@�O�E"��az�_���_ C.yKcH{����!��n�8G$�XF	��E�l������g��r�	:�-?<u��q���NE�WԏD T�Bb�%�Ks��/���"��8��Xy������^yod���ǯ����S��\j�O�V��_�j���
/��l�nB��b��ڲו%~�8��aqI��,�K�v�ݸ�ѣ�il�?>�j�A.l�%,Kϐ3ɲ܇�j�����kMJ���	�����
fq�ǉq����Ŵ���m�����K�u��8]G~o�FɪmKX�}��47m8�����[��F|�g�Σa`S�ҧ|�u1���}a3ޢ	Jޑ-$���(*��DG������DE�����{J��;Ƃ�,����M��^d7���.�qz
�k�/e�>�wuX��'=Ġ����k@��s?F�T����/L�s��{g�A8����X@�g)"�x�J�U���� @�����S�ש�t��m�p����x-b"�(>j�ϫ�Lr^��CQ�<B<E����la�
W��F�hW6�x�8�z�Yθ%'��z�3�(6�v�j����I��F[��Z��{�m�?#)ƺ��">q?D���sB�
'ü�^k �%q�J���g�tO���JIH�$����^n��Zs9���W��z�۔�gL�qc~��f���?���Sb炈W���`�4o���9�ٵ�d͗G���w����q	ʫ�~y3�IZIN�ub�&�Ъ��7X80���ω�~���(�"�'���A�į"�������jɶI,�Az:o�	�QЙ�x�D;�s}O���ʋ���Q�k{��ǈkG�
fs/¬ȿn��h=_�i�5@ί��+�
���Y���sY�@�)P��s[r��j8�˱�&5�c;eB���L1oK�e����z�'8e�.1�4L��}8.F�}i70� K��;�%�lͨ�s�+���?S�"��ɾ$4,̠��z��u�n�{�3W���JQ+>����3��H�a9|�A�알(�F�d#2�x���@��x�F�4���Lѵjw����Ǣ�j���,�~=���
RL�,��h���#�Iǯ4��uxP�\����R*[6B�lZw��	;�B;���Tt��^
I[�Rk���rj+�.d2�7^�J�E��j�L�E����m�f�0fpN�^iQk�8��N�\���z��h�Zn�2r\��Zf��x�(��LR[��hM��ΎBm�Q�3e��o	��C��[q'܏��&f���j�gc�Qw�ا
���l�VA���h���?�:#��<��b�e�k�ϧJE<����ʩ �8F�*��dSP��aPO�;�-�>ѯ�}���H���a��¨����*�X~%C
��<�@�՜K'�몹H�����l>�)=�{$%�gV��)�v"{CM��5���*l�q������Q�m��zTOr�'���h��8K�jX��(�ڱ�U�u���"I��� ��@�IU�%P��xG�/��a@��iZקl�*nAj��YIR�M{O����P�C����|&�j��ˏn;s"S7�gc�Vy-�4v�Y�I�V�:ջi�-�0?�-�����s�������Y����,N�oj��j�%Ru��E��ޓ��6�<�BQwe_퀐(`��3eu�+�����7���w�n"Un���\Qb.2I�Y���E�W��R�3�g�b�x�;;ݱ��8G׏�`�Л���{޺VD^�g��Z�}�'!j�5�|K�PK��[�\����v�.�M���bg�fhX�]Ja�� �-��% ��5��l�/�����ܼ8M~J�Ȳ�`y�qNlu�Fϩ����m36Ft6O
�+!r�'c�8O�X"L����S���!�&�{v5��lO������k.g+��֚��d�����?�.ֺ��٢8_�Z/l#�z[��_D 2������jz��x�;�q�(b�I��`��Ƈ�b�l׵���tjM�]��_Z��;��G�2�*�=���p�
�hSoS��N�]���%.R�vN�TAI�q�{H�ڭF:����S�V��w3y�G�fth��/���#�]l%�*�%�������eu�tU:�}�:��U���4zn$󌍸8��C��6�����B���5����4W# �31״�o#-Td	�y�mM�=	�նs���M�ѳ��2��p�Lm�lQԸ�1�Qތ�_¢�M��b�^���Y��rK A��dr/�|�]�|�Cl�N��hK�i�f��x�X[1��
ܠ���0�@H����AVNoNnȓA�U@P�;���.�>?FX��"y���	g$ש	\���C�z���؝}8G�o"pGP��W9��z�7 5�ۮPH�����J#,|�H'ͧ�*�,�o?��V�D�9(���f��8����0+�-��nAǸ={�'6������S}�
����`V�e_�!�3@��"�SW��ɽ͸�5�j���c�4�K�^3��S`7��8��4mW^�l�;7"���$DT{o3�ʷ��9y��X���#�Z�aԣ�7cH�	���Q�s\zmVj���/T[w0�������Wf;�ةɴ�$�#�"�6&rE�o�l��\��8F~����졋��y��C���ä܏f��(�"k�=��^�C+Dc��Wqє���S4�g�/�X�j��h]ˤ��}@��zO�z\�(��@$_}	�����8BqH�h����fL�-�#�瞿�tM8m�${�?j��M�7R�HE�DU�;��7��:"%�*��am�*O߫�D��6ܾa2�����u��/�֎���l�J/��͐MYgI�����M��u�*`���S�!����W���g���a��e��p����$�Z��]�IES8C�ۖ�y�t�^�װK1���q�Oyb�Cxeh�LE>�g_Pjj!����H�����P���#�.8�B������Z��N���iP�'�1�u�����h�"۬��P(�ᷲ��:�$|���6I��Ur �[s-��U|Z|������ZJFݳ��I��b��l�`[��]�\ƿ��_��4��>�n8l�{&�֋�&oԇ0	[xH��.��=d]1�#�@�B�N\�O"DGV��xﳲ�珔�V�v���b+.�sA�Y�l�0�f(L%�:�,�W�ϓj�~�0ؠ�'���Dۧ^�
)������	�t�p�׮�c;��/�5�O]�K#�D'����0��0�J8�dEiRnrm�L'�^V<k���{�F����c��~gI�M6E�#�z�Q�g����� �m�˶ȕ�"�qKe�9]�o$m�����C��v �GLi6}����u����ㆠ��K%W�ub��Ejt+�.o��B,q0ע,M�ބf��0�̾�&��&e=��}���lv�y���o+� �J�[ʣ��0�_ծ���6�.�L����$���V��j��%?�#|I�9b�Ҹk_j"��*���*�/�T9�Z7���]����+��r���n٥��]�����x U"@�l|���D�F��G�����JP�� �[Bgl
#��q���<z̆��^�x0!���1�	Y���4���I���(c|;��@tJȈ~��W����9ꖂ��&)_撤���;��m�\���S�.;���Jɸ	�����[U��uea�q(Nq�U�0w���eXqv��ߔ�0�ݧ���� � WV1�u�ӵ5�^�.y�Ե����1� p�_� �"�ظ�]�&�r���(�7|�q�V��o�d�'��$�(�چɹ���D�qq]d1���� �y��;�j���gŦ�6#U^w&����MQt��/p,��Q��*Dz���uN���ӝs|�T$��`�����QM���N���s�IW��VH��t��H�=�;&�K�S�.Am�2�BZ�Yds������c��&��mQ���N~�(ߞ�'>g�1��}��}m>I8�#�Aѳ��&|H򴝮���a3?[�j};J��ﺱ��J�&!0∆��������Tc��
 }s���N|�8fD�M[N�,n�H�$+[}m<��<af�����.�d��%�>�v�ϓ`2\�$q�م�v��{�W5�;��}��e��Z��f��n�6��/\�>�-�ͻ�޸S>=d~M�_a�|����cӦW\�Gsi����x�1S@�9��"�N$z�B���o?����׾;^�7/�'V`1.4��t 5ao�oA�Y�(�t}���q�`$������H���j����%u���V ��t��1
W��jc9�B��&�b�Fw;`J��i�Q^��څE:p�Ԅ��C�O}iF5��ã�u9�m;��%W�T�6�tV��}��0�V�xa��3;������,�������BLz0� �뤕zө��&���#�C��6f,����7x�<�'YQ��D��ʿ���S���vPf�k5f��m�nu��P��R�b��pR��TnM��l�uU���
�D`ʣD�^���鲵G�"�N�D�ĳFI�Pձ���lڒ�?�b����U��x_����a`S��B?qo@L�j֔�V����W���$����|��P1F"5����D�b��i��STb$h�qO:��l~#�]�e�#�-�O}�ΨA�C}�zX��P�#��F0 ~0A�S����+r�e�/Ǖ_�&��s�i��}W�9o���݉��Y�R|X�W�S<�m�cS��Z�{���r�(*�(.�&��R�B��pjQ�@.^�' k��r��
�����xT�j
>SjFaZ=����I	�ŕ�� G�#���_-h=F�j*�9H-� Q5��Zla�u��7��b|"K�w�y��-y�a95na�\���}�Fgm��n�����s ���O��{�ҽ�ɾb4�]��Q����U2`UX�M�]T9��w˘I503�/Ix�7vL���O�Ǿ�r,���*�pEG��&*�����kjq��U�����m��`��Ԝ(�?�"0�S��c��}���B"�Mk�s>�E�Q4c�l�F�/�N��Maeг��DG���^��o�^2 �t_�сj� �3�+����ڝ�g�F�D¶�(���1��G�ꍒ�W�U �Ew>%d���@0��`��kK�َ5�Сӡ=���Sz��Ԧ',�R���敭��&5I��}I$b�HՅ]R��� �x�}��8� /��t���^�eN˒W�*��$|��2�!��AUR��?�T����	��sP�t�(j_`a�	�^ƣPkTx�;��Ê.P���z��E)�{��SL�?
l��v�?�/�����m���is>�jilF�_S�D��v�Qz�6՚������������C$>��L^��(�+2�(P��J�p��2�[b�S��℁���T�&�(47�;~ҳ��A�Nl��lm+�k�MVb���df�.*/N�^e���w��~� P�����eF ��%_i��f�P��f+0aQ8�� Zڡ�k�q����0~'$	WW4(_=��/Y�����Ҧ^����'Q}�?=��zi4�c��g���o��;תiZ�a���/T��"q�d���ݯ��F�_��7�e M��w{>�¸�v�LM����j�N˷���	Z������cY*= �n<.�a�|-�`Oq�\ӫpF�_�N��ƃ��M!+����η�)T��ߠ%Z��tX�x�2�Rk;�H�u��޾��Zl2�o�c:��c����` 1��l���o��9p�y���
�|�囗�ThgХ��8��^��9V�I��tOl���/�(i"�<��}�z��Yt����H'v������+|�n�!ݹ,����~*JWB�ji�]	�����H��<�Z:�w�^������{�V�.;��["�$>*^���<N�s���8��b�w-�1�?x2�&�P%�.^�"�qeҚ��as�f;�m��&���g4"#n���N�%�!::�p���rksZTn��n}<�(r��4�by\Ny�u�*|�IU��8�&���.�*Ҋ\B��VC�-VU+�xZB@�_kN�.N:A��u�rRK�%C�� '26��k?B�f�B�Y|lߒO���n�PJ�E�����&�˴�/`��������M	��G&�L�jܨ�/En�tC$#��<���LWY3es���������h�E����fܰ6���^�m��\qqc� �x�w����6pԄ��e�$�:U�l����[�J<��5��Ɂ.	K�o�{`�"�Ta��������g�Rox�U$)��է#���8�49�ĳ$��O�7Y]�.�|����3�F�$����ZǑ���𞹳�f;u��������u�Rb���Eqc�HOnD�����Xfo��a�/hBJڵa`h�Tn����_�o�[�"�}�u���l)�z�°rQY�� �E?GN��W<E
��������,��k�E�<,��f�*�mnQ��J� x��s�����\!I�h�F��!�M[6��͋S�����0�gRm*9�s����>��O��1��GY~R�4N���r+��uu,���ފ�3C�0�=���(M�6����/�{!�����q�ի�AϷ'�a0՘`N)_S����Or��6����<����,�qeY�;d*=�r�Ǐ��D��
��%����S@�\n����r�\����e{`���>,/�@��Q������*t�v�}�/��=��1�As�\4��J�Є��=
% ����k���
�Z��\�M@޽��a�ix�9%0��<����S^
ª\���j�kc���w��{8X�o�1��#h�E=6]i=�T�s]$���|r$�CӖ�U�y�>|�>��)V�X�g�{
�P,�k�aS�ƛ%lg���\��L5`ca�zҩ��ݥ�RQ��m2��nY)t>�Q4�y"�٬�""�OU Hk��Fzي ��?̙V_=�R>�/�n�ףZY���_��۝1�^դ�_$���Hk�ƪ{gGr+!���L�����F`���^��� ���7��T�{��W#���L���*�1���)](��U��h���l����(���淋1t�Y���Z������k�9�s��]��}ǩ.���mp8OH�@#oQ�EC<���z)�O�i;nU�B؀��S��xG��I�c���k'��^1��XxS���H?r�Qi�W:�c����7.����LI�n^&4*����Ad�wڻ|(�̋P�����x/պA�?�H?��If����4��W\����[;,ܙ��=ഌC�!xF�F��fׯU9q��P�h�'���5dȞzJ��=�.�D;�g~��\穵d�I���~u,�R�. �S>��	lL����WZ��$��mp�*:��&ۍ� ��;�J��_�Wܭ��R��4��� �`C�	|dy�v=]�f��h
�W��|pZ����@ݙ��e���vi(��"N���x�W��isp�'��!�7��;��I��}���P�M�U�_�$$Ђ�n�Ód��A�s*/���vZC	��<��p�-����l�1V�Y�󽪌�B��@N�����z�oz��td+. 6<I�S>�fԭ���t����n�4I��7H ���L�U�4/��CY��.l��۷q*�g"�޼�q�=� � ǿ� ��0��ߴ����
ɩi��t
�ـ�v���˲�/4`��avW����x��r��)�GQ󖛢K`�0�U�"������i�R�y�x��ص�?"~�Ϝ�U�sA<��ơ������z���	�����]
0͐�]��&���	S��:�[�ow����A?��>װg�!�FJ�YՆ�SD�O�!�����a�q(��w�R�0�����,���&x�K��
�����/������/�Ң	D=�6�M�&�Wp�0�zi����d<L��aH���7;}��U,˴���� ���M�������z�� �@=b} ޏn�gR�MA�{g�:�iսd�c��P��g�~�Ҽ�ݲb�K3|��f�-!�КG�;(�Q}�u}�ͤJ�ZH�:�Y��t��BA���H�/4����N+��a����Q�¤��H%�ڎ}n+�z��9��ē��� S�5����q�Mё�H��\8<�|y�x�<�����˟R���/*`_�9��>{s$6�v���R� �Ӷ�c�Bo�8j���b��y[�v��y�Y;�Fvڃ(}�Y;�\��Ư�������a����;ʥ��vdi&�H�5�Jc~��� e^�Nl��$�����U*v���bG�!P)�I?��hrs� ��fx��m�(�l�9��R��'�0�(�'�HY�=��@�%^��ڏ�PL����G��tj�֧�DW�|�5JR������ h���;U�Hɦ�G�L}������S1��C28���U��-e3��`�Υ�sE��{��9塿��z�0f ý���m���5<���@_���<�s�<��MӢ�	����p�A_{ve]ȡ�s�Hd߀X,�flb�@��^�S�?�VcG�k���P�')})����'4�å�J��p��}S�Z_�a��iK��d��S,q�M�a�U��h��8�ّ��	ϻj�5~9����2ֵ��oܗs�⿿��(���Y�	-r9���Y�2��h\��5��aq���<a��XgNr�;ݠ�47Nn��8�j\Bߣ�W�Xv��?94Jۦ̥�T�(��ʅ��	��T<��EɾL̂;�����#�1Z�(:t�)�* ���e94����T_8�a� ����Y3ﰧ�Ud�f��Җe�5�Ȱ�#�$?:$���?�d��B��I��я*UlYB�p���v��6j/.�����V+1�R96�n8���y.��W��O�6r)��Θ��@��x����J�~����q]�R5<�^[*��X2��CX&�O6x��� _#���g��μ
,1��&g�.��ኾ@Յ�U��^rr��n3=��o�rɛ΀�T��Y�Ԯ��C��  �O
���j�VX��45%R���a�/de=�vK�zj�
4���g���_mW��T��`)��%W�U���ۿמfa!����ha�p�L��*�ӀF�T]�5v��E�l�h���	��b�x��9��~[`|6�5��eѨ�j�#�EC�Bc�2|$��q���}4�1�J��X�("�K���A��^+^�i�VN���ȶ�#�"��ޜ9�_���l)�0kV����aN�_��Y�*{1��k+,��l{�E2"��.�e��\ۆ�G�C���9,&:���D�E2�񝌔C&M\a�z��{�f4���?��yL}����O�Ϻ`�'ܛ"X���Ka����F���G�k�
����i�	|7w�����sDhї��npI�^���j�pR�h)OTy�H����A��j(�z�uD���Il�`���[""�y���Y��j��mA� ����}�ޥ(��ʕ�R�@��o��6��4g�N���6��2?m�-�ж��쀯%Ƭ�o�����������M�{���MK�$��ݓ�����)�T���O;jC�x��]Lp �fv[���~�^漙�1�	���H���w�8�4��u��R�p$���/�����B�b�����I�-T�U�L�&j������O��آ�8���tg���J�ф;�HΣJz6��B�mݘ/�'�?��f1��G�i� �{������i��	y��ѝ���г�_�C�틗Q�������C�T?)�C�D^��0��3㺪�� ���^p��@��ۛz�F )��*��k��}�����Xe?��X�(���.����ӒV����_����P*�v���b��?ŭm���&�x�8EB�p��а[�M��7�ʽR�rui�����n~���Q�^x��2D�f@�J�4�DG*���PS�[�s�K�����Z$ţ8������|?ra���2�ݽ���*7*���&����S��J 8-�U�|f����|?!�2�x:�ɔ<��je�A�0�]->���>�1�� �u.�=%h6����`W#��)��q�:���3CM���NA��$ �Ǚk4���s���$�d$�lRV1٨EO-?�r��A�G�5�tt����}������p�	i�Qie��	FA,�NLC�*[_� `�-�~nW�Y� Ye�e*�+�6&�ɷ5�K���Yf\�ME���'��X��JK���ɶ�fA�\	)�+8mV�N�����}��n��o�6mV�5,|Ĕ�.PN�?d�t1�b}_���c�&J?x"��m��2��V<��Yz�Z�7�Y[qb�n�]�T���z���)�1|�d��ev@�챬lK��	���?��2��
�8�y��MA�S�oK�M�j"ϼf1��nJU-��*yRߎCdN� P���hr���6���*������`��-{D�S�l���΃���ڬU��n���� iI!��9E�<�=�M}W�!�����z���o^"�I�ԣ��cG�fPu�:���q�{aTK�뫆���AÅ>��+����1��EU�-C�h�����\5����h� S�E˰SZW#����5�J`꫺m����8l��[��}��Xv\���U�U����!�O%�eq��V%}��5w��.)��>��"9^&�~���,�(7H�J�v�|�J<н��8���ח���d��5�/�| _]��S��ȸ�Z�zS���Zk��'9�����)��4�{�Α����HccCBv��5�r�q��
/y5