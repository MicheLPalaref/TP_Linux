��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������-��
1����yr1FUb��q�ej�IϢE^U�nA��a��"��� �AMF'�k-���޷n;m�o�}Z?��$Ĕ��L�h������g�Y]�)�}�"��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�?2zֺ�i�UCv�~��t_.> �KX����Q�!�N���k�
]�[�a���5�~��ѥ~�_!-�Ǵu�k0��s��@�b�L��Ih�.@4��I�~�l�*K��o��6Y{��� �U����rʽ��=�%�B��)� *z�h�	�ɳ�UN�I���yF��EԄxA?�·��0� ��٩E���$�z�����ϜE���
z3C���F�Q��
 D�=�*r�Ů�ߤ͔h��� �C��>'�K�j&�����i�'x�$��,�}>��	���~G�����+���og�b�Q}ȼ��l�GUX���讶�Qȹ��8�ɨ+9�Ф�P���� U�@s�p`�B�@�ob��Qٖ�d�� ])KOr�3��u�:f��
�N� �KЧ������\0Q�����w��Lk�}x���cBRo����@S��m����Ƹ��H'��JU�G�Leh�\Y �U2m���S���Q��$�G��X�R� 7)�6;;C���:�YSG�������S��pU˼��p�f'�Ȏ�6�Fe���k$J��������0L��#Л���Z��V�VW�*�24���4�E0?�$�)V����;�)�z�ϯ��?���y)�# 9@ ~�}{��'��G�8�0�<�y<��P�o٥�B�C�haZW�8���c��(�Q�%0ES�=�y�g��Q��m6%�"�ژJ��T������=/��¿꾄F@%]tS��2z8�\���D���۾��5�:��U���eWϠ�!s~*��I��X�Y�C��5Ů�љIt�����	o�D�`eO�pds&���J�RTv�U�Z�VX�O��4�N梻��X�Ǒ�^�fBP�)��¼��x:�>��:������-��+u��<��^��V�9�H��_M� ��A���9����:�W���3�C&֞��k`{�z��VH%]����:ղ��࿈eoY�ۧ�f&��#v0&V���wa��
qS��m���W.����>�r��!�=N��lFq��J`�r�Ap�`�!7��	�����*��r'�'.u�j�82��r^�x]���D���W�6��Z1'�@T(TD�i�N��׷=J}�($�� ��p�ۀ�x�������x�����%��c�����q��H��ນ����L#�>��qy��?�-(g�[_�?L7��皔�QR딁�Ś*�T.8��]N���]�c�}�M:� �r��"����b��8�?>���i��������ȴ���5l⣤���9�)�D��@Ō�u�-<�_8�O؈L�g�d2��POp#�R��(�v�?��V8ƅ6��b���#v�SI�#�Udo����?��x)�d�"~ps��{���U�|�+�4�X�}`��eAW�m���< u�c�S����s�&��F%2f��V�=C�c��YQq�-|�g���`�|tc�������E�s�n��`pM��C����M�B��SE�<{�Mw�Q�Z�-�u�J��A
�;b>�x��=��{���B�-ew3�#�;��,��ŕ���L�]�E{c�� �J�
��{�w�E�T{���Ϋ�!�h��^���;tq$�n��T���D���cuOyX��g���
Z`�wOJz+&bC�r�v^	��p9�8_8���A�3@-�>2�h��x]�L�w�Dbd��K�S5�qq-���N���S)��3�����_���`�W�Qqǵ|�		������	�x_�Md,X�J����v#�!���Cz1q��m��@�c_�Qѹ�U�&����r��kl������@�����3A��{'��6b�g�o�{\���gƂ�>�`ߎ�k���;ſ,,�r9v����պ��$ɽ/��$o�� ﵅�rEu�i~���{��Z����mP�T��	��j�fR�r��>M0��E�KBE��H�iC��
s����\]���3�g����e������?�f*ST�+��>��%�)y�dNR;^��?���D��m���>��Ko>�.�t�Dj�V�4Ol��q��'�@�{6�&O�)�!���"a1Tu��o9�=��8y�4�lW����k�D�� :h���&��<��/:?��`_�L�}���Ѿ�������>g�IEA�z�ڎ�	V���qS��sY�o�YԦq9Ğ�4���or�(�^��o&I?����M�=R�����7��W��}4N/�.�XމFy��-W�g�1}�Ud����z3�%&��M��Qd��S<3[�E�@�e&�L���<��4Uo���+d�~�X��i��]�gzv#_B�Ί���ڮ�4����ddS�^��Bi��N�M�N�
��mʋr.׊O=ϰޚT;�g���S�@���3����%�El#o���T�ڌ���C��
���?Zؤ*���'�h� r�a� �MgJƧ� |����ё��2�ԐA��*���}����kEW�~p&�wVL}nivjM?Ag��y�N13�EMXV
��9�d�z
t�7��G��e��D	�Ͳ7� 3�$�P����5��tfm�����Mz%�z����L���>��¾ғ���:�
��D2����:���D \�Ff;稣#��:8nwP���Zh�x?Γ���{;j�U���~B���k�ƾe;�tɔ������a����o.���E�S�&��^���A9���*�������l�p�_v��N��g���e^�$�!�R�?�_�X:0��SKq��@�i�w �1�Ŗ�W�3LF�[�����p�,�� n/QYY��'���M�
ޒ�Ap�b���}~,�ˆg��u����
�1!N���ZN�zHg��`��ս���%�?���Tm�>�)kK�
���%��X�.U+��n��C�"��K�v�nX��wa>�ϥ!A��┇g���^s,
�b�N"u��CC*��<�'A)�Uv��^�Nְ�&�@/\4&���;4�mN;��-�c-�2,�����o��T��������M2E>��yݦ_������3��^:�=S��rf�̻y��3]Qa�M�j4�%�Ǯ��Y�"~�Bc�<�����/�c!\�Y��1�sj�E܁�*��Y�v̮��(�"w�.X/u�n^]t�<��]�v��7�R�c�%�����;�t�[��M�	rL��1`\N0^o���]��6�.�<״��=����@pXP�Ց}�тͱ&�I�&�m@��}t�W1�©T.�q*(�6����أ�&���Mş������BΒ#�NI�C���A4B2��7 ��>����.^�<��Ƅ�8��E@gY�{.�0�˿����D!t�| �������i���W~�?��D�-��q���U�0#c}C�Ym���
�Y;@
1���[�ƇHM2N��觊��S0QѤ�]1-���hH�n@�P�I����������u�b�勆^�!�)B﹕D��Z)wqV�]�$�z�<&BN�������i�plEg���@�:2[�!��Z*��s��i�N�I����L���E� �FKv����q��߰�~S�g>|J�\�Ը�{�S����OQ?�e�W�v�A�{'6��<t�&{-?�E��� n~� �b�p��w�Ց
��*�E5���{��ҙl���Lu�3� )�zp��+����F'}Rܗ�e;6,AxA.��~������'�<�OH�K�Ώ���Dr"	S k�/��Li��k���E)��ӊ���t3�g[vPfc����ھ�8a��I����f�C���*"1a{��6B>�c�i}h���c�)���4�m���>cK�5<��_MÛ���@����{m\v��~�)KA�;Ak��a���dg!1��}q� �Z>�.�\eFI��_cRX�6Rdͅ�r�rJa��7����m|nUc~G�����<�O�p�:Ei�;��ܪ�'1q���8���7$��/�Aٙ �OG{��Ӧ�
��bVanЮ:���&�W��20�C3�*�l�~�:�Z���``+�m�]X�`1w�(;<'���Hz������������!E7�;G〯�اE��D����J�6�<.#�a,V��=c_[�-g���=����\Ȑ�ĞEL��=φ��T���vek�s:g#�z)%�pC������ȑ��I�ز:5@R+�I��	�������wb���K)��At��&����Ǧ*�-��|7@�� ����'�g���{� g�����|3��à�6�`�عso~(�I������t�#B�nA�+��K�+��`f״�#J�$n_�J�:�O��cPԢ��;FQ����q����r�X��Hf�n��'�w�v(9t0�ĉ�3;�@�i}�N4 އ��	�+�a<}m��;��#�k�r���2%Ee����������G���N<������7����jc~H=B�g]� ��a��S���F��*y�{��`��	�Zoq�.�W�
����$�OO�y!!�R��7����釦*R�}ȞӇE�KPB"(��{O츁S��_�	�J^��t9�T��m�Ő����Z~�=\���ch��v�e	�\1�([��}�(�j�eO#��B"�&���8�QIv#=hp
��7A�R3u��j����z�DډJ��t�I�;�J�"��M��\	ͺ���L���׀ld	��/��;�I�c�Q?�m#<���*oxEpAS��|a.�w�����hsq���u/�&�	�Ek�A��i�����3�v�69\����!�Ј-�V�Lru�r$�j`H{�O�.������$��'��]7K8{q֔��A�Lכs�K0�Db�7�J���\��-�P5T�YG�ڌ�&��Jj�dhd�u���午�\E���<mb�r)@~�x~��<����9/*B�e�j2?�J-�EL�8\�*Yfz��;{����.�?�
,[ejG]�`j���0���M��v���Sp��������.���^Po��:�Yf��s�bK�~Ě���t����W��h(���Z;R�.D�0P�.��8[4�-��ȫ� O���W�w0P�h��Z7c��۔]���m�j&c�%)w�=�z�eA�=��ݶ�a%ڔ�Cd�%�����=Բ�8��81��1��u'�+RG��08O�g0]jX��3/��r0��c�	`\�"[*ut�0�6KEn��C�zpw��� �WD���4hA��*i������`}������Ȏ���:��[3�3r�c�S|�o).Gw	���STɔ vﯘ��vv�����L`��w��|����֎�x��<��* nG�˙A���|�CA:�	#w/X)�8��#�¥��L�o�ߩ�0b&�JR%U XQ����إ!6����E� B��L��3`��I����][_��mю��|x��_*W䩓{�����~��[p�ޑ�ZTla�2�γ��Ac��}��wC[�RA�7T�vT"�C���[q��p���F��.�R�_ɀ�wZ3F�T�G��f4�TI�Jtm71�=j�Y%�#~#��L;-�ӻ� &�8���"s���I�l��+�����7>��N7�0לƝ���,�{�i�)N�!��P����#!���zH�o#µ<hMlI���ыV�IF>e�u+q��"���-���`
��ʌ%�+e��)� >�bnf7h/��p��F-�x����!]��^>X_�͠&�I hL�N)�O*7aw�:��9p�����o!J��� �ȆM� v�/ﾗ�uAн�1�ޚ֭",���I�� Y��p[4;���Mh���H�ʒO
u�Tm)y�+�6��{�W�*�
}��	�0^͵Yv�"�@S�p�0A>WfAZ�N�#��Г�X��	��o�2Bڢ�z`fACl(`��)�5/�u\�M,b�`S��ٙ(�A�j�����vw��*�9�a��/��*@s#I u+�*��nRG���x*�x
)2���������;p(7L|a���pv�ܒ�A���B�>=�Z��6��"7�PЂ��b�-0t�F����ۮ9�n`���)�Pc�&C�$⨒\,|bRȮ�Դ
�ʁu�?*f�~>Z�DxTq�t�ץ�=���ዸ �r�P��l�Y���8h��!SzT\����Uة��D~>���ɔ5A��s��Y��� �v�Hfj�1u���/c�xs-[�V"Ϗ�^�\4C��kt���)�80�UϜ�U/�H �a�L��xWn�9���H"\�\"�vg�u5O�	��YYRk�]��\�Z�O��	NF�q��c�'�v�D8hB�o��r*��FY@Iw�:?���L������#�M��������A�/������Ti����[��,INhx!&J2|f&�g�C�����<�=t{��Ä��4��]�k�D=?�9k�X�I\c��7WHI�������a��Pz�%#n�qj	7����w�yS6l��}�9��t�Ⱦ��A����o�u �酭��<�@����3�2I%�c�5�W���İ�O�h٠��( \���(��G8����(bc�Iy;~��,ll{���<�@�-���+#V||5�}�o���Fm�A�a�L���O`k��@m��?�%�����iq�tl��H��r!�.Qr�B�6��C����4_�^P��$�僨P�x��u���<��~+
LpV���}�z�����5�	0�RoG�͙YbI���%�*⬚���ƾF�J(�,��)����G�L�)�y�ILrWkKn_��2He�+7~,�NЖ)�q9���%�C	�N���4d�M�L��5��V~��LF�l@`շ������~K��%��u�cX��]b�����N���H^[s�$H��1Ж���֨Hj���q�P5Hĺ�
���vo3\LJ�J*
���/�c��^�_��݂r_�V�����6W���R�� �-,#���l ��U�v*��t`fa�A�A��ˤ,��|��¦=)?Y�]�)��󾁼��	i"t�r��:�z���+���)�SK3e����� T�����E��pxH��$$�m�$8D�\\�`��J��%��ȱ�O�Q��j�+;U̫~'�>�gn;�W�B��}[V���G�͒�o��vE����t���0���,���-�˼���	me=�؋*Ej��������h��Q��Y��*R��}I:l�Xp�A�)ͻ�}C�����4�� �A�me���ga�Y�ԗ-At�_�U8�&��3�G萏��o̶��%����{4�I���cD-.��n��K@(����%�,@�2�F�'-[�+�N!��quTjXjW閗Y<��+�Ĩ��Ba�T���̏ߍ��p����5g0R\ػ��?��Nd��~Cr}�\�;8�jv!��v�oT���?α�	[���ͪ�����A��ϴ�i�x��w�-�����s����eGV7[��/=���-o]�'�h�	�j����G<2�$nD�������ē�;�铀�a�m/�ߕc�0@\�qvR�|��b�*/(�H��m�99"�<��^�<{]��6[���X�i��u4��-�w�lck�s����a�ʑ�3?��^���n�f��y���؆-�l�Ȁ��63~h����^�p�l@7q�6凛na�f��úm��ue���<�5JU.,[�9�R�����C/X�$�s�\,��No�[4+�����lb��~yy���P	�d��1c�����E!����G
Lhl���'�ǁ����� ��ѨD��[�J��3�.�c��U� |��0������o����ԁ1=|���[�pX���A<.� =߸�Ӟ�d���\#_e|
�	Ns�_��Y¶y�y�����_lE��k����܈:�U����lupIj�,ge�s;y"$�K�{�Ŗ��0��i���p�*]p���w&�3��<祾잵�����?�^�*�%pG���#�@NÎx��z^s]p̛��.�[����&��������c�-��}^��rn�-�� �=�&����V,s-́�p��:��s!�l��Iz�[�h�Mn�_v ��q����!k	[$���E'�g�W���(�o����Q�e$L�qf�L��hpz.^�5T�ۣ�cu�su.L����[�#p�y�r��y๊�!ʀi���T̲�Wo�:�w�e4d1<��9���$n�d$�}X���I��ܛ����|Nh����Ow�P®�&�8��V�];�J�L�/~�R��QÖ+�o�^��~�M('�xW((7�uc�����B�E�1ULؽe �F�E*kK��c2��CC�Y;�lE�����<�OH'N�4B�VE�S�*���E�m�"D��%�����}�������Z�$���;��aF��a,�a�l/�c�V׃;��z�9�il�>&�>���jO�K� z��Ă�`�c���7�P��UP� �iv�md�������P?��7�L]�e��A5D��>|�2���dq�J�5�JT��^K`9(����u�p�\V(s$�v���+���_��ތ��`���9Ab�';9�Ư��$�����/�P��s8?>ǳ|B���n3rh�!�9k�L��9��=�ʶ�<<Hp�h]�Xek4q��@2Q���~�,�H���pq!�bu��V�z��~�~���a��2��pҰ��ms�ؐ�>��<��T���_���cp#�|u��i��|'���h����ă��4]�X��d�d��&!�2i�U�ADH�R�+c5YE�j��eE�OC� J��I�5�qd�ۜ�I5m���`��T�	oOt�_O��szr}Ȝ�V�|xU.[%U�X�C�l��*Q^}�y���K�}��V�9ȸ�[ MJ���a�.�_����fX<2�����b�lu�.��k���lg9<SX�ɜv��2�}MD���2��6	�ά5b��?���0��֏uiD���~��{\ �MbT�
g8L�$'�;�ȋ�e&�t����GA(i���,�p&��o�B"��'��CW��|��dˊ���%`�$�C�L���=�R����C˖��-����.�M&ك0Q:o���ت�1VG��dI����ɴ�GI��u�ߪU.|��W��M�g$�h�M�R�ֆ�����n哖r"WZ��*�]Q��K3�}6�0fH�Wq�W��lBH���B���J��z�O"qt�䷬gցW�i��~��
>F ��)A`�����&D�>k��[�<e���@��xev��vs�u������:����u\b�t���O;��>
Z�6�A�Q|����f�����JG����	r�2R�BL�wݎ���p4Mq���5���ʜbҴ��I5t�C���&���P��w����VF�~<��n����ͬ�,��2C���>���T���gy1�1��u�,��x����E��>��}��@K"�~�������BP��0��?jF<���.yc-R
C�ڸ���D����Z��<�a�P~�8������GJv�LL��q�"��p ��ج�8�����_+�a2%�v�ҝ���ڤK����ګ>�o��+}	s�쒿�4��Q+�!쥼��m)⼎&���X߰K�"t��z��Q�Z W���G�"��*k�eئw���T�0�HwP�s#rD�S-��+wH\i�K�b_��)����<��]H������$��".]'�̹U �'~|$�����D��>��"�8��/�S[�Y{Կ������5z�{{b!>� =�^�Ɋ�C���� ��&��NA��_n���%��M��	
ٛ��,�@�Z�J=7nV;Z�*�v�\�qm�a�TBy���D��	g��]�@duTv7hKP���]�Z3[�7��3ȇqǨЯw�#�p5Y-㧋n�}y�K���K�H��p��v���JN�UD;�Ӿ�K��-�~{�Ё`��ט�HqzOlf@5�>��ػKsUI���7k�d
�J�2)8=U;rT9�T�=�	U؜���LN$i�ʷ|�@K��nA8�m"aEbig�����/���)��V砓gL���H�v�U�K��Z���H�9��L��#$ۉL)�C�Z1�w�B��V@�<��$���r��n�9��c��g�(��	@���5+�=;4|�Ur�/����.Q�W�ԅ�"O����u�f�n[����04Z:(�x�k��#��%�}l���YdBni����ma-$?,�c* (��[���j�7���lWr༨ڨ��j��gəF��H������>���P��2\G�h��#nCY���p��9֏t�$F+�uB�k^���<-�Cv���涣t�X�ZL�m'��.*	V����t�Sס-��,/�X�)�Aw�y9֔��ҹi>����p4���1V�]ǲ��k������8�&����Q��c#��<�5"�i���l����DWش�U���͛5(�ճ��$�[B�T^&̯�	;��T n�����>8��4c]�F\���PN��bL t��;.A�:�!�������Y>�v�m��HAF�^b/� &j��{���7b���y^�e��F�}����,ka]�D	�:]"�����#���LM�a����hv��2�O$;�
2���"��^������Gz����d?T6"	�7�r�J��B��P]��A��؁��������D��`�8��&��	���lB}��'�~ko ��J�!YN�W�knL�N��j*��vgqDoHw�Z[<��2�����r2�[�u�Й��=/�O<�FSn���V�>�����e����Nt�� �#V���݅�'�9���(r�gjn�XĜL	R\@Ew�2��ި����<�?`�s�
�����T���b߹N(F',OG�e�}�Z�R�������]	.#%B9	Q���K�wsBZߤ��»��wќ��)���,!@�}7���Z�C�U��vu_C~U�e �.��R�����7Ǎ��y ��0��Tp-�LO���3��F��#�'S��9#��sO<X�e����^�Ckcj#��f�f0�l��%�e�%��@�-��꾪ZVԀ��΍����&n�&�q��2�j@�܉I��_ɣ<�[�˶T|�n!��Q���E>�"�(s+�=bir\Y����*� ��ͣ��!�|���/�p�!�<�n��;���X���2	�)QB?l�s�P�P� 7���
����SQfQ>2���V&�g�X@�u�M���#����	^;���စ����8:���
-�w��M�0�P��e�X�^�Ih�0L�]I�J����O�OI!��Y!��#c��TR|(�/oɑ��E%+['�N�`'���*Sx��~?��ݣuG�{����m��3ZW"�]ע�p$<y���	<���b�	���r?<�,Rd��l�G��Y�K��mL�pF�W��'�2v:��~f��	��԰�C��nO�~�FU���1��j�׾��p�V�n���E�sQu���}��}�ߴ�.\��O��fr�c��q�ʆ�W
�J�m�F !�+���=3Lb7`x]�{����*����hw7�R�Oؼ0V���`Y#�;犮�R���f�	��>ǐ����N�^�q��)D����*���ޘ%&��4(�ڤ��	:�I�����!X-q�-퀱�p�	����.8�#��4c^ ��v�RE�&�x/�~4�1�ߩ�l�U��u�#]t`�[��<XTGn5~~��qh]�J4�'�u�@���L�*�yS=�R��m���*�?��*��`H���W)�)��3uQ顉&�-=�!��HQ?�H�3�v}�K`�P��H����*&,1�q��4?�YA~4�Y�YW��~��:36��qv���=�i�GH�}���|�U�Y�� (�?�"쉱�/>1;�B��ءIG"\��!�]�H��#����EeUT[�*ޫ���>g�#��յIB�Cd[��p̔"f&�n��Ǭ]7P��sKOx�3��X��$�%�g�L�`��Ng�>���F�T� R'�B�J/c3�>��fNg����"��'���.j1��i>ϻes�u��{��rA16�<�M�_P�f
Y��8+2L(HQ�ʌ�3�����UaYk\}�@���R��1��i��,c�i� Pt�u8
�r�+媛P�MG�͟�Ic��`��'J��΀�L$D�r�x�'��k|@�Uy�lue`m����D���O���a��C|䝮.����I���I�Z��,�S
pUK	}��c��?\�ߤ��%�[�VA7U3dbA�!6�?/�踨��x"�D�}]L����3/k��T�Ȼ.�F������-��������NZ�6B+��I�G��%]���z1
��Ӷ��$/��f��ЪR(6�:X�[fy ..!k�@I~j�G�b�9:�<�İ�0ݝ!���s
K�T8K6��ᮽ`��_)�g�*�E�CX��t2�b9�o���n	�@�:R�w�8ן5�^�1��Y���/��m�Jx�#�8�z쨟��un�����rp�@�jh���lZI�d�߶i.��n�<���[�#V+X����<+���a��ɤ::�����jut�c�4�X��!E��@ �&�f�Q�*(*Z^���E���9&u=�]f5dǷ�D?�	�ۧ	&�����r�����������X�&��<��Q��P~Kz�Eli;��B�0Cg<
!���Ox�f��>е�ߪ�(�0yTY�T\+-	��G.��ݽ�wS����+��W~�qk���~� ڔVV$l`H��	M�q3J�Y�>�'|�a�\@���y���9���:�m�@��:���md������y���hHy:��fQ\�v�pa��e[�:[w[���Y�A���2KEx�$�E4cӝ���CBv�2�Ӛ��tQ=�"]��F�����3d�%�aUVg<����g ӝ�ɭ1ڛ����@�J�>�H���hڗBK�ү��ӯq�%E3��7�`+�%Udۻ/0kFk,Xm&j[?	��?G%�਒�I���[X����vHH�$�N�-A
Zc�O����xm�6Ԋ3J`Y�f5�A_&x����uw��[��ϔ�	~�aK� G�`p<Eq�~���,
��'�yFR�Kȃٗ~�3�Ql���-��kP~~���]q*����N�z�i�k��\\�%6�s��g��W/!d?��a��".|xPQ�;��Aλ�~�/��/��̸o��p��?A�D.���o\�H���l�r0����.�f��~��z�n���p&O�X���<6q�%m F�;��]C]�m��Ҝ|�P�ȋ�Bs�W>�cf��g����ŋ�RZ�˲��I3s�Qڰ�U�@����q�3U���C��H�F���-��	�Rr(����-���.�`%�L�zB8ˣ�
Hµo�W���zn��wT_Z�|�y�˯Q�nݩCgJJ���&v�U���C&�V�,�y1�όؼ�vg�o��ƶ�Q�{����$��E�ʵ2rl�-?��N��UӍ���2z�X��X�TD�v���!yT%Mo�i+K�z�1���h[�$a��ݨ&�cݢ4+�?v}�o3?����C��9?�PgFe���hbw͌2g\wQP�	8��~��l(z�!j�ܫ'�$��M}�ӛ_(�W�:�������Ԓ�V�,�u�4V���x�{���-f���,7�NHmc�-�i�Ԩ+m��JC]����E��Х#v�X�<��Zs7'CJI3�xDp�<P`X��̀[��o���W&;��2S���5�
�%� j�y'gN������f!�P:�SG���*��YEJ�qo�?q)'��a���[�� )��k{��X�r	$=>X�V5�v��Hf:�Tu�rI?�߁Ϯ�,l�^�M��"O�"�CdN�8�xä�=E��5���Ykƃ�?�^��5��wO� Lw-
s���,�7m{�j*#�T1ۘ�?���!fj����s�M[��Q>>�2Å�¼�6����Nc�Kb� 
��}�Y���4
�%��(��XZyթf������3
�:D&X��o?Z�x���*8��:֣�n?������2#�t��	E��JZ.E��[]�:�Sx8��\y?r�|���<'@�O�?W�˦�t��������$��ہ��S�u��k�w�"�����r���+�>�ؠ-�-�U>�`z9�g�an]���W�����oT<����{�ɨiS�r�!�bQ�w��w�KU��2;�?�Biѭj��*Ja�b�[E=��ar���
�+�d�#�^���'���e�
/I�J���|�(Up�n��i��	@�oojf�w�)���&DO�;�2�@���H��ݔ��	7�O;;��������۲,�9ꀆt�Nj���e��P�~u�l�O"VV�Lf�|�tD}��B��$QF��b%$��@���~d3��sA�s�E��Yx���p��1��MM���������얼	���z�T/k�r0�7��a��r�D�
߷���LY�jSc��x�H*@��ɉj^��,�ϸ�N��"��U`g���3�e�dkPW�.qi#3�e��d8N�F���-(������:�ߥ�z���`�Õ7��S?) 껠�Y{	Xd��g��Uw�z�=�ߙ��!Ǫ�TA�|�"�CWT���;���Z��^�WdM�b�W�6db��pH��f�TD��ⵣ����T0���A���1)^!ڒϨY�d])�CB�]+�dlt�uՠ��te��0�t�o	��+�B�I
 (&��ȋ�L�K+8/T}�j�Je���#��l7K ���S��p�Ķ�n͓&G��0�$����A1Ik�`y J<���BTo���!��YZ��RAq5�_�ԍ�Ki���V��D��L�nЀʊ�Pw'�$Xguô�ŉ���X�g-����wc~�+��7V�{oB��>5�>Z�nKk9�ː�ʜ�=�D��ǅ���19s1حx٤����N͘4��	�[؇Ҋ�I���7"d`Ie�
���:J�]s�l�T3y��o�|�g�Ջ����T������`�'������{讋���+;⒇�m�
����TU���Ά$��G/�B����,��4K�O3}�ը|3��Φ	tCA�Ϯ�!�wzIT�S7�S��x��G-�3�sDE�U} �p�)D�U�0Ū|t��^gf;~k��!Į@��H87���j�)��TeR=LG2BEj���k���� ^����z>��p"4rE��	{a2���vCE�9,�|K�j�E�Upq����`���U��SE2�2��k'[y3��E0��coW�i�Ûo�ɶ�Ԡ]00a>�L�#�a�����(�i���_��UƸD���yx���U�Z��t��!Й��º����x qo=vc���k����]��g��̣�V)�����É�nm��ʝ��%N�r�(m��M����E{ќ��0� -ǐ�Ē!���ɠ�X�RW�W��k@��`�}��z)j���碆�d_�c�o*���J�����mʖ<ت?##���S��~0��*���}|z>�N/��]�
�W�hh����1Mv��K\�v岧�^�0�]�T�[Kx�l�Ɩ:)�@�b�n�%��dq*�d�W5�h�Uh���_!h<kmg�R�.�[|������!�	vd���q�ႋ��h�q�D^����䚊$�2�4.*�h@c[-�*�q�ߢ�z�ȳV�V�8:1�jQ����}�Z��T<���Մ^�m:�uT��D`=2�n��A%�F
}�m=�@�׻��L)7ɱ��Y��#R~���8�ϰ�x�t��je���J�C��e��b[��<e�g�D��<Z�K�_h�t��F��"V_���$�Z���!)VH^���h�s����h��m�<s��^Mz�����H�nT�{3^:�t�����e�$W�_�:��?�E�9GI�#H�M?_�c�	�:��e��i�#s�Yۏ�껼�O*,��95�e(a5���.���ZJR:"N����ݭ0
'ߕq�ST��v �B+��	�&��u����%�]���r#���2d�0m<pY����Xbs*q��.�{���Ebܩ����L������RC���\�]���Nj��w��5����[)����#\@�9�Zo�ū@}�ջ�_ S:!.�EQ�P+��lħ�7R�H�R��6	��}#�<)��������)-�Bȯ�ۡ��2��ɹ�Kb.�������C{Rm5)
�@�z�1�����Ǯ��4t*[ ���]��9��Pe���7x��q-��1"�x�겣5�z�5�:F��>y;�6�@�&3�름։qů�)x�޾���,�r���2��h�ZX���.6EW�E�Bs�O��o\�Cv�)eM� 0i��"y�T&va��2мk�8ObG��A��M�^W��-� � �۳�|��MH�QkUj��?o��,���jb��MT<r�
���8IC����_�P����o��a�����m|:���6�m���:�Ŏ�$}�_-���3G"J�:���su�[KyԲʖ'�3lɯƍ�f�]��.F�E���dC<C�������r��b��XgY3���#�5�|��R� H9��g�\�Q �^J$�r��{�L
n�o)����j��F�k���S�����g��ފD�oq
�ٽ��b*IyU;O&����!�JJ������n�昜�"0�0��p�h��7{�
^��v���� =����P����ǴC���W�=��EU3�KY�,�.��	���Z� ڞ���G@�����z8�Q���D)���Mp,ip�|��
jl4j�o��W��v�:*v Z�&�����d�J�6ڬ��To}��c�l$�}Ȇ� ���,V+���{���J=�94����wj��4��>y�ӹ4˾��6����2$54�:�Xy!6�q���T������+uMuk�D�n	�fX��x�
a�Q��	b�o݅%X�W;MQ������|uJ���F�G�r�c�aD*I��-;�^[ȅAqO(�	���=��'g��\oe�X#�C�����ܘQ$��.ĉ�'�����4"
~���!�US=$X������7X�����Z���4�_�s�`�mT��v5��,�)��ڶ׹A����v�3�@�0�ٷ�+۷e̾�t4`�(BX�����q�I�H?'���9����?��Ǟ��T[����\��C�!尧H��m�u�1UO���pۣ��i��GR�4�s��N�z*�
/!��΋w���_��=k"}xoK$�Nx�@��D�
�nX�0�����;pG�?������?���s)D_#,�w���j�cا4�K��yv�-�5y,B	Zt"���!�r}�k;��[Ɂ8R3݀ ,;��b���С;_�8�v^�ѵͻ�p?�۸��QE��������@��ɑ9� �"92� lj�OxɑZO�w�L�� ^��ω�r:�E��5��L^�&��ߗ$m�A=,���^����k~�P��l��|��$�B�6�jQ��Y�l�8�p@,�������^�A[τ��� u�)ս��Z��
3�,i�޲ݭE#(EsY��Z��,LI(�>���qk���~��<�F�����0T|�:�z�j\t԰�e8�o����)�\�с�o͗]������"�B�r1��"�[l��ǭ��=��iܶ�^^������5�����~b��e�x��(��<�+��"nƆ_���yFj��t�V�p׳�"��}E�./�d� ��p�@�a�����S ٛ�;wQ���'fc���U�^a�pV��O.�٠�f�y��p�Z��fJZ1��)v�e��2�K��ԥd R<X'U��)���;47�A5 ��Lf�?)6���B;Y���E&�椨�J����%�4y�c �l����7��"��t"�C��w7�	$����a��`NK�4�	������w}��ގìA�N�o>wn�7[�2
�dq{Iݎ���[!�g��Z����j��)~W�Y�C%4�As�,H�k�X�M��1N�;1�8UX�Anu'��Ga��hJ�X��3~�_y���%A_���F'��ٰ�Vo��; SDc*#x��(��Ye�l/n�IjqSkÐ[?8D�G����[
AN	}�,W��`�ӏ-�� �S���S{�i9#F/~�:j#Y�pL���9��ҸR��9�{�k�������@;��h`(�M8�P}=����&������i��o�3�����{#�P���\�(���4����/�	�H��m�4�	޺��@��r�F��N>f�Y��y!�&H OTj��1���.�# ��XlT1�'g��1�Pޕ3� ���n<����#D#��db�D�>Τ�,㤛GSe!Sftk?U[��~�u��i���q"��`�cΠ\����2��p�ݲ���-gt������O�c�VX�Xq�fp%2�9*{��Y���i��6V�u∱�v��͌��P�U��O}I��_K�l��gHM������E���S�9�2�75��5
��Mk��ĕ��9�;.+�C���:�#y�
���MYxz27�d�Qv�|�l|��5�1ť�k.�ض}���X��J�^g�z�	{ �����T��֡�^�����7R#��a�Ұ���O�b��?N�S��C}(�Cr�I�Y�]ܓ��4�W5i��kz*" �8�#��a:�o��,�.qE�%ϲ�_�ː����z'U[�C�b��.f��rXˠ������xԋt"0��ɞG��2xeMJ�0ݵG���]�����=yP�����f������:ݷ*��RJ��{`�!�	K���Q,�.����K�B���_�(孝�R
r#t�j�`8�X���;
��(f�lv8_���P����(������5��&�ʗ=����&f��P��gN�(sz @�����YWƲ���c�=>�S�~�zެK��3�����ʛ����b��@O>;���j.w1��Gŝ����ă�)W�1j���:�-��p���� � f�z	�����Qbh'1�mpe���0���[�b��Q�PntH���r"�5��UaT>ɷDK�]X����[���� �}�^���U}'`9������j6��T�yF����o9��f`}f`��_����_��{>dqY���Y�+��سј���NuTbL�(�����LFGȼ���2r��?0o��w��/�� ��煮���I�����? ����,gԐh��V#u������pClh�4H��-�Be?��nl dt�#���@�{5�l��������H�����/���23K'��(��tu����ig��­�:h`���VX���JG��V�.}y��lz��\�6����jhqu9'|o��h9��D_X�yk�F)BEӢ�U�����582vQL�K˚�r =�	?[� ǎ�!��ްW�{K��6�x	�Q<��mf�Έ�4r��W3�b��Q�{Z��f��̕�0rLk�c���猹�h��βR��\�b]�*���$���_���_�rԽ0�%���j��8�f�d|��7]��G5��6i�B���ylg�%H`[I��%�0�i%Y�9<+�)��|�t�;�DA�w� ���}��5�4Z�W=l^�$J����J�f�8el�o�L����J�ܤ|��I�����|@LWu<q�6�-Z%�r�R�=΄�VИ	�2�xKt^{c�pC��'�f�01KCu6#%ۣ��/���E[�PR���ɤ��	׆�%Y0z�����N�@�n(��,��pt�|���4�\��,C����Ւ����\t��6�a����d+,�"=�#������x�>�!�nq��7�E2��I���� ����`�7A6n޶��8⼄[����\%�"����IY	�H�T��Iv�����`K5��������v��q���
�����sqs
Y|݇�0c䰕���xx�&<e�K��ÚDs�?���%3=�$Op#�t��KQ���n���Ρ+��VM��STKR��)S̈/3r H��,����\$2�cVb�輦U����.q^��z�Ql��#��:�1z��G��[:�����$��,���hT��	��N�p{��9�%@��Z�x�UI� �XuO`�޻6r�x�jSM�� =t���r�Ɏ��:AfP�Ǣ&%۸נ �nVȪr����`�s�4��	%���\C�v������B}#���W�u���0mIX�h��M�;��Z���c�y~>r,,�e� P��g�,z���}�� ��N3`�4�<0��00�޾4����$���$/ub�V	�ե��a���$���`!��S�R=,`
�	�<���X!N=�a��A���9иBk^g(]��tr#d�r�*���P��OXP�Uf8�S>�(������/��+n������o��WNm�UΑ��s����o˾^��"TX%�N�W��t6	j��h��U�zf�-�4�&���~�P�_���^�`{O-�T䚁姕�}IB+ss��t� Ŗ�gO����YM��2�s�����hM'�ϵ��q�kE��/�N4a ٬1l]T.���n&[m�3�"� 17K P�����I�w�r�=�2/^'���#b��\�T��r�1n���Mc�q
�i�C�*"Ӽ�DF%�M*؝�V]X.��Q��Q�E��SVT)X�B���{�W�Z��0oK�@V���`Q ,w5bf��r5��_`�����0R�J4��/U��"�eO� w�C-Ot<dAZ���Aľ��g$��i��r.c�Q��l*�z�����՜)�!��8����f�ܑ�(��ħ���NZЦ��tC�PÊ��z����2-�0�Gu&lG���?�T��ZL�xDt\ϯ���2����X����:��[�O� p�>b�c8&�ƹ-��g4�=C,�.��\N:b-�ƀQ���7�A��.l̳cO��x��&x�,0��N�Ӛ�7�Sh����K�m=� �Z}�5°�j���E�k謁�%Ա���}�z.�tϞ��5lIlf���j�*ZJ�͒Ɍ�P�g�y@��h���f��6��)�b��a��ʑ����m��(VX�F��ޓ��u�I�ߋ��d�x�Ҿ��̆�r�����=?��jLǥ�058��V�xPSV�F�نd�mpo�"R�4��nOL�A n'��I��^T�<y̵�/��-̎;&ԃ��=-'�{L�w?�u�@q����2Lyn��R0Uf��! ��hAݠ1~��$L�nj˓o-��Ǯ�����ǫet�2n�/L�!��o]#Ժ��1�!Uhì�(1P�QM��t�𞒔քhT"f��҃K�5�UO%?ՙ��ZtBM����f��\�0���-����uL���O��.���N#��X/F�\��l[�%쿿[�z�m�X�����4���b��[���M�j�lLy8�Gg���s*���ɤR:$Ř���mN^���p��%ĸ/���St����L�����M�hF��a�yHcc�����l���l�����l�-vQ �#��I�w��<���ռ^νѫ��`W�B�O��ϩu�Wyҿ�z�)"��K���ͮ)��	!\���=לD����/nլ"� u��B��CZe��7��kC����N}�����xF���ƶ[z�)=P�P�5O�3&L�V~��~�
��Z����>Iʹ���`u16��[�xU^VҼ�o�P�h�'_�q�����A�xA������]���i�G@왘�j�ݥ��`n�V��/m�o&�9��r���E�Y����e㱬���8i������)g8Y���e�K���LZD��a��7qx&dA���}�4, �0G���7�`��j����<��L�������-�o6��!&>�Q0�Wz�Sbk��T���*�̬)S��%�h����
�ylcxF%ǡp���vZ/I��$�k�ꛊ]O����~�9H���6�dH��	v�VyM))�u�� 	w;�"��Ne���M�W��*2�f��UMU �H������ؚ��z�%����W3�X��}ZN1��s�@Tv����AZ�]�K�</K�A�6/uv%'ׯ��z��-����R����Jj+J����g��ڍ\��sؾ���,�^��"�O�K)��1Bϥ��0� Yk���9��L;]P1��=�r6|wF+?�ܸ��
�}c�]�R�/��p��1	��$�����nx�ݬ�}T���,�)I������,���)�_�D�����r}k����8'�8s�.��4]�ʠ����� ���F�@���%�Gm���;���m��<L��C����Qi�-w�b�X=���RE��`ČͶs�Ov�R��&~#KƄ�Nz!-���8Y�r#�4��G��`:V9ԣtݭ�R~ʋ(ٷp�w""��'��l���ca��`{$3��H��p���%4��f�c��
j�r���	"�*ƇC\�	Mf)L�(|)�w��w���-5�܈~t�&FwA���#��lف�;�����T]�ɦ��[�ץa��ĭ�?F+љ��js����G�N�/�c�"�U��j�-C������ӆ���J}%_4�tI[!����XF���cB�g}��{5�SO"�=�Co]�u��8m�b�Is�VaC7����K��_�V�̪A��C�sj����l���]���s���<�x�J�:�s��:�F���{��97���cT�����(���� h�;�;D�}/uN�nv�	�Ef�-%&}\ڟ����󜈓��Wqp':��Ƃ��#��
	��];�Rl�ߺ�9SH�ç�����N�Y�3td�V���X���S�� �زbꏔ0�i�9dOUe���U��پ��U�I��@��{����4lؔ�1q�p�s�I�q$�qu��'���7�0����������"L!�?��)EC+CR��#�G���B�����?L)`�`Q��r�EO{��qI�s=g��Sá,i���SAs��\��[Z%��D��O���i���BE��C=�L��+	�H�Eh@�ى)�V��(X����Ma��*���8�I��=�fc�q�+P,ƈ@k;3�S�O�w���9����/iA�� ����P�$f���T��l^R��b�˙�(���SD�P�����j��a�K@8�q3B���3掵��b�!G�M����^g�L�<?-U�}c*l�K��TK�����ޕP�eM�HpV��G&Ҿ֞@�pyІ�}��7}��iȂ'�]_4#K%�6�������������	�>��F�������b�.���Sh&���.���y��hIx	p$$2{
���-��3���QI���$�8%���Cg ��IQ����Y�v���X��t�&���]x��.�W��.�ܖ�m5��g������~�sf�SC�|��Ƶ�k@����r��h	��Ul��s�.ԆǦ]^S����K��ʄ:g��f`t�$���M~Rj��I)���^���;	����so֏�y��|���;��;OA�����X�U�8�
���I�H.9���p�J�n�F�G7�6��O�������Wf�t�������-�h��b�;c��q�M�sf,){�?�R��2�c�v�ߓ(���e��3�z&g8W�s�G}�hd�]�3y�#�������Le��XLSv�4X��lL���@�~U9q�Ͼ�6���+�h�J�Æ�NI�פ������5=����ht��Ƒч��W����7���2��%T�C��ʖ/�1�?lU.�EQӖj��;��b��7�*�3\���,���&�IxPͿ�➇I.r�7�40��ב]����_i��=�C$2�p����w|���&�4^XӲ�V��4�53A�ݨ
p�t�]M��8<3�)QWVv^�-�p��e�C��V���X���z�=U��d��+�=���Y�
I��;NwV.#�>V�N��ezٺ*�G|^����N����q��-������}�-r�+;��_D�
��$�csbS)��^��Ҧª;tjt��u��1#��y� _O�1��I֤)���}�6F�+S��z-�g �WPi�^��Q��2��YG��5��E�Kk֘�u `a������l����L�0�K���KZ�B3�TX�:%�,p�3����b�	�O����R6Kw��ȸ6���qA��9믬����^_�(`�mw�	� n��ʱ���%�5uy�162?'�x
U����d����j	��~U_�ê݅mMQ8w8��6�ldz����g~�sT����T�.��^-rtko��#5��D��?��6������r��:�����L@vE3:�U�1��I�Z��`Q!L!��)L�<�f�X���]�Je�Y%��|��i�ƣ�n$(j�]�̅�x_���o�6
s�a������;bEa�-�)����Gז�EO��<��>�5�9�ϋq����L
\f(���Ig3���^- Ul�2�w�"m�>
��*��4�Vr�VLT=��25$����/HՑ� ,87ɀ�:6��7{�HE7�]0�L�I����>͍��Ns�@h�g�����０�y��2�<0>@3�ʤR�A�(������l|� ����7J�U��fm2�U���c/��7��N�8w��{W3�*�]���~��<��a�|���t�,��"D�&Ȫ�'�}m5�JGLݚ�Kjש�~�y����i�==ۢpg�bahIE���
�Å>*��-���@4#m�ت�����ݢ#x��G*x�$G�6�mBѥv�<��]�g;�#����	��ﲮ���E5E����\�A3֓⛎t�D�
��\�[�������M�kι�����8�����(��wm���ǨŐo����,ך��X�����k�K"��,-{�� �d����U�:p�yb�1�,W�P��K&�'��Pz2��������D���R��MA�!{���f�Q|F����P.rA�(�4�v9��g�ͮ���*`�����_�o砰�^y�"�"=���H� ?��z�3�x�gi���<�{�ٴ��	V���ʤ�����Ur	W�r0�'�,y�UJ���3�ZɡM�c��v/�@��X�����*(.��;���n?4��j��Y<j�`LC[��S����n��Ė����#�
i^j�3��v��r�y��{c49��ѱ��	���uG�	b�ņ�_[}z��=���i`�p���X�Ve����#����.ob�$2�E.�cF�����=��"�+�J�t#M�p��9�vN�M�GHA��SF�e�5鎯Np.2����!n���Z�3z;;��b��4J=_i�D�B����9�!�}�=x� '�����MO�%�0�^E4T�{���v��#X[��� '��5��Å��'�DdB!^xG]?� �`n/U���Z`Z�=�c�X^"�|J�X�n0F�+g`�a�&�S<4�){ds9�����+���^sm��)s!�r�͕h��_�L���߼���?g��{�a�z�:�j%�7����OG�h%�����vI���4X���?��[<@&�t�����?E+o�,�%�a�A'B2��ղo���� ^Clm���E��#�qJ�F)/�kn[����Nע����0{L�����Z�����pI�����(\�_�U�z�%�1-xP�s���=ɼ��$.y����K-u�]l�n3{ܒJJ�B(��L�?��P`}`�9s�愺"�ɡ0������_Y���T������ʅ �F���͖��nG=�@Q�Z"�|��O$��	m&�]r����DyЪeB�,��D�$�n[�w��L�Ǚ(6M5K,�=���E0w���o�B�pW~�#����fu޻(�Ǫ9N��w�=�ք%9��w���/�ɿ-�4����xcdWi�*�)}�,/����Ġ*3��(@�R�g1����p����Z�,z�nKo��,��\�E^s��R[HG���=v��<b��Pr��-j�Ov��'՚��/�)�p꿎]�����]�$v�@W��x�6��v�O�}�Z�2�rK������w m�D*�\N,�4�yމs�d~�h��R�y���.��`����K�w[�4���("ł�[�
�;�J�u4��
���m�zLn��G�t'A)路K�����|<���3�`d����xX>sX�M<ea
e3i�#�mʒ@�5��a�,~M�����aO���4�����4�=
�n|V�4�-���rJ)62tV���RK(�?߯��⦚�"�4���H	,XB�K��Bċ��4�m�+$IU�s_v��}���M��Ta�L9��|���jR�ӆ���x��m�4���}J����㰊r�W�(6a��9ƶj��÷��(ua���>`)�\\��J��U+�ZB�,M$F��q-��3Z�D��ʉ���7�(&��)��=��T�U8�e�D����
k��Q��|M�-��>��{�!�'븪/�����'��耈'�jn�55�����˽:�	�&�j���/�ew6C�g���� k�.[Fzx��\����o��x3�@-��_�m�*?�1����_��W��J"���l=L:�&��?�>�����j���������6p��P��ϰ���k%s�/�i��p�����)���[��ؠ��;�ΏSA�����%�g��5�4`�(w�)�\쬼��޼h���������ؘ�����j,R+.5q��i2j���!Z�҉.�ˢ{���N#�²-�Q"��7v�#JD��&U�����p0 �u���>]0М!^����t;�l�
�Gr�9.���S�W�p�f,dJ֦����%r};j	L�/�^|�Or��t`"o�����O �h����"9���;���4_��/�F���]�%N:_�q��0�:f���?�����pWb)6wbC�M���ڹV�Q�&io��g|�#[oIrE� ��I��� Ah,��nw��E��mX=w
$�~͘��F��iԌ(���I�y��!�������������"F0�]�g����	���^�x�T-���ȀJ�2#p�}��1�=j���b�����>�����-�쥁ɷ]�eZB�ru��%�~R � J|�Z��4>5���^]Hd�p�=�~���|jC�o�(�fo��|+�?��A@S4��j����]�v�qJu��o�@�*�N>��N~��UT�ጒ����w��~�	P ̢θ�uK_�	x#
�͐`?MP������í�4�rD��ݞU5��#�E����eǖl:Hb�MH��d���	�W�|�gt��c�Z�F{��YEk�rN��ݯ��ݙc3f�/X�-O�.HF�u]���	�e�]ۮmn+Umh�6k�a	�	�8�л�{�>��"��r��^�Jy ���=Uߖ�I��fF���1J������I	�G>�����+cEg����$@�)�Y��@ �M�]�/2�L��L1����2���&M'ڤ(�)���u��N0�mh?��&���6����@���I=�|��ʐ��ŎTͣG��;�j.W�����y\��QD��EE��5�Q ��A���V���&W�U���a���HN9�y���+��H#�u�a5�P�X�������dʐ�v����5���g��3��t.3�?�!.U1]���gL�m�c�������i�#��n�p/��-��ϙ}��b��"*gTU؏���\�b�$��:J�D3�=�����y�n�_JCc+A��.'r�BG���Q0g
�	��X� E3ƨ��v�K G�e��@&jFJY�NC���o��d�����_���#��8I�ND�c��ՐD��Yy�=m$�]�ĩ	��9��Q���߈9įs@p��������!�%�9~���Jf=�۴�&�m����3ш)~6l?|�z�<�C{p���W���Ɏ�77NҨ�e
w=Ҝu�i��>m6��u��d��1u�P߇�Xߣ��8o�H�K�/G�AM�~!�\�v��PcAj�CY�F{"V��+C������3�JK, i$��Z��Bl�HD#�&/M��93���:R�w�tҝۆűϵ�������o"�1���N��.�`[� p��K�ݱ{idV�������r9�?��$���w�-����퉕������X8���7�����[��!�d;f�#�g��/�����I���c����8�a��{�O���c԰��I�u��oW:I<6R����)��
�m�Ƶ����7�A��ɃNTy���00mz�&"�)5O��~�y)� <�u���c�����Un'JrǱ�v�Q��D�>��OF����rq��Nc�`5+��a�ab
�DuI�����r�7Ԛ���t�u3�%Ob�@`M�e�
[���\yV	��u��s͗Ga������Q����4Bjy��A	��3��J��S����V���ġ����*<핯i+����y��wW�(�����y���'����#�R�|ܸ��zWȿ����W?����C&��,��P`;�(,�����ˀQ��P����gC`k�aK%&��G�A�-1���;��ֹ�������aږ�<�Ӓ;ֆ�Bh�+u�1����i�A�?�C����a��������Ye4y�����Ć�Bc	֖*��-����v(�����f�*��s���T��ݱdݪ��w��$]m�/��(�p��
��᜾\��-�6�U��9PO���%��ã�ض���%�n��7����ex3��^��p��>o�%�U�]��N4��X�aJ�߶���(8'���r E�x�Ŧ	!�4,l>?D�����g�(�)"��%�n�?B�zMI�hM%�b1 i0btQ�ӓ% �4(<�<�AA3A"�{m]�C�>�������o����i0j-�0�|���{�Et������f�!ۅ� =�*4�ד7�;��('�M������)m��k���6<Zfs�6�ŋva^p��GD������E�w]]Fj� '�h?����*E����'߁�~��
�׋.{/	ٙ����Y�N2������m9|J��s�SE